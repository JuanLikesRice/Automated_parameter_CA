module BRAM_AUTO (
    input wire clk,           // Clock signal 
    input wire [15:0] addr,    // Address input (8 bits)
     input wire we,            // Write enable signal
    input wire [7:0] write_data, // Data input (8 bits)
    input wire enable,        // Enable signal for read and write operations
    output reg [7:0] read_data // Data output (9 bits)
);
  reg [7:0] memory [0:65535]; // 65536x8-bit Block RAM

    reg [7:0] read_data_buff1, read_data_buff2, reg_last_written_data, reg_last_written_addr;
    initial begin
reg_last_written_data <= 8'b0;
reg_last_written_addr <= 8'b0;
read_data_buff1 <= 8'h00;
read_data_buff2 <= 8'h00;
read_data <=   8'h00;


    memory[0] <=  8'h77;        memory[1] <=  8'h6f;        memory[2] <=  8'h72;        memory[3] <=  8'h64;        memory[4] <=  8'h31;        memory[5] <=  8'h4b;        memory[6] <=  8'h68;        memory[7] <=  8'h67;        memory[8] <=  8'h76;        memory[9] <=  8'h73;        memory[10] <=  8'h64;        memory[11] <=  8'h62;        memory[12] <=  8'h6e;        memory[13] <=  8'h73;        memory[14] <=  8'h6a;        memory[15] <=  8'h61;        memory[16] <=  8'h61;        memory[17] <=  8'h79;        memory[18] <=  8'h67;        memory[19] <=  8'h76;        memory[20] <=  8'h62;        memory[21] <=  8'h6e;        memory[22] <=  8'h61;        memory[23] <=  8'h74;        memory[24] <=  8'h6f;        memory[25] <=  8'h6b;        memory[26] <=  8'h6a;        memory[27] <=  8'h68;        memory[28] <=  8'h63;        memory[29] <=  8'h67;        memory[30] <=  8'h76;        memory[31] <=  8'h64;        memory[32] <=  8'h73;        memory[33] <=  8'h77;        memory[34] <=  8'h6f;        memory[35] <=  8'h72;        memory[36] <=  8'h64;        memory[37] <=  8'h34;        memory[38] <=  8'h73;        memory[39] <=  8'h63;        memory[40] <=  8'h76;        memory[41] <=  8'h63;        memory[42] <=  8'h62;        memory[43] <=  8'h61;        memory[44] <=  8'h62;        memory[45] <=  8'h61;        memory[46] <=  8'h62;        memory[47] <=  8'h61;        memory[48] <=  8'h62;        memory[49] <=  8'h61;        memory[50] <=  8'h62;        memory[51] <=  8'h62;        memory[52] <=  8'h61;        memory[53] <=  8'h62;        memory[54] <=  8'h61;        memory[55] <=  8'h62;        memory[56] <=  8'h61;        memory[57] <=  8'h62;        memory[58] <=  8'h2c;        memory[59] <=  8'h6d;        memory[60] <=  8'h73;        memory[61] <=  8'h6b;        memory[62] <=  8'h64;        memory[63] <=  8'h6c;        memory[64] <=  8'h70;        memory[65] <=  8'h5b;        memory[66] <=  8'h3b;        memory[67] <=  8'h73;        memory[68] <=  8'h6c;        memory[69] <=  8'h64;        memory[70] <=  8'h70;        memory[71] <=  8'h76;        memory[72] <=  8'h63;        memory[73] <=  8'h5b;        memory[74] <=  8'h78;        memory[75] <=  8'h76;        memory[76] <=  8'h63;        memory[77] <=  8'h5b;        memory[78] <=  8'h78;        memory[79] <=  8'h70;        memory[80] <=  8'h6f;        memory[81] <=  8'h20;        memory[82] <=  8'h62;        memory[83] <=  8'h61;        memory[84] <=  8'h72;        memory[85] <=  8'h74;        memory[86] <=  8'h74;        memory[87] <=  8'h62;        memory[88] <=  8'h61;        memory[89] <=  8'h72;        memory[90] <=  8'h74;        memory[91] <=  8'h78;        memory[92] <=  8'h61;        memory[93] <=  8'h74;        memory[94] <=  8'h6b;        memory[95] <=  8'h73;        memory[96] <=  8'h68;        memory[97] <=  8'h63;        memory[98] <=  8'h66;        memory[99] <=  8'h69;        memory[100] <=  8'h77;        memory[101] <=  8'h68;        memory[102] <=  8'h61;        memory[103] <=  8'h69;        memory[104] <=  8'h6a;        memory[105] <=  8'h78;        memory[106] <=  8'h5d;        memory[107] <=  8'h65;        memory[108] <=  8'h6b;        memory[109] <=  8'h6f;        memory[110] <=  8'h39;        memory[111] <=  8'h64;        memory[112] <=  8'h75;        memory[113] <=  8'h38;        memory[114] <=  8'h79;        memory[115] <=  8'h20;        memory[116] <=  8'h61;        memory[117] <=  8'h64;        memory[118] <=  8'h76;        memory[119] <=  8'h73;        memory[120] <=  8'h65;        memory[121] <=  8'h66;        memory[122] <=  8'h77;        memory[123] <=  8'h65;        memory[124] <=  8'h64;        memory[125] <=  8'h63;        memory[126] <=  8'h37;        memory[127] <=  8'h63;        memory[128] <=  8'h67;        memory[129] <=  8'h78;        memory[130] <=  8'h63;        memory[131] <=  8'h75;        memory[132] <=  8'h68;        memory[133] <=  8'h69;        memory[134] <=  8'h6a;        memory[135] <=  8'h77;        memory[136] <=  8'h69;        memory[137] <=  8'h64;        memory[138] <=  8'h66;        memory[139] <=  8'h68;        memory[140] <=  8'h75;        memory[141] <=  8'h76;        memory[142] <=  8'h64;        memory[143] <=  8'h62;        memory[144] <=  8'h66;        memory[145] <=  8'h6a;        memory[146] <=  8'h6e;        memory[147] <=  8'h6b;        memory[148] <=  8'h6a;        memory[149] <=  8'h65;        memory[150] <=  8'h38;        memory[151] <=  8'h66;        memory[152] <=  8'h37;        memory[153] <=  8'h67;        memory[154] <=  8'h79;        memory[155] <=  8'h76;        memory[156] <=  8'h63;        memory[157] <=  8'h68;        memory[158] <=  8'h69;        memory[159] <=  8'h6a;        memory[160] <=  8'h33;        memory[161] <=  8'h65;        memory[162] <=  8'h67;        memory[163] <=  8'h79;        memory[164] <=  8'h72;        memory[165] <=  8'h64;        memory[166] <=  8'h62;        memory[167] <=  8'h6e;        memory[168] <=  8'h63;        memory[169] <=  8'h7a;        memory[170] <=  8'h6a;        memory[171] <=  8'h6f;        memory[172] <=  8'h66;        memory[173] <=  8'h78;        memory[174] <=  8'h6a;        memory[175] <=  8'h69;        memory[176] <=  8'h63;        memory[177] <=  8'h68;        memory[178] <=  8'h62;        memory[179] <=  8'h6e;        memory[180] <=  8'h6d;        memory[181] <=  8'h63;        memory[182] <=  8'h73;        memory[183] <=  8'h6c;        memory[184] <=  8'h6b;        memory[185] <=  8'h6a;        memory[186] <=  8'h69;        memory[187] <=  8'h68;        memory[188] <=  8'h76;        memory[189] <=  8'h75;        memory[190] <=  8'h69;        memory[191] <=  8'h64;        memory[192] <=  8'h68;        memory[193] <=  8'h75;        memory[194] <=  8'h67;        memory[195] <=  8'h79;        memory[196] <=  8'h62;        memory[197] <=  8'h68;        memory[198] <=  8'h65;        memory[199] <=  8'h6a;        memory[200] <=  8'h72;        memory[201] <=  8'h6b;        memory[202] <=  8'h6a;        memory[203] <=  8'h6f;        memory[204] <=  8'h64;        memory[205] <=  8'h67;        memory[206] <=  8'h69;        memory[207] <=  8'h75;        memory[208] <=  8'h69;        memory[209] <=  8'h67;        memory[210] <=  8'h76;        memory[211] <=  8'h79;        memory[212] <=  8'h75;        memory[213] <=  8'h67;        memory[214] <=  8'h78;        memory[215] <=  8'h68;        memory[216] <=  8'h63;        memory[217] <=  8'h20;        memory[218] <=  8'h20;        memory[219] <=  8'h20;        memory[220] <=  8'h78;        memory[221] <=  8'h76;        memory[222] <=  8'h20;        memory[223] <=  8'h63;        memory[224] <=  8'h78;        memory[225] <=  8'h67;        memory[226] <=  8'h79;        memory[227] <=  8'h63;        memory[228] <=  8'h75;        memory[229] <=  8'h68;        memory[230] <=  8'h6a;        memory[231] <=  8'h6b;        memory[232] <=  8'h61;        memory[233] <=  8'h6c;        memory[234] <=  8'h78;        memory[235] <=  8'h76;        memory[236] <=  8'h70;        memory[237] <=  8'h6f;        memory[238] <=  8'h69;        memory[239] <=  8'h6a;        memory[240] <=  8'h69;        memory[241] <=  8'h68;        memory[242] <=  8'h6a;        memory[243] <=  8'h62;        memory[244] <=  8'h77;        memory[245] <=  8'h65;        memory[246] <=  8'h6e;        memory[247] <=  8'h61;        memory[248] <=  8'h66;        memory[249] <=  8'h6d;        memory[250] <=  8'h64;        memory[251] <=  8'h6b;        memory[252] <=  8'h6d;        memory[253] <=  8'h76;        memory[254] <=  8'h6c;        memory[255] <=  8'h63;        memory[256] <=  8'h6f;        memory[257] <=  8'h64;        memory[258] <=  8'h69;        memory[259] <=  8'h75;        memory[260] <=  8'h68;        memory[261] <=  8'h73;        memory[262] <=  8'h66;        memory[263] <=  8'h65;        memory[264] <=  8'h62;        memory[265] <=  8'h6e;        memory[266] <=  8'h64;        memory[267] <=  8'h73;        memory[268] <=  8'h63;        memory[269] <=  8'h6b;        memory[270] <=  8'h20;        memory[271] <=  8'h78;        memory[272] <=  8'h6a;        memory[273] <=  8'h78;        memory[274] <=  8'h63;        memory[275] <=  8'h73;        memory[276] <=  8'h64;        memory[277] <=  8'h66;        memory[278] <=  8'h6b;        memory[279] <=  8'h64;        memory[280] <=  8'h6e;        memory[281] <=  8'h6d;        memory[282] <=  8'h64;        memory[283] <=  8'h73;        memory[284] <=  8'h63;        memory[285] <=  8'h6b;        memory[286] <=  8'h78;        memory[287] <=  8'h6c;        memory[288] <=  8'h6f;        memory[289] <=  8'h66;        memory[290] <=  8'h6a;        memory[291] <=  8'h69;        memory[292] <=  8'h61;        memory[293] <=  8'h62;        memory[294] <=  8'h6e;        memory[295] <=  8'h20;        memory[296] <=  8'h78;        memory[297] <=  8'h6b;        memory[298] <=  8'h6d;        memory[299] <=  8'h20;        memory[300] <=  8'h6f;        memory[301] <=  8'h63;        memory[302] <=  8'h76;        memory[303] <=  8'h73;        memory[304] <=  8'h64;        memory[305] <=  8'h69;        memory[306] <=  8'h66;        memory[307] <=  8'h68;        memory[308] <=  8'h65;        memory[309] <=  8'h71;        memory[310] <=  8'h6a;        memory[311] <=  8'h77;        memory[312] <=  8'h62;        memory[313] <=  8'h65;        memory[314] <=  8'h6e;        memory[315] <=  8'h20;        memory[316] <=  8'h6d;        memory[317] <=  8'h64;        memory[318] <=  8'h73;        memory[319] <=  8'h6c;        memory[320] <=  8'h76;        memory[321] <=  8'h6b;        memory[322] <=  8'h63;        memory[323] <=  8'h78;        memory[324] <=  8'h20;        memory[325] <=  8'h6f;        memory[326] <=  8'h78;        memory[327] <=  8'h69;        memory[328] <=  8'h63;        memory[329] <=  8'h6a;        memory[330] <=  8'h76;        memory[331] <=  8'h64;        memory[332] <=  8'h66;        memory[333] <=  8'h65;        memory[334] <=  8'h71;        memory[335] <=  8'h6e;        memory[336] <=  8'h20;        memory[337] <=  8'h64;        memory[338] <=  8'h6d;        memory[339] <=  8'h73;        memory[340] <=  8'h6c;        memory[341] <=  8'h63;        memory[342] <=  8'h78;        memory[343] <=  8'h6b;        memory[344] <=  8'h20;        memory[345] <=  8'h6f;        memory[346] <=  8'h78;        memory[347] <=  8'h63;        memory[348] <=  8'h76;        memory[349] <=  8'h6a;        memory[350] <=  8'h64;        memory[351] <=  8'h62;        memory[352] <=  8'h71;        memory[353] <=  8'h77;        memory[354] <=  8'h65;        memory[355] <=  8'h6e;        memory[356] <=  8'h6d;        memory[357] <=  8'h64;        memory[358] <=  8'h6c;        memory[359] <=  8'h73;        memory[360] <=  8'h2c;        memory[361] <=  8'h76;        memory[362] <=  8'h63;        memory[363] <=  8'h78;        memory[364] <=  8'h20;        memory[365] <=  8'h63;        memory[366] <=  8'h6f;        memory[367] <=  8'h69;        memory[368] <=  8'h76;        memory[369] <=  8'h68;        memory[370] <=  8'h73;        memory[371] <=  8'h64;        memory[372] <=  8'h62;        memory[373] <=  8'h71;        memory[374] <=  8'h77;        memory[375] <=  8'h65;        memory[376] <=  8'h6e;        memory[377] <=  8'h64;        memory[378] <=  8'h6b;        memory[379] <=  8'h73;        memory[380] <=  8'h76;        memory[381] <=  8'h6f;        memory[382] <=  8'h63;        memory[383] <=  8'h20;        memory[384] <=  8'h76;        memory[385] <=  8'h69;        memory[386] <=  8'h75;        memory[387] <=  8'h69;        memory[388] <=  8'h68;        memory[389] <=  8'h63;        memory[390] <=  8'h78;        memory[391] <=  8'h69;        memory[392] <=  8'h6f;        memory[393] <=  8'h76;        memory[394] <=  8'h73;        memory[395] <=  8'h64;        memory[396] <=  8'h61;        memory[397] <=  8'h64;        memory[398] <=  8'h6e;        memory[399] <=  8'h77;        memory[400] <=  8'h71;        memory[401] <=  8'h6b;        memory[402] <=  8'h6c;        memory[403] <=  8'h73;        memory[404] <=  8'h76;        memory[405] <=  8'h6e;        memory[406] <=  8'h62;        memory[407] <=  8'h20;        memory[408] <=  8'h64;        memory[409] <=  8'h66;        memory[410] <=  8'h6a;        memory[411] <=  8'h6b;        memory[412] <=  8'h71;        memory[413] <=  8'h64;        memory[414] <=  8'h77;        memory[415] <=  8'h65;        memory[416] <=  8'h6e;        memory[417] <=  8'h62;        memory[418] <=  8'h20;        memory[419] <=  8'h64;        memory[420] <=  8'h73;        memory[421] <=  8'h76;        memory[422] <=  8'h68;        memory[423] <=  8'h64;        memory[424] <=  8'h61;        memory[425] <=  8'h71;        memory[426] <=  8'h77;        memory[427] <=  8'h6a;        memory[428] <=  8'h65;        memory[429] <=  8'h6e;        memory[430] <=  8'h64;        memory[431] <=  8'h20;        memory[432] <=  8'h61;        memory[433] <=  8'h63;        memory[434] <=  8'h62;        memory[435] <=  8'h68;        memory[436] <=  8'h64;        memory[437] <=  8'h61;        memory[438] <=  8'h77;        memory[439] <=  8'h71;        memory[440] <=  8'h6e;        memory[441] <=  8'h20;        memory[442] <=  8'h62;        memory[443] <=  8'h73;        memory[444] <=  8'h76;        memory[445] <=  8'h61;        memory[446] <=  8'h67;        memory[447] <=  8'h76;        memory[448] <=  8'h68;        memory[449] <=  8'h67;        memory[450] <=  8'h61;        memory[451] <=  8'h73;        memory[452] <=  8'h6a;        memory[453] <=  8'h6b;        memory[454] <=  8'h63;        memory[455] <=  8'h78;        memory[456] <=  8'h76;        memory[457] <=  8'h6e;        memory[458] <=  8'h73;        memory[459] <=  8'h64;        memory[460] <=  8'h20;        memory[461] <=  8'h66;        memory[462] <=  8'h62;        memory[463] <=  8'h64;        memory[464] <=  8'h61;        memory[465] <=  8'h73;        memory[466] <=  8'h76;        memory[467] <=  8'h67;        memory[468] <=  8'h63;        memory[469] <=  8'h79;        memory[470] <=  8'h7a;        memory[471] <=  8'h78;        memory[472] <=  8'h79;        memory[473] <=  8'h75;        memory[474] <=  8'h20;        memory[475] <=  8'h69;        memory[476] <=  8'h6a;        memory[477] <=  8'h64;        memory[478] <=  8'h66;        memory[479] <=  8'h6b;        memory[480] <=  8'h61;        memory[481] <=  8'h64;        memory[482] <=  8'h63;        memory[483] <=  8'h78;        memory[484] <=  8'h68;        memory[485] <=  8'h20;        memory[486] <=  8'h67;        memory[487] <=  8'h61;        memory[488] <=  8'h68;        memory[489] <=  8'h75;        memory[490] <=  8'h64;        memory[491] <=  8'h73;        memory[492] <=  8'h69;        memory[493] <=  8'h6a;        memory[494] <=  8'h61;        memory[495] <=  8'h6b;        memory[496] <=  8'h63;        memory[497] <=  8'h62;        memory[498] <=  8'h61;        memory[499] <=  8'h72;        memory[500] <=  8'h73;        memory[501] <=  8'h68;        memory[502] <=  8'h64;        memory[503] <=  8'h66;        memory[504] <=  8'h67;        memory[505] <=  8'h73;        memory[506] <=  8'h68;        memory[507] <=  8'h64;        memory[508] <=  8'h66;        memory[509] <=  8'h68;        memory[510] <=  8'h64;        memory[511] <=  8'h6a;        memory[512] <=  8'h68;        memory[513] <=  8'h62;        memory[514] <=  8'h67;        memory[515] <=  8'h63;        memory[516] <=  8'h61;        memory[517] <=  8'h66;        memory[518] <=  8'h73;        memory[519] <=  8'h79;        memory[520] <=  8'h67;        memory[521] <=  8'h6b;        memory[522] <=  8'h75;        memory[523] <=  8'h64;        memory[524] <=  8'h68;        memory[525] <=  8'h62;        memory[526] <=  8'h77;        memory[527] <=  8'h76;        memory[528] <=  8'h67;        memory[529] <=  8'h61;        memory[530] <=  8'h66;        memory[531] <=  8'h64;        memory[532] <=  8'h74;        memory[533] <=  8'h75;        memory[534] <=  8'h66;        memory[535] <=  8'h79;        memory[536] <=  8'h67;        memory[537] <=  8'h69;        memory[538] <=  8'h75;        memory[539] <=  8'h68;        memory[540] <=  8'h6c;        memory[541] <=  8'h6a;        memory[542] <=  8'h62;        memory[543] <=  8'h6b;        memory[544] <=  8'h68;        memory[545] <=  8'h76;        memory[546] <=  8'h67;        memory[547] <=  8'h63;        memory[548] <=  8'h66;        memory[549] <=  8'h78;        memory[550] <=  8'h64;        memory[551] <=  8'h74;        memory[552] <=  8'h75;        memory[553] <=  8'h79;        memory[554] <=  8'h69;        memory[555] <=  8'h75;        memory[556] <=  8'h68;        memory[557] <=  8'h6c;        memory[558] <=  8'h6a;        memory[559] <=  8'h6b;        memory[560] <=  8'h67;        memory[561] <=  8'h6a;        memory[562] <=  8'h63;        memory[563] <=  8'h66;        memory[564] <=  8'h68;        memory[565] <=  8'h64;        memory[566] <=  8'h67;        memory[567] <=  8'h72;        memory[568] <=  8'h79;        memory[569] <=  8'h74;        memory[570] <=  8'h66;        memory[571] <=  8'h75;        memory[572] <=  8'h79;        memory[573] <=  8'h69;        memory[574] <=  8'h68;        memory[575] <=  8'h6c;        memory[576] <=  8'h62;        memory[577] <=  8'h6d;        memory[578] <=  8'h76;        memory[579] <=  8'h6e;        memory[580] <=  8'h63;        memory[581] <=  8'h66;        memory[582] <=  8'h68;        memory[583] <=  8'h64;        memory[584] <=  8'h74;        memory[585] <=  8'h75;        memory[586] <=  8'h67;        memory[587] <=  8'h79;        memory[588] <=  8'h69;        memory[589] <=  8'h68;        memory[590] <=  8'h75;        memory[591] <=  8'h6a;        memory[592] <=  8'h6c;        memory[593] <=  8'h62;        memory[594] <=  8'h6d;        memory[595] <=  8'h76;        memory[596] <=  8'h6e;        memory[597] <=  8'h63;        memory[598] <=  8'h66;        memory[599] <=  8'h68;        memory[600] <=  8'h67;        memory[601] <=  8'h79;        memory[602] <=  8'h68;        memory[603] <=  8'h75;        memory[604] <=  8'h6a;        memory[605] <=  8'h6e;        memory[606] <=  8'h2c;        memory[607] <=  8'h77;        memory[608] <=  8'h6f;        memory[609] <=  8'h72;        memory[610] <=  8'h64;        memory[611] <=  8'h34;        memory[612] <=  8'h20;        memory[613] <=  8'h6e;        memory[614] <=  8'h76;        memory[615] <=  8'h63;        memory[616] <=  8'h61;        memory[617] <=  8'h64;        memory[618] <=  8'h73;        memory[619] <=  8'h67;        memory[620] <=  8'h79;        memory[621] <=  8'h68;        memory[622] <=  8'h75;        memory[623] <=  8'h61;        memory[624] <=  8'h6a;        memory[625] <=  8'h6b;        memory[626] <=  8'h78;        memory[627] <=  8'h62;        memory[628] <=  8'h20;        memory[629] <=  8'h6e;        memory[630] <=  8'h76;        memory[631] <=  8'h63;        memory[632] <=  8'h61;        memory[633] <=  8'h73;        memory[634] <=  8'h67;        memory[635] <=  8'h68;        memory[636] <=  8'h75;        memory[637] <=  8'h6a;        memory[638] <=  8'h6c;        memory[639] <=  8'h6b;        memory[640] <=  8'h63;        memory[641] <=  8'h78;        memory[642] <=  8'h20;        memory[643] <=  8'h6a;        memory[644] <=  8'h6b;        memory[645] <=  8'h68;        memory[646] <=  8'h61;        memory[647] <=  8'h73;        memory[648] <=  8'h76;        memory[649] <=  8'h64;        memory[650] <=  8'h6e;        memory[651] <=  8'h20;        memory[652] <=  8'h62;        memory[653] <=  8'h6e;        memory[654] <=  8'h6d;        memory[655] <=  8'h6b;        memory[656] <=  8'h77;        memory[657] <=  8'h64;        memory[658] <=  8'h6f;        memory[659] <=  8'h77;        memory[660] <=  8'h69;        memory[661] <=  8'h6f;        memory[662] <=  8'h75;        memory[663] <=  8'h69;        memory[664] <=  8'h68;        memory[665] <=  8'h62;        memory[666] <=  8'h6e;        memory[667] <=  8'h6b;        memory[668] <=  8'h77;        memory[669] <=  8'h69;        memory[670] <=  8'h6f;        memory[671] <=  8'h75;        memory[672] <=  8'h71;        memory[673] <=  8'h69;        memory[674] <=  8'h79;        memory[675] <=  8'h67;        memory[676] <=  8'h6a;        memory[677] <=  8'h64;        memory[678] <=  8'h61;        memory[679] <=  8'h76;        memory[680] <=  8'h62;        memory[681] <=  8'h6e;        memory[682] <=  8'h6b;        memory[683] <=  8'h6f;        memory[684] <=  8'h70;        memory[685] <=  8'h64;        memory[686] <=  8'h76;        memory[687] <=  8'h69;        memory[688] <=  8'h6f;        memory[689] <=  8'h75;        memory[690] <=  8'h69;        memory[691] <=  8'h48;        memory[692] <=  8'h42;        memory[693] <=  8'h6b;        memory[694] <=  8'h64;        memory[695] <=  8'h6e;        memory[696] <=  8'h6c;        memory[697] <=  8'h71;        memory[698] <=  8'h6b;        memory[699] <=  8'h6d;        memory[700] <=  8'h6a;        memory[701] <=  8'h70;        memory[702] <=  8'h69;        memory[703] <=  8'h6f;        memory[704] <=  8'h68;        memory[705] <=  8'h65;        memory[706] <=  8'h66;        memory[707] <=  8'h75;        memory[708] <=  8'h67;        memory[709] <=  8'h69;        memory[710] <=  8'h73;        memory[711] <=  8'h61;        memory[712] <=  8'h62;        memory[713] <=  8'h64;        memory[714] <=  8'h6b;        memory[715] <=  8'h6a;        memory[716] <=  8'h6b;        memory[717] <=  8'h6c;        memory[718] <=  8'h6a;        memory[719] <=  8'h69;        memory[720] <=  8'h73;        memory[721] <=  8'h6f;        memory[722] <=  8'h71;        memory[723] <=  8'h68;        memory[724] <=  8'h77;        memory[725] <=  8'h67;        memory[726] <=  8'h69;        memory[727] <=  8'h79;        memory[728] <=  8'h6a;        memory[729] <=  8'h64;        memory[730] <=  8'h76;        memory[731] <=  8'h62;        memory[732] <=  8'h6e;        memory[733] <=  8'h61;        memory[734] <=  8'h73;        memory[735] <=  8'h66;        memory[736] <=  8'h6c;        memory[737] <=  8'h6b;        memory[738] <=  8'h64;        memory[739] <=  8'h6a;        memory[740] <=  8'h68;        memory[741] <=  8'h63;        memory[742] <=  8'h67;        memory[743] <=  8'h6a;        memory[744] <=  8'h76;        memory[745] <=  8'h73;        memory[746] <=  8'h64;        memory[747] <=  8'h62;        memory[748] <=  8'h62;        memory[749] <=  8'h61;        memory[750] <=  8'h72;        memory[751] <=  8'h62;        memory[752] <=  8'h62;        memory[753] <=  8'h73;        memory[754] <=  8'h62;        memory[755] <=  8'h67;        memory[756] <=  8'h73;        memory[757] <=  8'h66;        memory[758] <=  8'h67;        memory[759] <=  8'h61;        memory[760] <=  8'h68;        memory[761] <=  8'h66;        memory[762] <=  8'h73;        memory[763] <=  8'h68;        memory[764] <=  8'h61;        memory[765] <=  8'h66;        memory[766] <=  8'h73;        memory[767] <=  8'h66;        memory[768] <=  8'h68;        memory[769] <=  8'h61;        memory[770] <=  8'h69;        memory[771] <=  8'h64;        memory[772] <=  8'h75;        memory[773] <=  8'h67;        memory[774] <=  8'h64;        memory[775] <=  8'h77;        memory[776] <=  8'h62;        memory[777] <=  8'h61;        memory[778] <=  8'h62;        memory[779] <=  8'h72;        memory[780] <=  8'h62;        memory[781] <=  8'h61;        memory[782] <=  8'h62;        memory[783] <=  8'h62;        memory[784] <=  8'h74;        memory[785] <=  8'h62;        memory[786] <=  8'h62;        memory[787] <=  8'h62;        memory[788] <=  8'h62;        memory[789] <=  8'h62;        memory[790] <=  8'h62;        memory[791] <=  8'h62;        memory[792] <=  8'h62;        memory[793] <=  8'h61;        memory[794] <=  8'h62;        memory[795] <=  8'h62;        memory[796] <=  8'h72;        memory[797] <=  8'h74;        memory[798] <=  8'h62;        memory[799] <=  8'h62;        memory[800] <=  8'h61;        memory[801] <=  8'h62;        memory[802] <=  8'h72;        memory[803] <=  8'h62;        memory[804] <=  8'h74;        memory[805] <=  8'h62;        memory[806] <=  8'h62;        memory[807] <=  8'h62;        memory[808] <=  8'h63;        memory[809] <=  8'h61;        memory[810] <=  8'h72;        memory[811] <=  8'h74;        memory[812] <=  8'h73;        memory[813] <=  8'h62;        memory[814] <=  8'h61;        memory[815] <=  8'h72;        memory[816] <=  8'h74;        memory[817] <=  8'h74;        memory[818] <=  8'h62;        memory[819] <=  8'h61;        memory[820] <=  8'h72;        memory[821] <=  8'h74;        memory[822] <=  8'h78;        memory[823] <=  8'h61;        memory[824] <=  8'h74;        memory[825] <=  8'h6b;        memory[826] <=  8'h73;        memory[827] <=  8'h68;        memory[828] <=  8'h63;        memory[829] <=  8'h66;        memory[830] <=  8'h69;        memory[831] <=  8'h77;        memory[832] <=  8'h68;        memory[833] <=  8'h61;        memory[834] <=  8'h74;        memory[835] <=  8'h61;        memory[836] <=  8'h6e;        memory[837] <=  8'h61;        memory[838] <=  8'h62;        memory[839] <=  8'h61;        memory[840] <=  8'h63;        memory[841] <=  8'h61;        memory[842] <=  8'h74;        memory[843] <=  8'h61;        memory[844] <=  8'h62;        memory[845] <=  8'h61;        memory[846] <=  8'h72;        memory[847] <=  8'h63;        memory[848] <=  8'h61;        memory[849] <=  8'h68;        memory[850] <=  8'h64;        memory[851] <=  8'h75;        memory[852] <=  8'h63;        memory[853] <=  8'h74;        memory[854] <=  8'h61;        memory[855] <=  8'h64;        memory[856] <=  8'h61;        memory[857] <=  8'h61;        memory[858] <=  8'h63;        memory[859] <=  8'h61;        memory[860] <=  8'h72;        memory[861] <=  8'h63;        memory[862] <=  8'h74;        memory[863] <=  8'h72;        memory[864] <=  8'h63;        memory[865] <=  8'h61;        memory[866] <=  8'h74;        memory[867] <=  8'h72;        memory[868] <=  8'h63;        memory[869] <=  8'h61;        memory[870] <=  8'h74;        memory[871] <=  8'h63;        memory[872] <=  8'h62;        memory[873] <=  8'h61;        memory[874] <=  8'h74;        memory[875] <=  8'h62;        memory[876] <=  8'h72;        memory[877] <=  8'h63;        memory[878] <=  8'h61;        memory[879] <=  8'h74;        memory[880] <=  8'h72;        memory[881] <=  8'h6e;        memory[882] <=  8'h62;        memory[883] <=  8'h61;        memory[884] <=  8'h63;        memory[885] <=  8'h61;        memory[886] <=  8'h74;        memory[887] <=  8'h79;        memory[888] <=  8'h73;        memory[889] <=  8'h6e;        memory[890] <=  8'h63;        memory[891] <=  8'h74;        memory[892] <=  8'h61;        memory[893] <=  8'h6e;        memory[894] <=  8'h62;        memory[895] <=  8'h61;        memory[896] <=  8'h63;        memory[897] <=  8'h72;        memory[898] <=  8'h6e;        memory[899] <=  8'h74;        memory[900] <=  8'h61;        memory[901] <=  8'h62;        memory[902] <=  8'h74;        memory[903] <=  8'h6e;        memory[904] <=  8'h61;        memory[905] <=  8'h72;        memory[906] <=  8'h62;        memory[907] <=  8'h78;        memory[908] <=  8'h74;        memory[909] <=  8'h61;        memory[910] <=  8'h72;        memory[911] <=  8'h62;        memory[912] <=  8'h61;        memory[913] <=  8'h72;        memory[914] <=  8'h74;        memory[915] <=  8'h74;        memory[916] <=  8'h62;        memory[917] <=  8'h61;        memory[918] <=  8'h72;        memory[919] <=  8'h74;        memory[920] <=  8'h78;        memory[921] <=  8'h61;        memory[922] <=  8'h74;        memory[923] <=  8'h6b;        memory[924] <=  8'h73;        memory[925] <=  8'h68;        memory[926] <=  8'h63;        memory[927] <=  8'h66;        memory[928] <=  8'h69;        memory[929] <=  8'h77;        memory[930] <=  8'h68;        memory[931] <=  8'h61;        memory[932] <=  8'h74;        memory[933] <=  8'h61;        memory[934] <=  8'h6e;        memory[935] <=  8'h61;        memory[936] <=  8'h62;        memory[937] <=  8'h61;        memory[938] <=  8'h63;        memory[939] <=  8'h61;        memory[940] <=  8'h74;        memory[941] <=  8'h61;        memory[942] <=  8'h62;        memory[943] <=  8'h61;        memory[944] <=  8'h72;        memory[945] <=  8'h63;        memory[946] <=  8'h61;        memory[947] <=  8'h68;        memory[948] <=  8'h64;        memory[949] <=  8'h75;        memory[950] <=  8'h63;        memory[951] <=  8'h74;        memory[952] <=  8'h61;        memory[953] <=  8'h64;        memory[954] <=  8'h61;        memory[955] <=  8'h61;        memory[956] <=  8'h63;        memory[957] <=  8'h61;        memory[958] <=  8'h72;        memory[959] <=  8'h63;        memory[960] <=  8'h74;        memory[961] <=  8'h72;        memory[962] <=  8'h63;        memory[963] <=  8'h61;        memory[964] <=  8'h74;        memory[965] <=  8'h72;        memory[966] <=  8'h63;        memory[967] <=  8'h61;        memory[968] <=  8'h74;        memory[969] <=  8'h63;        memory[970] <=  8'h62;        memory[971] <=  8'h61;        memory[972] <=  8'h74;        memory[973] <=  8'h62;        memory[974] <=  8'h72;        memory[975] <=  8'h63;        memory[976] <=  8'h61;        memory[977] <=  8'h74;        memory[978] <=  8'h72;        memory[979] <=  8'h6e;        memory[980] <=  8'h62;        memory[981] <=  8'h61;        memory[982] <=  8'h63;        memory[983] <=  8'h61;        memory[984] <=  8'h74;        memory[985] <=  8'h79;        memory[986] <=  8'h73;        memory[987] <=  8'h6e;        memory[988] <=  8'h63;        memory[989] <=  8'h74;        memory[990] <=  8'h61;        memory[991] <=  8'h6e;        memory[992] <=  8'h62;        memory[993] <=  8'h61;        memory[994] <=  8'h63;        memory[995] <=  8'h72;        memory[996] <=  8'h6e;        memory[997] <=  8'h74;        memory[998] <=  8'h61;        memory[999] <=  8'h62;        memory[1000] <=  8'h74;        memory[1001] <=  8'h6e;        memory[1002] <=  8'h61;        memory[1003] <=  8'h72;        memory[1004] <=  8'h62;        memory[1005] <=  8'h78;        memory[1006] <=  8'h74;        memory[1007] <=  8'h61;        memory[1008] <=  8'h72;        memory[1009] <=  8'h62;        memory[1010] <=  8'h61;        memory[1011] <=  8'h72;        memory[1012] <=  8'h74;        memory[1013] <=  8'h74;        memory[1014] <=  8'h62;        memory[1015] <=  8'h61;        memory[1016] <=  8'h72;        memory[1017] <=  8'h74;        memory[1018] <=  8'h78;        memory[1019] <=  8'h61;        memory[1020] <=  8'h74;        memory[1021] <=  8'h6b;        memory[1022] <=  8'h73;        memory[1023] <=  8'h68;        memory[1024] <=  8'h63;        memory[1025] <=  8'h66;        memory[1026] <=  8'h69;        memory[1027] <=  8'h77;        memory[1028] <=  8'h68;        memory[1029] <=  8'h61;        memory[1030] <=  8'h74;        memory[1031] <=  8'h61;        memory[1032] <=  8'h6e;        memory[1033] <=  8'h61;        memory[1034] <=  8'h62;        memory[1035] <=  8'h61;        memory[1036] <=  8'h63;        memory[1037] <=  8'h61;        memory[1038] <=  8'h74;        memory[1039] <=  8'h61;        memory[1040] <=  8'h62;        memory[1041] <=  8'h61;        memory[1042] <=  8'h72;        memory[1043] <=  8'h63;        memory[1044] <=  8'h61;        memory[1045] <=  8'h68;        memory[1046] <=  8'h64;        memory[1047] <=  8'h75;        memory[1048] <=  8'h63;        memory[1049] <=  8'h74;        memory[1050] <=  8'h61;        memory[1051] <=  8'h64;        memory[1052] <=  8'h61;        memory[1053] <=  8'h61;        memory[1054] <=  8'h63;        memory[1055] <=  8'h61;        memory[1056] <=  8'h72;        memory[1057] <=  8'h63;        memory[1058] <=  8'h74;        memory[1059] <=  8'h72;        memory[1060] <=  8'h63;        memory[1061] <=  8'h61;        memory[1062] <=  8'h74;        memory[1063] <=  8'h72;        memory[1064] <=  8'h63;        memory[1065] <=  8'h61;        memory[1066] <=  8'h74;        memory[1067] <=  8'h63;        memory[1068] <=  8'h62;        memory[1069] <=  8'h61;        memory[1070] <=  8'h74;        memory[1071] <=  8'h62;        memory[1072] <=  8'h72;        memory[1073] <=  8'h63;        memory[1074] <=  8'h61;        memory[1075] <=  8'h74;        memory[1076] <=  8'h72;        memory[1077] <=  8'h6e;        memory[1078] <=  8'h62;        memory[1079] <=  8'h61;        memory[1080] <=  8'h63;        memory[1081] <=  8'h61;        memory[1082] <=  8'h74;        memory[1083] <=  8'h79;        memory[1084] <=  8'h73;        memory[1085] <=  8'h6e;        memory[1086] <=  8'h63;        memory[1087] <=  8'h74;        memory[1088] <=  8'h61;        memory[1089] <=  8'h6e;        memory[1090] <=  8'h62;        memory[1091] <=  8'h61;        memory[1092] <=  8'h63;        memory[1093] <=  8'h72;        memory[1094] <=  8'h6e;        memory[1095] <=  8'h74;        memory[1096] <=  8'h61;        memory[1097] <=  8'h62;        memory[1098] <=  8'h74;        memory[1099] <=  8'h6e;        memory[1100] <=  8'h61;        memory[1101] <=  8'h72;        memory[1102] <=  8'h62;        memory[1103] <=  8'h78;        memory[1104] <=  8'h74;        memory[1105] <=  8'h61;        memory[1106] <=  8'h72;        memory[1107] <=  8'h5d;        memory[1108] <=  8'h5d;        memory[1109] <=  8'h65;        memory[1110] <=  8'h66;        memory[1111] <=  8'h77;        memory[1112] <=  8'h65;        memory[1113] <=  8'h5d;        memory[1114] <=  8'h65;        memory[1115] <=  8'h67;        memory[1116] <=  8'h73;        memory[1117] <=  8'h67;        memory[1118] <=  8'h66;        memory[1119] <=  8'h62;        memory[1120] <=  8'h61;        memory[1121] <=  8'h72;        memory[1122] <=  8'h74;        memory[1123] <=  8'h74;        memory[1124] <=  8'h62;        memory[1125] <=  8'h61;        memory[1126] <=  8'h72;        memory[1127] <=  8'h74;        memory[1128] <=  8'h78;        memory[1129] <=  8'h61;        memory[1130] <=  8'h74;        memory[1131] <=  8'h6b;        memory[1132] <=  8'h73;        memory[1133] <=  8'h68;        memory[1134] <=  8'h63;        memory[1135] <=  8'h66;        memory[1136] <=  8'h69;        memory[1137] <=  8'h77;        memory[1138] <=  8'h68;        memory[1139] <=  8'h61;        memory[1140] <=  8'h74;        memory[1141] <=  8'h61;        memory[1142] <=  8'h6e;        memory[1143] <=  8'h61;        memory[1144] <=  8'h62;        memory[1145] <=  8'h61;        memory[1146] <=  8'h63;        memory[1147] <=  8'h61;        memory[1148] <=  8'h74;        memory[1149] <=  8'h61;        memory[1150] <=  8'h62;        memory[1151] <=  8'h61;        memory[1152] <=  8'h72;        memory[1153] <=  8'h63;        memory[1154] <=  8'h61;        memory[1155] <=  8'h68;        memory[1156] <=  8'h64;        memory[1157] <=  8'h75;        memory[1158] <=  8'h63;        memory[1159] <=  8'h74;        memory[1160] <=  8'h61;        memory[1161] <=  8'h64;        memory[1162] <=  8'h61;        memory[1163] <=  8'h61;        memory[1164] <=  8'h63;        memory[1165] <=  8'h61;        memory[1166] <=  8'h72;        memory[1167] <=  8'h63;        memory[1168] <=  8'h74;        memory[1169] <=  8'h72;        memory[1170] <=  8'h63;        memory[1171] <=  8'h61;        memory[1172] <=  8'h74;        memory[1173] <=  8'h72;        memory[1174] <=  8'h63;        memory[1175] <=  8'h61;        memory[1176] <=  8'h74;        memory[1177] <=  8'h63;        memory[1178] <=  8'h62;        memory[1179] <=  8'h61;        memory[1180] <=  8'h74;        memory[1181] <=  8'h62;        memory[1182] <=  8'h72;        memory[1183] <=  8'h63;        memory[1184] <=  8'h61;        memory[1185] <=  8'h74;        memory[1186] <=  8'h72;        memory[1187] <=  8'h6e;        memory[1188] <=  8'h62;        memory[1189] <=  8'h61;        memory[1190] <=  8'h63;        memory[1191] <=  8'h61;        memory[1192] <=  8'h74;        memory[1193] <=  8'h79;        memory[1194] <=  8'h73;        memory[1195] <=  8'h6e;        memory[1196] <=  8'h63;        memory[1197] <=  8'h74;        memory[1198] <=  8'h61;        memory[1199] <=  8'h6e;        memory[1200] <=  8'h62;        memory[1201] <=  8'h61;        memory[1202] <=  8'h63;        memory[1203] <=  8'h72;        memory[1204] <=  8'h6e;        memory[1205] <=  8'h74;        memory[1206] <=  8'h61;        memory[1207] <=  8'h62;        memory[1208] <=  8'h74;        memory[1209] <=  8'h6e;        memory[1210] <=  8'h61;        memory[1211] <=  8'h72;        memory[1212] <=  8'h62;        memory[1213] <=  8'h78;        memory[1214] <=  8'h74;        memory[1215] <=  8'h61;        memory[1216] <=  8'h72;        memory[1217] <=  8'h62;        memory[1218] <=  8'h61;        memory[1219] <=  8'h72;        memory[1220] <=  8'h74;        memory[1221] <=  8'h74;        memory[1222] <=  8'h62;        memory[1223] <=  8'h61;        memory[1224] <=  8'h72;        memory[1225] <=  8'h74;        memory[1226] <=  8'h78;        memory[1227] <=  8'h61;        memory[1228] <=  8'h74;        memory[1229] <=  8'h6b;        memory[1230] <=  8'h73;        memory[1231] <=  8'h68;        memory[1232] <=  8'h63;        memory[1233] <=  8'h66;        memory[1234] <=  8'h69;        memory[1235] <=  8'h77;        memory[1236] <=  8'h68;        memory[1237] <=  8'h61;        memory[1238] <=  8'h74;        memory[1239] <=  8'h61;        memory[1240] <=  8'h6e;        memory[1241] <=  8'h61;        memory[1242] <=  8'h62;        memory[1243] <=  8'h61;        memory[1244] <=  8'h63;        memory[1245] <=  8'h61;        memory[1246] <=  8'h74;        memory[1247] <=  8'h61;        memory[1248] <=  8'h62;        memory[1249] <=  8'h61;        memory[1250] <=  8'h72;        memory[1251] <=  8'h63;        memory[1252] <=  8'h61;        memory[1253] <=  8'h68;        memory[1254] <=  8'h64;        memory[1255] <=  8'h75;        memory[1256] <=  8'h63;        memory[1257] <=  8'h74;        memory[1258] <=  8'h61;        memory[1259] <=  8'h64;        memory[1260] <=  8'h61;        memory[1261] <=  8'h61;        memory[1262] <=  8'h63;        memory[1263] <=  8'h61;        memory[1264] <=  8'h72;        memory[1265] <=  8'h63;        memory[1266] <=  8'h74;        memory[1267] <=  8'h72;        memory[1268] <=  8'h63;        memory[1269] <=  8'h61;        memory[1270] <=  8'h74;        memory[1271] <=  8'h72;        memory[1272] <=  8'h63;        memory[1273] <=  8'h61;        memory[1274] <=  8'h74;        memory[1275] <=  8'h63;        memory[1276] <=  8'h62;        memory[1277] <=  8'h61;        memory[1278] <=  8'h71;        memory[1279] <=  8'h74;        memory[1280] <=  8'h74;        memory[1281] <=  8'h62;        memory[1282] <=  8'h72;        memory[1283] <=  8'h63;        memory[1284] <=  8'h61;        memory[1285] <=  8'h74;        memory[1286] <=  8'h72;        memory[1287] <=  8'h6e;        memory[1288] <=  8'h62;        memory[1289] <=  8'h61;        memory[1290] <=  8'h63;        memory[1291] <=  8'h61;        memory[1292] <=  8'h74;        memory[1293] <=  8'h79;        memory[1294] <=  8'h73;        memory[1295] <=  8'h6e;        memory[1296] <=  8'h63;        memory[1297] <=  8'h74;        memory[1298] <=  8'h61;        memory[1299] <=  8'h6e;        memory[1300] <=  8'h62;        memory[1301] <=  8'h61;        memory[1302] <=  8'h63;        memory[1303] <=  8'h72;        memory[1304] <=  8'h6e;        memory[1305] <=  8'h74;        memory[1306] <=  8'h61;        memory[1307] <=  8'h62;        memory[1308] <=  8'h74;        memory[1309] <=  8'h6e;        memory[1310] <=  8'h61;        memory[1311] <=  8'h72;        memory[1312] <=  8'h62;        memory[1313] <=  8'h78;        memory[1314] <=  8'h74;        memory[1315] <=  8'h61;        memory[1316] <=  8'h72;        memory[1317] <=  8'h64;        memory[1318] <=  8'h66;        memory[1319] <=  8'h73;        memory[1320] <=  8'h67;        memory[1321] <=  8'h76;        memory[1322] <=  8'h68;        memory[1323] <=  8'h62;        memory[1324] <=  8'h6b;        memory[1325] <=  8'h6a;        memory[1326] <=  8'h6e;        memory[1327] <=  8'h6d;        memory[1328] <=  8'h62;        memory[1329] <=  8'h76;        memory[1330] <=  8'h78;        memory[1331] <=  8'h63;        memory[1332] <=  8'h73;        memory[1333] <=  8'h66;        memory[1334] <=  8'h72;        memory[1335] <=  8'h74;        memory[1336] <=  8'h79;        memory[1337] <=  8'h75;        memory[1338] <=  8'h6a;        memory[1339] <=  8'h6e;        memory[1340] <=  8'h62;        memory[1341] <=  8'h76;        memory[1342] <=  8'h63;        memory[1343] <=  8'h64;        memory[1344] <=  8'h74;        memory[1345] <=  8'h79;        memory[1346] <=  8'h75;        memory[1347] <=  8'h69;        memory[1348] <=  8'h6b;        memory[1349] <=  8'h6d;        memory[1350] <=  8'h6e;        memory[1351] <=  8'h62;        memory[1352] <=  8'h76;        memory[1353] <=  8'h63;        memory[1354] <=  8'h78;        memory[1355] <=  8'h73;        memory[1356] <=  8'h64;        memory[1357] <=  8'h72;        memory[1358] <=  8'h74;        memory[1359] <=  8'h79;        memory[1360] <=  8'h75;        memory[1361] <=  8'h69;        memory[1362] <=  8'h6b;        memory[1363] <=  8'h6d;        memory[1364] <=  8'h6e;        memory[1365] <=  8'h62;        memory[1366] <=  8'h76;        memory[1367] <=  8'h63;        memory[1368] <=  8'h73;        memory[1369] <=  8'h77;        memory[1370] <=  8'h33;        memory[1371] <=  8'h34;        memory[1372] <=  8'h35;        memory[1373] <=  8'h36;        memory[1374] <=  8'h37;        memory[1375] <=  8'h38;        memory[1376] <=  8'h69;        memory[1377] <=  8'h6b;        memory[1378] <=  8'h6d;        memory[1379] <=  8'h6e;        memory[1380] <=  8'h62;        memory[1381] <=  8'h76;        memory[1382] <=  8'h63;        memory[1383] <=  8'h64;        memory[1384] <=  8'h65;        memory[1385] <=  8'h72;        memory[1386] <=  8'h36;        memory[1387] <=  8'h37;        memory[1388] <=  8'h38;        memory[1389] <=  8'h69;        memory[1390] <=  8'h6f;        memory[1391] <=  8'h6b;        memory[1392] <=  8'h6a;        memory[1393] <=  8'h6e;        memory[1394] <=  8'h62;        memory[1395] <=  8'h76;        memory[1396] <=  8'h63;        memory[1397] <=  8'h64;        memory[1398] <=  8'h72;        memory[1399] <=  8'h74;        memory[1400] <=  8'h79;        memory[1401] <=  8'h75;        memory[1402] <=  8'h73;        memory[1403] <=  8'h6a;        memory[1404] <=  8'h63;        memory[1405] <=  8'h6e;        memory[1406] <=  8'h62;        memory[1407] <=  8'h64;        memory[1408] <=  8'h66;        memory[1409] <=  8'h73;        memory[1410] <=  8'h74;        memory[1411] <=  8'h79;        memory[1412] <=  8'h75;        memory[1413] <=  8'h61;        memory[1414] <=  8'h69;        memory[1415] <=  8'h6b;        memory[1416] <=  8'h78;        memory[1417] <=  8'h6d;        memory[1418] <=  8'h6e;        memory[1419] <=  8'h73;        memory[1420] <=  8'h6a;        memory[1421] <=  8'h6f;        memory[1422] <=  8'h64;        memory[1423] <=  8'h6c;        memory[1424] <=  8'h63;        memory[1425] <=  8'h78;        memory[1426] <=  8'h62;        memory[1427] <=  8'h61;        memory[1428] <=  8'h72;        memory[1429] <=  8'h74;        memory[1430] <=  8'h78;        memory[1431] <=  8'h61;        memory[1432] <=  8'h74;        memory[1433] <=  8'h6b;        memory[1434] <=  8'h73;        memory[1435] <=  8'h68;        memory[1436] <=  8'h63;        memory[1437] <=  8'h66;        memory[1438] <=  8'h69;        memory[1439] <=  8'h77;        memory[1440] <=  8'h68;        memory[1441] <=  8'h61;        memory[1442] <=  8'h74;        memory[1443] <=  8'h61;        memory[1444] <=  8'h6e;        memory[1445] <=  8'h61;        memory[1446] <=  8'h62;        memory[1447] <=  8'h61;        memory[1448] <=  8'h63;        memory[1449] <=  8'h61;        memory[1450] <=  8'h74;        memory[1451] <=  8'h61;        memory[1452] <=  8'h62;        memory[1453] <=  8'h61;        memory[1454] <=  8'h72;        memory[1455] <=  8'h63;        memory[1456] <=  8'h61;        memory[1457] <=  8'h68;        memory[1458] <=  8'h64;        memory[1459] <=  8'h75;        memory[1460] <=  8'h63;        memory[1461] <=  8'h74;        memory[1462] <=  8'h61;        memory[1463] <=  8'h64;        memory[1464] <=  8'h61;        memory[1465] <=  8'h61;        memory[1466] <=  8'h63;        memory[1467] <=  8'h61;        memory[1468] <=  8'h72;        memory[1469] <=  8'h62;        memory[1470] <=  8'h61;        memory[1471] <=  8'h72;        memory[1472] <=  8'h74;        memory[1473] <=  8'h78;        memory[1474] <=  8'h61;        memory[1475] <=  8'h74;        memory[1476] <=  8'h6b;        memory[1477] <=  8'h73;        memory[1478] <=  8'h68;        memory[1479] <=  8'h63;        memory[1480] <=  8'h66;        memory[1481] <=  8'h69;        memory[1482] <=  8'h77;        memory[1483] <=  8'h68;        memory[1484] <=  8'h61;        memory[1485] <=  8'h74;        memory[1486] <=  8'h61;        memory[1487] <=  8'h6e;        memory[1488] <=  8'h61;        memory[1489] <=  8'h62;        memory[1490] <=  8'h61;        memory[1491] <=  8'h63;        memory[1492] <=  8'h61;        memory[1493] <=  8'h74;        memory[1494] <=  8'h61;        memory[1495] <=  8'h62;        memory[1496] <=  8'h61;        memory[1497] <=  8'h72;        memory[1498] <=  8'h63;        memory[1499] <=  8'h61;        memory[1500] <=  8'h68;        memory[1501] <=  8'h64;        memory[1502] <=  8'h75;        memory[1503] <=  8'h63;        memory[1504] <=  8'h74;        memory[1505] <=  8'h61;        memory[1506] <=  8'h64;        memory[1507] <=  8'h61;        memory[1508] <=  8'h61;        memory[1509] <=  8'h63;        memory[1510] <=  8'h61;        memory[1511] <=  8'h72;        memory[1512] <=  8'h62;        memory[1513] <=  8'h61;        memory[1514] <=  8'h72;        memory[1515] <=  8'h74;        memory[1516] <=  8'h78;        memory[1517] <=  8'h61;        memory[1518] <=  8'h74;        memory[1519] <=  8'h6b;        memory[1520] <=  8'h73;        memory[1521] <=  8'h68;        memory[1522] <=  8'h63;        memory[1523] <=  8'h66;        memory[1524] <=  8'h69;        memory[1525] <=  8'h77;        memory[1526] <=  8'h68;        memory[1527] <=  8'h61;        memory[1528] <=  8'h74;        memory[1529] <=  8'h61;        memory[1530] <=  8'h6e;        memory[1531] <=  8'h61;        memory[1532] <=  8'h62;        memory[1533] <=  8'h61;        memory[1534] <=  8'h63;        memory[1535] <=  8'h61;        memory[1536] <=  8'h74;        memory[1537] <=  8'h61;        memory[1538] <=  8'h62;        memory[1539] <=  8'h61;        memory[1540] <=  8'h72;        memory[1541] <=  8'h63;        memory[1542] <=  8'h61;        memory[1543] <=  8'h68;        memory[1544] <=  8'h64;        memory[1545] <=  8'h75;        memory[1546] <=  8'h63;        memory[1547] <=  8'h74;        memory[1548] <=  8'h61;        memory[1549] <=  8'h64;        memory[1550] <=  8'h61;        memory[1551] <=  8'h61;        memory[1552] <=  8'h63;        memory[1553] <=  8'h61;        memory[1554] <=  8'h72;        memory[1555] <=  8'h62;        memory[1556] <=  8'h61;        memory[1557] <=  8'h72;        memory[1558] <=  8'h74;        memory[1559] <=  8'h78;        memory[1560] <=  8'h61;        memory[1561] <=  8'h74;        memory[1562] <=  8'h6b;        memory[1563] <=  8'h73;        memory[1564] <=  8'h68;        memory[1565] <=  8'h63;        memory[1566] <=  8'h66;        memory[1567] <=  8'h69;        memory[1568] <=  8'h77;        memory[1569] <=  8'h68;        memory[1570] <=  8'h61;        memory[1571] <=  8'h74;        memory[1572] <=  8'h61;        memory[1573] <=  8'h6e;        memory[1574] <=  8'h61;        memory[1575] <=  8'h62;        memory[1576] <=  8'h61;        memory[1577] <=  8'h63;        memory[1578] <=  8'h61;        memory[1579] <=  8'h74;        memory[1580] <=  8'h61;        memory[1581] <=  8'h62;        memory[1582] <=  8'h61;        memory[1583] <=  8'h72;        memory[1584] <=  8'h63;        memory[1585] <=  8'h61;        memory[1586] <=  8'h68;        memory[1587] <=  8'h64;        memory[1588] <=  8'h75;        memory[1589] <=  8'h63;        memory[1590] <=  8'h74;        memory[1591] <=  8'h61;        memory[1592] <=  8'h64;        memory[1593] <=  8'h61;        memory[1594] <=  8'h61;        memory[1595] <=  8'h63;        memory[1596] <=  8'h61;        memory[1597] <=  8'h72;        memory[1598] <=  8'h62;        memory[1599] <=  8'h61;        memory[1600] <=  8'h72;        memory[1601] <=  8'h74;        memory[1602] <=  8'h78;        memory[1603] <=  8'h61;        memory[1604] <=  8'h74;        memory[1605] <=  8'h6b;        memory[1606] <=  8'h73;        memory[1607] <=  8'h68;        memory[1608] <=  8'h63;        memory[1609] <=  8'h66;        memory[1610] <=  8'h69;        memory[1611] <=  8'h77;        memory[1612] <=  8'h68;        memory[1613] <=  8'h61;        memory[1614] <=  8'h74;        memory[1615] <=  8'h61;        memory[1616] <=  8'h6e;        memory[1617] <=  8'h61;        memory[1618] <=  8'h62;        memory[1619] <=  8'h61;        memory[1620] <=  8'h63;        memory[1621] <=  8'h61;        memory[1622] <=  8'h74;        memory[1623] <=  8'h61;        memory[1624] <=  8'h62;        memory[1625] <=  8'h61;        memory[1626] <=  8'h72;        memory[1627] <=  8'h63;        memory[1628] <=  8'h61;        memory[1629] <=  8'h68;        memory[1630] <=  8'h64;        memory[1631] <=  8'h75;        memory[1632] <=  8'h63;        memory[1633] <=  8'h74;        memory[1634] <=  8'h61;        memory[1635] <=  8'h64;        memory[1636] <=  8'h61;        memory[1637] <=  8'h61;        memory[1638] <=  8'h63;        memory[1639] <=  8'h61;        memory[1640] <=  8'h72;        memory[1641] <=  8'h62;        memory[1642] <=  8'h61;        memory[1643] <=  8'h72;        memory[1644] <=  8'h74;        memory[1645] <=  8'h78;        memory[1646] <=  8'h61;        memory[1647] <=  8'h74;        memory[1648] <=  8'h6b;        memory[1649] <=  8'h73;        memory[1650] <=  8'h68;        memory[1651] <=  8'h63;        memory[1652] <=  8'h66;        memory[1653] <=  8'h69;        memory[1654] <=  8'h77;        memory[1655] <=  8'h68;        memory[1656] <=  8'h61;        memory[1657] <=  8'h74;        memory[1658] <=  8'h61;        memory[1659] <=  8'h6e;        memory[1660] <=  8'h61;        memory[1661] <=  8'h62;        memory[1662] <=  8'h61;        memory[1663] <=  8'h63;        memory[1664] <=  8'h61;        memory[1665] <=  8'h74;        memory[1666] <=  8'h61;        memory[1667] <=  8'h62;        memory[1668] <=  8'h61;        memory[1669] <=  8'h72;        memory[1670] <=  8'h63;        memory[1671] <=  8'h61;        memory[1672] <=  8'h68;        memory[1673] <=  8'h64;        memory[1674] <=  8'h75;        memory[1675] <=  8'h63;        memory[1676] <=  8'h74;        memory[1677] <=  8'h61;        memory[1678] <=  8'h64;        memory[1679] <=  8'h61;        memory[1680] <=  8'h61;        memory[1681] <=  8'h63;        memory[1682] <=  8'h61;        memory[1683] <=  8'h72;        memory[1684] <=  8'h62;        memory[1685] <=  8'h61;        memory[1686] <=  8'h72;        memory[1687] <=  8'h74;        memory[1688] <=  8'h78;        memory[1689] <=  8'h61;        memory[1690] <=  8'h74;        memory[1691] <=  8'h6b;        memory[1692] <=  8'h73;        memory[1693] <=  8'h68;        memory[1694] <=  8'h63;        memory[1695] <=  8'h66;        memory[1696] <=  8'h69;        memory[1697] <=  8'h77;        memory[1698] <=  8'h68;        memory[1699] <=  8'h61;        memory[1700] <=  8'h74;        memory[1701] <=  8'h61;        memory[1702] <=  8'h6e;        memory[1703] <=  8'h61;        memory[1704] <=  8'h62;        memory[1705] <=  8'h61;        memory[1706] <=  8'h63;        memory[1707] <=  8'h61;        memory[1708] <=  8'h74;        memory[1709] <=  8'h61;        memory[1710] <=  8'h62;        memory[1711] <=  8'h61;        memory[1712] <=  8'h72;        memory[1713] <=  8'h63;        memory[1714] <=  8'h61;        memory[1715] <=  8'h68;        memory[1716] <=  8'h64;        memory[1717] <=  8'h75;        memory[1718] <=  8'h63;        memory[1719] <=  8'h74;        memory[1720] <=  8'h61;        memory[1721] <=  8'h64;        memory[1722] <=  8'h61;        memory[1723] <=  8'h61;        memory[1724] <=  8'h63;        memory[1725] <=  8'h61;        memory[1726] <=  8'h72;        memory[1727] <=  8'h62;        memory[1728] <=  8'h61;        memory[1729] <=  8'h72;        memory[1730] <=  8'h74;        memory[1731] <=  8'h78;        memory[1732] <=  8'h61;        memory[1733] <=  8'h74;        memory[1734] <=  8'h6b;        memory[1735] <=  8'h73;        memory[1736] <=  8'h68;        memory[1737] <=  8'h63;        memory[1738] <=  8'h66;        memory[1739] <=  8'h69;        memory[1740] <=  8'h77;        memory[1741] <=  8'h68;        memory[1742] <=  8'h61;        memory[1743] <=  8'h74;        memory[1744] <=  8'h61;        memory[1745] <=  8'h6e;        memory[1746] <=  8'h61;        memory[1747] <=  8'h62;        memory[1748] <=  8'h61;        memory[1749] <=  8'h63;        memory[1750] <=  8'h61;        memory[1751] <=  8'h74;        memory[1752] <=  8'h61;        memory[1753] <=  8'h62;        memory[1754] <=  8'h61;        memory[1755] <=  8'h72;        memory[1756] <=  8'h63;        memory[1757] <=  8'h61;        memory[1758] <=  8'h68;        memory[1759] <=  8'h64;        memory[1760] <=  8'h75;        memory[1761] <=  8'h63;        memory[1762] <=  8'h74;        memory[1763] <=  8'h61;        memory[1764] <=  8'h64;        memory[1765] <=  8'h61;        memory[1766] <=  8'h61;        memory[1767] <=  8'h63;        memory[1768] <=  8'h61;        memory[1769] <=  8'h72;        memory[1770] <=  8'h62;        memory[1771] <=  8'h61;        memory[1772] <=  8'h72;        memory[1773] <=  8'h74;        memory[1774] <=  8'h78;        memory[1775] <=  8'h61;        memory[1776] <=  8'h74;        memory[1777] <=  8'h6b;        memory[1778] <=  8'h73;        memory[1779] <=  8'h68;        memory[1780] <=  8'h63;        memory[1781] <=  8'h66;        memory[1782] <=  8'h69;        memory[1783] <=  8'h77;        memory[1784] <=  8'h68;        memory[1785] <=  8'h61;        memory[1786] <=  8'h74;        memory[1787] <=  8'h61;        memory[1788] <=  8'h6e;        memory[1789] <=  8'h61;        memory[1790] <=  8'h62;        memory[1791] <=  8'h61;        memory[1792] <=  8'h63;        memory[1793] <=  8'h61;        memory[1794] <=  8'h74;        memory[1795] <=  8'h61;        memory[1796] <=  8'h62;        memory[1797] <=  8'h61;        memory[1798] <=  8'h72;        memory[1799] <=  8'h63;        memory[1800] <=  8'h61;        memory[1801] <=  8'h68;        memory[1802] <=  8'h64;        memory[1803] <=  8'h75;        memory[1804] <=  8'h63;        memory[1805] <=  8'h74;        memory[1806] <=  8'h61;        memory[1807] <=  8'h64;        memory[1808] <=  8'h61;        memory[1809] <=  8'h61;        memory[1810] <=  8'h63;        memory[1811] <=  8'h61;        memory[1812] <=  8'h72;        memory[1813] <=  8'h62;        memory[1814] <=  8'h61;        memory[1815] <=  8'h72;        memory[1816] <=  8'h74;        memory[1817] <=  8'h74;        memory[1818] <=  8'h62;        memory[1819] <=  8'h61;        memory[1820] <=  8'h72;        memory[1821] <=  8'h74;        memory[1822] <=  8'h78;        memory[1823] <=  8'h61;        memory[1824] <=  8'h74;        memory[1825] <=  8'h6b;        memory[1826] <=  8'h73;        memory[1827] <=  8'h68;        memory[1828] <=  8'h63;        memory[1829] <=  8'h66;        memory[1830] <=  8'h69;        memory[1831] <=  8'h77;        memory[1832] <=  8'h68;        memory[1833] <=  8'h61;        memory[1834] <=  8'h74;        memory[1835] <=  8'h61;        memory[1836] <=  8'h6e;        memory[1837] <=  8'h61;        memory[1838] <=  8'h62;        memory[1839] <=  8'h61;        memory[1840] <=  8'h63;        memory[1841] <=  8'h61;        memory[1842] <=  8'h74;        memory[1843] <=  8'h61;        memory[1844] <=  8'h62;        memory[1845] <=  8'h61;        memory[1846] <=  8'h72;        memory[1847] <=  8'h63;        memory[1848] <=  8'h61;        memory[1849] <=  8'h68;        memory[1850] <=  8'h64;        memory[1851] <=  8'h75;        memory[1852] <=  8'h63;        memory[1853] <=  8'h74;        memory[1854] <=  8'h61;        memory[1855] <=  8'h64;        memory[1856] <=  8'h61;        memory[1857] <=  8'h61;        memory[1858] <=  8'h63;        memory[1859] <=  8'h61;        memory[1860] <=  8'h72;        memory[1861] <=  8'h63;        memory[1862] <=  8'h74;        memory[1863] <=  8'h72;        memory[1864] <=  8'h63;        memory[1865] <=  8'h61;        memory[1866] <=  8'h74;        memory[1867] <=  8'h72;        memory[1868] <=  8'h63;        memory[1869] <=  8'h61;        memory[1870] <=  8'h74;        memory[1871] <=  8'h63;        memory[1872] <=  8'h62;        memory[1873] <=  8'h61;        memory[1874] <=  8'h74;        memory[1875] <=  8'h62;        memory[1876] <=  8'h72;        memory[1877] <=  8'h63;        memory[1878] <=  8'h61;        memory[1879] <=  8'h72;        memory[1880] <=  8'h62;        memory[1881] <=  8'h78;        memory[1882] <=  8'h74;        memory[1883] <=  8'h61;        memory[1884] <=  8'h72;        memory[1885] <=  8'h64;        memory[1886] <=  8'h66;        memory[1887] <=  8'h73;        memory[1888] <=  8'h67;        memory[1889] <=  8'h76;        memory[1890] <=  8'h68;        memory[1891] <=  8'h62;        memory[1892] <=  8'h6b;        memory[1893] <=  8'h6a;        memory[1894] <=  8'h6e;        memory[1895] <=  8'h6d;        memory[1896] <=  8'h62;        memory[1897] <=  8'h76;        memory[1898] <=  8'h78;        memory[1899] <=  8'h63;        memory[1900] <=  8'h73;        memory[1901] <=  8'h66;        memory[1902] <=  8'h72;        memory[1903] <=  8'h74;        memory[1904] <=  8'h79;        memory[1905] <=  8'h75;        memory[1906] <=  8'h6a;        memory[1907] <=  8'h6e;        memory[1908] <=  8'h62;        memory[1909] <=  8'h76;        memory[1910] <=  8'h63;        memory[1911] <=  8'h64;        memory[1912] <=  8'h74;        memory[1913] <=  8'h79;        memory[1914] <=  8'h75;        memory[1915] <=  8'h69;        memory[1916] <=  8'h6b;        memory[1917] <=  8'h6d;        memory[1918] <=  8'h6e;        memory[1919] <=  8'h62;        memory[1920] <=  8'h76;        memory[1921] <=  8'h63;        memory[1922] <=  8'h78;        memory[1923] <=  8'h73;        memory[1924] <=  8'h64;        memory[1925] <=  8'h72;        memory[1926] <=  8'h74;        memory[1927] <=  8'h79;        memory[1928] <=  8'h75;        memory[1929] <=  8'h69;        memory[1930] <=  8'h6b;        memory[1931] <=  8'h6d;        memory[1932] <=  8'h6e;        memory[1933] <=  8'h62;        memory[1934] <=  8'h76;        memory[1935] <=  8'h63;        memory[1936] <=  8'h73;        memory[1937] <=  8'h77;        memory[1938] <=  8'h33;        memory[1939] <=  8'h34;        memory[1940] <=  8'h35;        memory[1941] <=  8'h36;        memory[1942] <=  8'h37;        memory[1943] <=  8'h38;        memory[1944] <=  8'h69;        memory[1945] <=  8'h6b;        memory[1946] <=  8'h6d;        memory[1947] <=  8'h6e;        memory[1948] <=  8'h62;        memory[1949] <=  8'h76;        memory[1950] <=  8'h63;        memory[1951] <=  8'h64;        memory[1952] <=  8'h65;        memory[1953] <=  8'h72;        memory[1954] <=  8'h36;        memory[1955] <=  8'h37;        memory[1956] <=  8'h38;        memory[1957] <=  8'h69;        memory[1958] <=  8'h6f;        memory[1959] <=  8'h6b;        memory[1960] <=  8'h6a;        memory[1961] <=  8'h6e;        memory[1962] <=  8'h62;        memory[1963] <=  8'h76;        memory[1964] <=  8'h63;        memory[1965] <=  8'h64;        memory[1966] <=  8'h72;        memory[1967] <=  8'h74;        memory[1968] <=  8'h79;        memory[1969] <=  8'h75;        memory[1970] <=  8'h73;        memory[1971] <=  8'h6a;        memory[1972] <=  8'h63;        memory[1973] <=  8'h6e;        memory[1974] <=  8'h62;        memory[1975] <=  8'h64;        memory[1976] <=  8'h66;        memory[1977] <=  8'h73;        memory[1978] <=  8'h74;        memory[1979] <=  8'h79;        memory[1980] <=  8'h75;        memory[1981] <=  8'h61;        memory[1982] <=  8'h69;        memory[1983] <=  8'h6b;        memory[1984] <=  8'h78;        memory[1985] <=  8'h6d;        memory[1986] <=  8'h6e;        memory[1987] <=  8'h73;        memory[1988] <=  8'h6a;        memory[1989] <=  8'h6f;        memory[1990] <=  8'h64;        memory[1991] <=  8'h6c;        memory[1992] <=  8'h63;        memory[1993] <=  8'h78;        memory[1994] <=  8'h2c;        memory[1995] <=  8'h6d;        memory[1996] <=  8'h73;        memory[1997] <=  8'h6b;        memory[1998] <=  8'h64;        memory[1999] <=  8'h6c;        memory[2000] <=  8'h70;        memory[2001] <=  8'h5b;        memory[2002] <=  8'h3b;        memory[2003] <=  8'h73;        memory[2004] <=  8'h6c;        memory[2005] <=  8'h64;        memory[2006] <=  8'h70;        memory[2007] <=  8'h76;        memory[2008] <=  8'h63;        memory[2009] <=  8'h5b;        memory[2010] <=  8'h78;        memory[2011] <=  8'h76;        memory[2012] <=  8'h63;        memory[2013] <=  8'h5b;        memory[2014] <=  8'h78;        memory[2015] <=  8'h70;        memory[2016] <=  8'h6f;        memory[2017] <=  8'h20;        memory[2018] <=  8'h62;        memory[2019] <=  8'h61;        memory[2020] <=  8'h72;        memory[2021] <=  8'h74;        memory[2022] <=  8'h74;        memory[2023] <=  8'h62;        memory[2024] <=  8'h61;        memory[2025] <=  8'h72;        memory[2026] <=  8'h74;        memory[2027] <=  8'h78;        memory[2028] <=  8'h61;        memory[2029] <=  8'h74;        memory[2030] <=  8'h6b;        memory[2031] <=  8'h73;        memory[2032] <=  8'h68;        memory[2033] <=  8'h63;        memory[2034] <=  8'h66;        memory[2035] <=  8'h69;        memory[2036] <=  8'h77;        memory[2037] <=  8'h68;        memory[2038] <=  8'h61;        memory[2039] <=  8'h69;        memory[2040] <=  8'h6a;        memory[2041] <=  8'h78;        memory[2042] <=  8'h5d;        memory[2043] <=  8'h65;        memory[2044] <=  8'h6b;        memory[2045] <=  8'h6f;        memory[2046] <=  8'h39;        memory[2047] <=  8'h64;        memory[2048] <=  8'h75;        memory[2049] <=  8'h38;        memory[2050] <=  8'h79;        memory[2051] <=  8'h20;        memory[2052] <=  8'h37;        memory[2053] <=  8'h63;        memory[2054] <=  8'h67;        memory[2055] <=  8'h78;        memory[2056] <=  8'h63;        memory[2057] <=  8'h75;        memory[2058] <=  8'h68;        memory[2059] <=  8'h69;        memory[2060] <=  8'h6a;        memory[2061] <=  8'h77;        memory[2062] <=  8'h69;        memory[2063] <=  8'h64;        memory[2064] <=  8'h66;        memory[2065] <=  8'h68;        memory[2066] <=  8'h75;        memory[2067] <=  8'h76;        memory[2068] <=  8'h64;        memory[2069] <=  8'h62;        memory[2070] <=  8'h66;        memory[2071] <=  8'h6a;        memory[2072] <=  8'h6e;        memory[2073] <=  8'h6b;        memory[2074] <=  8'h6a;        memory[2075] <=  8'h65;        memory[2076] <=  8'h38;        memory[2077] <=  8'h66;        memory[2078] <=  8'h37;        memory[2079] <=  8'h67;        memory[2080] <=  8'h79;        memory[2081] <=  8'h76;        memory[2082] <=  8'h63;        memory[2083] <=  8'h68;        memory[2084] <=  8'h69;        memory[2085] <=  8'h6a;        memory[2086] <=  8'h33;        memory[2087] <=  8'h65;        memory[2088] <=  8'h67;        memory[2089] <=  8'h79;        memory[2090] <=  8'h72;        memory[2091] <=  8'h64;        memory[2092] <=  8'h62;        memory[2093] <=  8'h6e;        memory[2094] <=  8'h63;        memory[2095] <=  8'h7a;        memory[2096] <=  8'h6a;        memory[2097] <=  8'h6f;        memory[2098] <=  8'h66;        memory[2099] <=  8'h78;        memory[2100] <=  8'h6a;        memory[2101] <=  8'h69;        memory[2102] <=  8'h63;        memory[2103] <=  8'h68;        memory[2104] <=  8'h62;        memory[2105] <=  8'h6e;        memory[2106] <=  8'h6d;        memory[2107] <=  8'h63;        memory[2108] <=  8'h73;        memory[2109] <=  8'h6c;        memory[2110] <=  8'h6b;        memory[2111] <=  8'h6a;        memory[2112] <=  8'h69;        memory[2113] <=  8'h68;        memory[2114] <=  8'h76;        memory[2115] <=  8'h75;        memory[2116] <=  8'h69;        memory[2117] <=  8'h64;        memory[2118] <=  8'h68;        memory[2119] <=  8'h75;        memory[2120] <=  8'h67;        memory[2121] <=  8'h79;        memory[2122] <=  8'h62;        memory[2123] <=  8'h68;        memory[2124] <=  8'h65;        memory[2125] <=  8'h6a;        memory[2126] <=  8'h72;        memory[2127] <=  8'h6b;        memory[2128] <=  8'h6a;        memory[2129] <=  8'h6f;        memory[2130] <=  8'h64;        memory[2131] <=  8'h67;        memory[2132] <=  8'h69;        memory[2133] <=  8'h75;        memory[2134] <=  8'h69;        memory[2135] <=  8'h67;        memory[2136] <=  8'h76;        memory[2137] <=  8'h79;        memory[2138] <=  8'h75;        memory[2139] <=  8'h67;        memory[2140] <=  8'h78;        memory[2141] <=  8'h68;        memory[2142] <=  8'h63;        memory[2143] <=  8'h20;        memory[2144] <=  8'h20;        memory[2145] <=  8'h20;        memory[2146] <=  8'h78;        memory[2147] <=  8'h76;        memory[2148] <=  8'h20;        memory[2149] <=  8'h63;        memory[2150] <=  8'h78;        memory[2151] <=  8'h67;        memory[2152] <=  8'h79;        memory[2153] <=  8'h63;        memory[2154] <=  8'h75;        memory[2155] <=  8'h68;        memory[2156] <=  8'h6a;        memory[2157] <=  8'h6b;        memory[2158] <=  8'h61;        memory[2159] <=  8'h6c;        memory[2160] <=  8'h78;        memory[2161] <=  8'h76;        memory[2162] <=  8'h70;        memory[2163] <=  8'h6f;        memory[2164] <=  8'h69;        memory[2165] <=  8'h6a;        memory[2166] <=  8'h69;        memory[2167] <=  8'h68;        memory[2168] <=  8'h6a;        memory[2169] <=  8'h62;        memory[2170] <=  8'h77;        memory[2171] <=  8'h65;        memory[2172] <=  8'h6e;        memory[2173] <=  8'h61;        memory[2174] <=  8'h66;        memory[2175] <=  8'h6d;        memory[2176] <=  8'h64;        memory[2177] <=  8'h6b;        memory[2178] <=  8'h6d;        memory[2179] <=  8'h76;        memory[2180] <=  8'h6c;        memory[2181] <=  8'h63;        memory[2182] <=  8'h6f;        memory[2183] <=  8'h64;        memory[2184] <=  8'h69;        memory[2185] <=  8'h75;        memory[2186] <=  8'h68;        memory[2187] <=  8'h73;        memory[2188] <=  8'h66;        memory[2189] <=  8'h65;        memory[2190] <=  8'h62;        memory[2191] <=  8'h6e;        memory[2192] <=  8'h64;        memory[2193] <=  8'h73;        memory[2194] <=  8'h63;        memory[2195] <=  8'h6b;        memory[2196] <=  8'h20;        memory[2197] <=  8'h78;        memory[2198] <=  8'h6a;        memory[2199] <=  8'h78;        memory[2200] <=  8'h63;        memory[2201] <=  8'h73;        memory[2202] <=  8'h64;        memory[2203] <=  8'h66;        memory[2204] <=  8'h6b;        memory[2205] <=  8'h64;        memory[2206] <=  8'h6e;        memory[2207] <=  8'h6d;        memory[2208] <=  8'h64;        memory[2209] <=  8'h73;        memory[2210] <=  8'h63;        memory[2211] <=  8'h6b;        memory[2212] <=  8'h78;        memory[2213] <=  8'h6c;        memory[2214] <=  8'h6f;        memory[2215] <=  8'h66;        memory[2216] <=  8'h6a;        memory[2217] <=  8'h69;        memory[2218] <=  8'h61;        memory[2219] <=  8'h62;        memory[2220] <=  8'h6e;        memory[2221] <=  8'h20;        memory[2222] <=  8'h78;        memory[2223] <=  8'h6b;        memory[2224] <=  8'h6d;        memory[2225] <=  8'h20;        memory[2226] <=  8'h6f;        memory[2227] <=  8'h63;        memory[2228] <=  8'h76;        memory[2229] <=  8'h73;        memory[2230] <=  8'h64;        memory[2231] <=  8'h69;        memory[2232] <=  8'h66;        memory[2233] <=  8'h68;        memory[2234] <=  8'h65;        memory[2235] <=  8'h71;        memory[2236] <=  8'h6a;        memory[2237] <=  8'h77;        memory[2238] <=  8'h62;        memory[2239] <=  8'h65;        memory[2240] <=  8'h6e;        memory[2241] <=  8'h20;        memory[2242] <=  8'h6d;        memory[2243] <=  8'h64;        memory[2244] <=  8'h73;        memory[2245] <=  8'h6c;        memory[2246] <=  8'h76;        memory[2247] <=  8'h6b;        memory[2248] <=  8'h63;        memory[2249] <=  8'h78;        memory[2250] <=  8'h20;        memory[2251] <=  8'h6f;        memory[2252] <=  8'h78;        memory[2253] <=  8'h69;        memory[2254] <=  8'h63;        memory[2255] <=  8'h6a;        memory[2256] <=  8'h76;        memory[2257] <=  8'h64;        memory[2258] <=  8'h66;        memory[2259] <=  8'h65;        memory[2260] <=  8'h71;        memory[2261] <=  8'h6e;        memory[2262] <=  8'h20;        memory[2263] <=  8'h64;        memory[2264] <=  8'h6d;        memory[2265] <=  8'h73;        memory[2266] <=  8'h6c;        memory[2267] <=  8'h63;        memory[2268] <=  8'h78;        memory[2269] <=  8'h6b;        memory[2270] <=  8'h20;        memory[2271] <=  8'h6f;        memory[2272] <=  8'h78;        memory[2273] <=  8'h63;        memory[2274] <=  8'h76;        memory[2275] <=  8'h6a;        memory[2276] <=  8'h64;        memory[2277] <=  8'h62;        memory[2278] <=  8'h71;        memory[2279] <=  8'h77;        memory[2280] <=  8'h65;        memory[2281] <=  8'h6e;        memory[2282] <=  8'h6d;        memory[2283] <=  8'h64;        memory[2284] <=  8'h6c;        memory[2285] <=  8'h73;        memory[2286] <=  8'h2c;        memory[2287] <=  8'h76;        memory[2288] <=  8'h63;        memory[2289] <=  8'h78;        memory[2290] <=  8'h20;        memory[2291] <=  8'h63;        memory[2292] <=  8'h6f;        memory[2293] <=  8'h69;        memory[2294] <=  8'h76;        memory[2295] <=  8'h68;        memory[2296] <=  8'h73;        memory[2297] <=  8'h64;        memory[2298] <=  8'h62;        memory[2299] <=  8'h71;        memory[2300] <=  8'h77;        memory[2301] <=  8'h65;        memory[2302] <=  8'h6e;        memory[2303] <=  8'h64;        memory[2304] <=  8'h6b;        memory[2305] <=  8'h73;        memory[2306] <=  8'h76;        memory[2307] <=  8'h6f;        memory[2308] <=  8'h63;        memory[2309] <=  8'h20;        memory[2310] <=  8'h76;        memory[2311] <=  8'h69;        memory[2312] <=  8'h75;        memory[2313] <=  8'h69;        memory[2314] <=  8'h68;        memory[2315] <=  8'h63;        memory[2316] <=  8'h78;        memory[2317] <=  8'h69;        memory[2318] <=  8'h6f;        memory[2319] <=  8'h76;        memory[2320] <=  8'h73;        memory[2321] <=  8'h64;        memory[2322] <=  8'h61;        memory[2323] <=  8'h64;        memory[2324] <=  8'h6e;        memory[2325] <=  8'h77;        memory[2326] <=  8'h71;        memory[2327] <=  8'h6b;        memory[2328] <=  8'h6c;        memory[2329] <=  8'h73;        memory[2330] <=  8'h76;        memory[2331] <=  8'h6e;        memory[2332] <=  8'h62;        memory[2333] <=  8'h20;        memory[2334] <=  8'h64;        memory[2335] <=  8'h66;        memory[2336] <=  8'h6a;        memory[2337] <=  8'h6b;        memory[2338] <=  8'h71;        memory[2339] <=  8'h64;        memory[2340] <=  8'h77;        memory[2341] <=  8'h65;        memory[2342] <=  8'h6e;        memory[2343] <=  8'h62;        memory[2344] <=  8'h20;        memory[2345] <=  8'h64;        memory[2346] <=  8'h73;        memory[2347] <=  8'h76;        memory[2348] <=  8'h68;        memory[2349] <=  8'h64;        memory[2350] <=  8'h61;        memory[2351] <=  8'h71;        memory[2352] <=  8'h77;        memory[2353] <=  8'h6a;        memory[2354] <=  8'h65;        memory[2355] <=  8'h6e;        memory[2356] <=  8'h64;        memory[2357] <=  8'h20;        memory[2358] <=  8'h61;        memory[2359] <=  8'h63;        memory[2360] <=  8'h62;        memory[2361] <=  8'h68;        memory[2362] <=  8'h64;        memory[2363] <=  8'h61;        memory[2364] <=  8'h77;        memory[2365] <=  8'h71;        memory[2366] <=  8'h6e;        memory[2367] <=  8'h20;        memory[2368] <=  8'h62;        memory[2369] <=  8'h73;        memory[2370] <=  8'h76;        memory[2371] <=  8'h61;        memory[2372] <=  8'h67;        memory[2373] <=  8'h76;        memory[2374] <=  8'h68;        memory[2375] <=  8'h67;        memory[2376] <=  8'h61;        memory[2377] <=  8'h73;        memory[2378] <=  8'h6a;        memory[2379] <=  8'h6b;        memory[2380] <=  8'h63;        memory[2381] <=  8'h78;        memory[2382] <=  8'h76;        memory[2383] <=  8'h6e;        memory[2384] <=  8'h73;        memory[2385] <=  8'h64;        memory[2386] <=  8'h20;        memory[2387] <=  8'h66;        memory[2388] <=  8'h62;        memory[2389] <=  8'h64;        memory[2390] <=  8'h61;        memory[2391] <=  8'h73;        memory[2392] <=  8'h76;        memory[2393] <=  8'h67;        memory[2394] <=  8'h63;        memory[2395] <=  8'h79;        memory[2396] <=  8'h7a;        memory[2397] <=  8'h78;        memory[2398] <=  8'h79;        memory[2399] <=  8'h75;        memory[2400] <=  8'h20;        memory[2401] <=  8'h69;        memory[2402] <=  8'h6a;        memory[2403] <=  8'h64;        memory[2404] <=  8'h66;        memory[2405] <=  8'h6b;        memory[2406] <=  8'h61;        memory[2407] <=  8'h64;        memory[2408] <=  8'h63;        memory[2409] <=  8'h78;        memory[2410] <=  8'h68;        memory[2411] <=  8'h20;        memory[2412] <=  8'h67;        memory[2413] <=  8'h61;        memory[2414] <=  8'h68;        memory[2415] <=  8'h75;        memory[2416] <=  8'h64;        memory[2417] <=  8'h73;        memory[2418] <=  8'h69;        memory[2419] <=  8'h6a;        memory[2420] <=  8'h61;        memory[2421] <=  8'h6b;        memory[2422] <=  8'h63;        memory[2423] <=  8'h62;        memory[2424] <=  8'h61;        memory[2425] <=  8'h72;        memory[2426] <=  8'h73;        memory[2427] <=  8'h68;        memory[2428] <=  8'h64;        memory[2429] <=  8'h66;        memory[2430] <=  8'h67;        memory[2431] <=  8'h73;        memory[2432] <=  8'h68;        memory[2433] <=  8'h64;        memory[2434] <=  8'h66;        memory[2435] <=  8'h68;        memory[2436] <=  8'h64;        memory[2437] <=  8'h6a;        memory[2438] <=  8'h68;        memory[2439] <=  8'h62;        memory[2440] <=  8'h67;        memory[2441] <=  8'h63;        memory[2442] <=  8'h61;        memory[2443] <=  8'h66;        memory[2444] <=  8'h73;        memory[2445] <=  8'h79;        memory[2446] <=  8'h67;        memory[2447] <=  8'h6b;        memory[2448] <=  8'h75;        memory[2449] <=  8'h64;        memory[2450] <=  8'h68;        memory[2451] <=  8'h62;        memory[2452] <=  8'h77;        memory[2453] <=  8'h76;        memory[2454] <=  8'h67;        memory[2455] <=  8'h61;        memory[2456] <=  8'h66;        memory[2457] <=  8'h64;        memory[2458] <=  8'h74;        memory[2459] <=  8'h75;        memory[2460] <=  8'h66;        memory[2461] <=  8'h79;        memory[2462] <=  8'h67;        memory[2463] <=  8'h69;        memory[2464] <=  8'h75;        memory[2465] <=  8'h68;        memory[2466] <=  8'h6c;        memory[2467] <=  8'h6a;        memory[2468] <=  8'h62;        memory[2469] <=  8'h6b;        memory[2470] <=  8'h68;        memory[2471] <=  8'h76;        memory[2472] <=  8'h67;        memory[2473] <=  8'h63;        memory[2474] <=  8'h66;        memory[2475] <=  8'h78;        memory[2476] <=  8'h64;        memory[2477] <=  8'h74;        memory[2478] <=  8'h75;        memory[2479] <=  8'h79;        memory[2480] <=  8'h69;        memory[2481] <=  8'h75;        memory[2482] <=  8'h68;        memory[2483] <=  8'h6c;        memory[2484] <=  8'h6a;        memory[2485] <=  8'h6b;        memory[2486] <=  8'h67;        memory[2487] <=  8'h6a;        memory[2488] <=  8'h63;        memory[2489] <=  8'h66;        memory[2490] <=  8'h68;        memory[2491] <=  8'h64;        memory[2492] <=  8'h67;        memory[2493] <=  8'h72;        memory[2494] <=  8'h79;        memory[2495] <=  8'h74;        memory[2496] <=  8'h66;        memory[2497] <=  8'h75;        memory[2498] <=  8'h79;        memory[2499] <=  8'h69;        memory[2500] <=  8'h68;        memory[2501] <=  8'h6c;        memory[2502] <=  8'h62;        memory[2503] <=  8'h6d;        memory[2504] <=  8'h76;        memory[2505] <=  8'h6e;        memory[2506] <=  8'h63;        memory[2507] <=  8'h66;        memory[2508] <=  8'h68;        memory[2509] <=  8'h64;        memory[2510] <=  8'h74;        memory[2511] <=  8'h75;        memory[2512] <=  8'h67;        memory[2513] <=  8'h79;        memory[2514] <=  8'h69;        memory[2515] <=  8'h68;        memory[2516] <=  8'h75;        memory[2517] <=  8'h6a;        memory[2518] <=  8'h6c;        memory[2519] <=  8'h62;        memory[2520] <=  8'h6d;        memory[2521] <=  8'h76;        memory[2522] <=  8'h6e;        memory[2523] <=  8'h63;        memory[2524] <=  8'h66;        memory[2525] <=  8'h68;        memory[2526] <=  8'h67;        memory[2527] <=  8'h79;        memory[2528] <=  8'h68;        memory[2529] <=  8'h75;        memory[2530] <=  8'h6a;        memory[2531] <=  8'h6e;        memory[2532] <=  8'h2c;        memory[2533] <=  8'h62;        memory[2534] <=  8'h6e;        memory[2535] <=  8'h6d;        memory[2536] <=  8'h76;        memory[2537] <=  8'h6e;        memory[2538] <=  8'h63;        memory[2539] <=  8'h66;        memory[2540] <=  8'h68;        memory[2541] <=  8'h74;        memory[2542] <=  8'h79;        memory[2543] <=  8'h69;        memory[2544] <=  8'h75;        memory[2545] <=  8'h6c;        memory[2546] <=  8'h6a;        memory[2547] <=  8'h62;        memory[2548] <=  8'h6d;        memory[2549] <=  8'h76;        memory[2550] <=  8'h6e;        memory[2551] <=  8'h63;        memory[2552] <=  8'h66;        memory[2553] <=  8'h74;        memory[2554] <=  8'h75;        memory[2555] <=  8'h79;        memory[2556] <=  8'h69;        memory[2557] <=  8'h68;        memory[2558] <=  8'h6b;        memory[2559] <=  8'h62;        memory[2560] <=  8'h76;        memory[2561] <=  8'h63;        memory[2562] <=  8'h66;        memory[2563] <=  8'h67;        memory[2564] <=  8'h74;        memory[2565] <=  8'h75;        memory[2566] <=  8'h79;        memory[2567] <=  8'h69;        memory[2568] <=  8'h75;        memory[2569] <=  8'h68;        memory[2570] <=  8'h6a;        memory[2571] <=  8'h6b;        memory[2572] <=  8'h62;        memory[2573] <=  8'h76;        memory[2574] <=  8'h63;        memory[2575] <=  8'h66;        memory[2576] <=  8'h74;        memory[2577] <=  8'h75;        memory[2578] <=  8'h79;        memory[2579] <=  8'h69;        memory[2580] <=  8'h75;        memory[2581] <=  8'h6a;        memory[2582] <=  8'h6b;        memory[2583] <=  8'h6e;        memory[2584] <=  8'h62;        memory[2585] <=  8'h76;        memory[2586] <=  8'h67;        memory[2587] <=  8'h66;        memory[2588] <=  8'h74;        memory[2589] <=  8'h79;        memory[2590] <=  8'h75;        memory[2591] <=  8'h75;        memory[2592] <=  8'h69;        memory[2593] <=  8'h6a;        memory[2594] <=  8'h6b;        memory[2595] <=  8'h68;        memory[2596] <=  8'h62;        memory[2597] <=  8'h6a;        memory[2598] <=  8'h67;        memory[2599] <=  8'h68;        memory[2600] <=  8'h66;        memory[2601] <=  8'h79;        memory[2602] <=  8'h74;        memory[2603] <=  8'h79;        memory[2604] <=  8'h69;        memory[2605] <=  8'h75;        memory[2606] <=  8'h64;        memory[2607] <=  8'h6a;        memory[2608] <=  8'h6b;        memory[2609] <=  8'h68;        memory[2610] <=  8'h63;        memory[2611] <=  8'h7a;        memory[2612] <=  8'h67;        memory[2613] <=  8'h68;        memory[2614] <=  8'h74;        memory[2615] <=  8'h75;        memory[2616] <=  8'h79;        memory[2617] <=  8'h69;        memory[2618] <=  8'h61;        memory[2619] <=  8'h73;        memory[2620] <=  8'h75;        memory[2621] <=  8'h6a;        memory[2622] <=  8'h6b;        memory[2623] <=  8'h62;        memory[2624] <=  8'h6e;        memory[2625] <=  8'h61;        memory[2626] <=  8'h76;        memory[2627] <=  8'h63;        memory[2628] <=  8'h66;        memory[2629] <=  8'h68;        memory[2630] <=  8'h75;        memory[2631] <=  8'h61;        memory[2632] <=  8'h73;        memory[2633] <=  8'h79;        memory[2634] <=  8'h64;        memory[2635] <=  8'h75;        memory[2636] <=  8'h69;        memory[2637] <=  8'h6a;        memory[2638] <=  8'h61;        memory[2639] <=  8'h6b;        memory[2640] <=  8'h62;        memory[2641] <=  8'h63;        memory[2642] <=  8'h78;        memory[2643] <=  8'h68;        memory[2644] <=  8'h67;        memory[2645] <=  8'h79;        memory[2646] <=  8'h75;        memory[2647] <=  8'h7a;        memory[2648] <=  8'h63;        memory[2649] <=  8'h61;        memory[2650] <=  8'h73;        memory[2651] <=  8'h69;        memory[2652] <=  8'h75;        memory[2653] <=  8'h6f;        memory[2654] <=  8'h69;        memory[2655] <=  8'h6a;        memory[2656] <=  8'h61;        memory[2657] <=  8'h6c;        memory[2658] <=  8'h63;        memory[2659] <=  8'h78;        memory[2660] <=  8'h62;        memory[2661] <=  8'h63;        memory[2662] <=  8'h20;        memory[2663] <=  8'h6e;        memory[2664] <=  8'h76;        memory[2665] <=  8'h63;        memory[2666] <=  8'h61;        memory[2667] <=  8'h64;        memory[2668] <=  8'h73;        memory[2669] <=  8'h67;        memory[2670] <=  8'h79;        memory[2671] <=  8'h68;        memory[2672] <=  8'h75;        memory[2673] <=  8'h61;        memory[2674] <=  8'h6a;        memory[2675] <=  8'h6b;        memory[2676] <=  8'h78;        memory[2677] <=  8'h62;        memory[2678] <=  8'h20;        memory[2679] <=  8'h6e;        memory[2680] <=  8'h76;        memory[2681] <=  8'h63;        memory[2682] <=  8'h61;        memory[2683] <=  8'h73;        memory[2684] <=  8'h67;        memory[2685] <=  8'h68;        memory[2686] <=  8'h75;        memory[2687] <=  8'h6a;        memory[2688] <=  8'h6c;        memory[2689] <=  8'h6b;        memory[2690] <=  8'h63;        memory[2691] <=  8'h78;        memory[2692] <=  8'h20;        memory[2693] <=  8'h6a;        memory[2694] <=  8'h6b;        memory[2695] <=  8'h68;        memory[2696] <=  8'h61;        memory[2697] <=  8'h73;        memory[2698] <=  8'h76;        memory[2699] <=  8'h64;        memory[2700] <=  8'h6e;        memory[2701] <=  8'h20;        memory[2702] <=  8'h62;        memory[2703] <=  8'h6e;        memory[2704] <=  8'h6d;        memory[2705] <=  8'h6b;        memory[2706] <=  8'h77;        memory[2707] <=  8'h64;        memory[2708] <=  8'h6f;        memory[2709] <=  8'h77;        memory[2710] <=  8'h69;        memory[2711] <=  8'h6f;        memory[2712] <=  8'h75;        memory[2713] <=  8'h69;        memory[2714] <=  8'h68;        memory[2715] <=  8'h62;        memory[2716] <=  8'h6e;        memory[2717] <=  8'h6b;        memory[2718] <=  8'h77;        memory[2719] <=  8'h69;        memory[2720] <=  8'h6f;        memory[2721] <=  8'h75;        memory[2722] <=  8'h71;        memory[2723] <=  8'h69;        memory[2724] <=  8'h79;        memory[2725] <=  8'h67;        memory[2726] <=  8'h6a;        memory[2727] <=  8'h64;        memory[2728] <=  8'h61;        memory[2729] <=  8'h76;        memory[2730] <=  8'h62;        memory[2731] <=  8'h6e;        memory[2732] <=  8'h6b;        memory[2733] <=  8'h6f;        memory[2734] <=  8'h70;        memory[2735] <=  8'h64;        memory[2736] <=  8'h76;        memory[2737] <=  8'h69;        memory[2738] <=  8'h6f;        memory[2739] <=  8'h75;        memory[2740] <=  8'h69;        memory[2741] <=  8'h48;        memory[2742] <=  8'h42;        memory[2743] <=  8'h6b;        memory[2744] <=  8'h64;        memory[2745] <=  8'h6e;        memory[2746] <=  8'h6c;        memory[2747] <=  8'h71;        memory[2748] <=  8'h6b;        memory[2749] <=  8'h6d;        memory[2750] <=  8'h6a;        memory[2751] <=  8'h70;        memory[2752] <=  8'h69;        memory[2753] <=  8'h6f;        memory[2754] <=  8'h68;        memory[2755] <=  8'h65;        memory[2756] <=  8'h66;        memory[2757] <=  8'h75;        memory[2758] <=  8'h67;        memory[2759] <=  8'h69;        memory[2760] <=  8'h73;        memory[2761] <=  8'h61;        memory[2762] <=  8'h62;        memory[2763] <=  8'h64;        memory[2764] <=  8'h6b;        memory[2765] <=  8'h6a;        memory[2766] <=  8'h6b;        memory[2767] <=  8'h6c;        memory[2768] <=  8'h6a;        memory[2769] <=  8'h69;        memory[2770] <=  8'h73;        memory[2771] <=  8'h6f;        memory[2772] <=  8'h71;        memory[2773] <=  8'h68;        memory[2774] <=  8'h77;        memory[2775] <=  8'h67;        memory[2776] <=  8'h69;        memory[2777] <=  8'h79;        memory[2778] <=  8'h6a;        memory[2779] <=  8'h64;        memory[2780] <=  8'h76;        memory[2781] <=  8'h62;        memory[2782] <=  8'h6e;        memory[2783] <=  8'h61;        memory[2784] <=  8'h73;        memory[2785] <=  8'h66;        memory[2786] <=  8'h6c;        memory[2787] <=  8'h6b;        memory[2788] <=  8'h64;        memory[2789] <=  8'h6a;        memory[2790] <=  8'h68;        memory[2791] <=  8'h63;        memory[2792] <=  8'h67;        memory[2793] <=  8'h6a;        memory[2794] <=  8'h76;        memory[2795] <=  8'h73;        memory[2796] <=  8'h64;        memory[2797] <=  8'h62;        memory[2798] <=  8'h62;        memory[2799] <=  8'h61;        memory[2800] <=  8'h72;        memory[2801] <=  8'h62;        memory[2802] <=  8'h62;        memory[2803] <=  8'h73;        memory[2804] <=  8'h62;        memory[2805] <=  8'h67;        memory[2806] <=  8'h73;        memory[2807] <=  8'h66;        memory[2808] <=  8'h67;        memory[2809] <=  8'h61;        memory[2810] <=  8'h68;        memory[2811] <=  8'h66;        memory[2812] <=  8'h73;        memory[2813] <=  8'h68;        memory[2814] <=  8'h61;        memory[2815] <=  8'h66;        memory[2816] <=  8'h73;        memory[2817] <=  8'h66;        memory[2818] <=  8'h68;        memory[2819] <=  8'h61;        memory[2820] <=  8'h69;        memory[2821] <=  8'h64;        memory[2822] <=  8'h75;        memory[2823] <=  8'h67;        memory[2824] <=  8'h64;        memory[2825] <=  8'h77;        memory[2826] <=  8'h62;        memory[2827] <=  8'h61;        memory[2828] <=  8'h62;        memory[2829] <=  8'h72;        memory[2830] <=  8'h62;        memory[2831] <=  8'h61;        memory[2832] <=  8'h62;        memory[2833] <=  8'h62;        memory[2834] <=  8'h74;        memory[2835] <=  8'h62;        memory[2836] <=  8'h62;        memory[2837] <=  8'h62;        memory[2838] <=  8'h62;        memory[2839] <=  8'h62;        memory[2840] <=  8'h62;        memory[2841] <=  8'h62;        memory[2842] <=  8'h62;        memory[2843] <=  8'h61;        memory[2844] <=  8'h62;        memory[2845] <=  8'h62;        memory[2846] <=  8'h72;        memory[2847] <=  8'h74;        memory[2848] <=  8'h62;        memory[2849] <=  8'h62;        memory[2850] <=  8'h61;        memory[2851] <=  8'h62;        memory[2852] <=  8'h72;        memory[2853] <=  8'h62;        memory[2854] <=  8'h74;        memory[2855] <=  8'h62;        memory[2856] <=  8'h62;        memory[2857] <=  8'h62;        memory[2858] <=  8'h63;        memory[2859] <=  8'h61;        memory[2860] <=  8'h72;        memory[2861] <=  8'h74;        memory[2862] <=  8'h73;        memory[2863] <=  8'h62;        memory[2864] <=  8'h61;        memory[2865] <=  8'h72;        memory[2866] <=  8'h74;        memory[2867] <=  8'h74;        memory[2868] <=  8'h62;        memory[2869] <=  8'h61;        memory[2870] <=  8'h72;        memory[2871] <=  8'h74;        memory[2872] <=  8'h78;        memory[2873] <=  8'h61;        memory[2874] <=  8'h74;        memory[2875] <=  8'h6b;        memory[2876] <=  8'h73;        memory[2877] <=  8'h68;        memory[2878] <=  8'h63;        memory[2879] <=  8'h66;        memory[2880] <=  8'h69;        memory[2881] <=  8'h77;        memory[2882] <=  8'h68;        memory[2883] <=  8'h61;        memory[2884] <=  8'h74;        memory[2885] <=  8'h61;        memory[2886] <=  8'h6e;        memory[2887] <=  8'h61;        memory[2888] <=  8'h62;        memory[2889] <=  8'h61;        memory[2890] <=  8'h63;        memory[2891] <=  8'h61;        memory[2892] <=  8'h74;        memory[2893] <=  8'h61;        memory[2894] <=  8'h62;        memory[2895] <=  8'h61;        memory[2896] <=  8'h72;        memory[2897] <=  8'h63;        memory[2898] <=  8'h61;        memory[2899] <=  8'h68;        memory[2900] <=  8'h64;        memory[2901] <=  8'h75;        memory[2902] <=  8'h63;        memory[2903] <=  8'h74;        memory[2904] <=  8'h61;        memory[2905] <=  8'h64;        memory[2906] <=  8'h61;        memory[2907] <=  8'h61;        memory[2908] <=  8'h63;        memory[2909] <=  8'h61;        memory[2910] <=  8'h72;        memory[2911] <=  8'h63;        memory[2912] <=  8'h74;        memory[2913] <=  8'h72;        memory[2914] <=  8'h63;        memory[2915] <=  8'h61;        memory[2916] <=  8'h74;        memory[2917] <=  8'h72;        memory[2918] <=  8'h63;        memory[2919] <=  8'h61;        memory[2920] <=  8'h74;        memory[2921] <=  8'h63;        memory[2922] <=  8'h62;        memory[2923] <=  8'h61;        memory[2924] <=  8'h74;        memory[2925] <=  8'h62;        memory[2926] <=  8'h72;        memory[2927] <=  8'h63;        memory[2928] <=  8'h61;        memory[2929] <=  8'h74;        memory[2930] <=  8'h72;        memory[2931] <=  8'h6e;        memory[2932] <=  8'h62;        memory[2933] <=  8'h61;        memory[2934] <=  8'h63;        memory[2935] <=  8'h61;        memory[2936] <=  8'h74;        memory[2937] <=  8'h79;        memory[2938] <=  8'h73;        memory[2939] <=  8'h6e;        memory[2940] <=  8'h63;        memory[2941] <=  8'h74;        memory[2942] <=  8'h61;        memory[2943] <=  8'h6e;        memory[2944] <=  8'h62;        memory[2945] <=  8'h61;        memory[2946] <=  8'h63;        memory[2947] <=  8'h72;        memory[2948] <=  8'h6e;        memory[2949] <=  8'h74;        memory[2950] <=  8'h61;        memory[2951] <=  8'h62;        memory[2952] <=  8'h74;        memory[2953] <=  8'h6e;        memory[2954] <=  8'h61;        memory[2955] <=  8'h72;        memory[2956] <=  8'h62;        memory[2957] <=  8'h78;        memory[2958] <=  8'h74;        memory[2959] <=  8'h61;        memory[2960] <=  8'h72;        memory[2961] <=  8'h62;        memory[2962] <=  8'h61;        memory[2963] <=  8'h72;        memory[2964] <=  8'h74;        memory[2965] <=  8'h74;        memory[2966] <=  8'h62;        memory[2967] <=  8'h61;        memory[2968] <=  8'h72;        memory[2969] <=  8'h74;        memory[2970] <=  8'h78;        memory[2971] <=  8'h61;        memory[2972] <=  8'h74;        memory[2973] <=  8'h6b;        memory[2974] <=  8'h73;        memory[2975] <=  8'h68;        memory[2976] <=  8'h63;        memory[2977] <=  8'h66;        memory[2978] <=  8'h69;        memory[2979] <=  8'h77;        memory[2980] <=  8'h68;        memory[2981] <=  8'h61;        memory[2982] <=  8'h74;        memory[2983] <=  8'h61;        memory[2984] <=  8'h6e;        memory[2985] <=  8'h61;        memory[2986] <=  8'h62;        memory[2987] <=  8'h61;        memory[2988] <=  8'h63;        memory[2989] <=  8'h61;        memory[2990] <=  8'h74;        memory[2991] <=  8'h61;        memory[2992] <=  8'h62;        memory[2993] <=  8'h61;        memory[2994] <=  8'h72;        memory[2995] <=  8'h63;        memory[2996] <=  8'h61;        memory[2997] <=  8'h68;        memory[2998] <=  8'h64;        memory[2999] <=  8'h75;        memory[3000] <=  8'h63;        memory[3001] <=  8'h74;        memory[3002] <=  8'h61;        memory[3003] <=  8'h64;        memory[3004] <=  8'h61;        memory[3005] <=  8'h61;        memory[3006] <=  8'h63;        memory[3007] <=  8'h61;        memory[3008] <=  8'h72;        memory[3009] <=  8'h63;        memory[3010] <=  8'h74;        memory[3011] <=  8'h72;        memory[3012] <=  8'h63;        memory[3013] <=  8'h61;        memory[3014] <=  8'h74;        memory[3015] <=  8'h72;        memory[3016] <=  8'h63;        memory[3017] <=  8'h61;        memory[3018] <=  8'h74;        memory[3019] <=  8'h63;        memory[3020] <=  8'h62;        memory[3021] <=  8'h61;        memory[3022] <=  8'h74;        memory[3023] <=  8'h62;        memory[3024] <=  8'h72;        memory[3025] <=  8'h63;        memory[3026] <=  8'h61;        memory[3027] <=  8'h74;        memory[3028] <=  8'h72;        memory[3029] <=  8'h6e;        memory[3030] <=  8'h62;        memory[3031] <=  8'h61;        memory[3032] <=  8'h63;        memory[3033] <=  8'h61;        memory[3034] <=  8'h74;        memory[3035] <=  8'h79;        memory[3036] <=  8'h73;        memory[3037] <=  8'h6e;        memory[3038] <=  8'h63;        memory[3039] <=  8'h74;        memory[3040] <=  8'h61;        memory[3041] <=  8'h6e;        memory[3042] <=  8'h62;        memory[3043] <=  8'h61;        memory[3044] <=  8'h63;        memory[3045] <=  8'h72;        memory[3046] <=  8'h6e;        memory[3047] <=  8'h74;        memory[3048] <=  8'h61;        memory[3049] <=  8'h62;        memory[3050] <=  8'h74;        memory[3051] <=  8'h6e;        memory[3052] <=  8'h61;        memory[3053] <=  8'h72;        memory[3054] <=  8'h62;        memory[3055] <=  8'h78;        memory[3056] <=  8'h74;        memory[3057] <=  8'h61;        memory[3058] <=  8'h72;        memory[3059] <=  8'h62;        memory[3060] <=  8'h61;        memory[3061] <=  8'h72;        memory[3062] <=  8'h74;        memory[3063] <=  8'h74;        memory[3064] <=  8'h62;        memory[3065] <=  8'h61;        memory[3066] <=  8'h72;        memory[3067] <=  8'h74;        memory[3068] <=  8'h78;        memory[3069] <=  8'h61;        memory[3070] <=  8'h74;        memory[3071] <=  8'h6b;        memory[3072] <=  8'h73;        memory[3073] <=  8'h68;        memory[3074] <=  8'h63;        memory[3075] <=  8'h66;        memory[3076] <=  8'h69;        memory[3077] <=  8'h77;        memory[3078] <=  8'h68;        memory[3079] <=  8'h61;        memory[3080] <=  8'h74;        memory[3081] <=  8'h61;        memory[3082] <=  8'h6e;        memory[3083] <=  8'h61;        memory[3084] <=  8'h62;        memory[3085] <=  8'h61;        memory[3086] <=  8'h63;        memory[3087] <=  8'h61;        memory[3088] <=  8'h74;        memory[3089] <=  8'h61;        memory[3090] <=  8'h62;        memory[3091] <=  8'h61;        memory[3092] <=  8'h72;        memory[3093] <=  8'h63;        memory[3094] <=  8'h61;        memory[3095] <=  8'h68;        memory[3096] <=  8'h64;        memory[3097] <=  8'h75;        memory[3098] <=  8'h63;        memory[3099] <=  8'h74;        memory[3100] <=  8'h61;        memory[3101] <=  8'h64;        memory[3102] <=  8'h61;        memory[3103] <=  8'h61;        memory[3104] <=  8'h63;        memory[3105] <=  8'h61;        memory[3106] <=  8'h72;        memory[3107] <=  8'h63;        memory[3108] <=  8'h74;        memory[3109] <=  8'h72;        memory[3110] <=  8'h63;        memory[3111] <=  8'h61;        memory[3112] <=  8'h74;        memory[3113] <=  8'h72;        memory[3114] <=  8'h63;        memory[3115] <=  8'h61;        memory[3116] <=  8'h74;        memory[3117] <=  8'h63;        memory[3118] <=  8'h62;        memory[3119] <=  8'h61;        memory[3120] <=  8'h74;        memory[3121] <=  8'h62;        memory[3122] <=  8'h72;        memory[3123] <=  8'h63;        memory[3124] <=  8'h61;        memory[3125] <=  8'h74;        memory[3126] <=  8'h72;        memory[3127] <=  8'h6e;        memory[3128] <=  8'h62;        memory[3129] <=  8'h61;        memory[3130] <=  8'h63;        memory[3131] <=  8'h61;        memory[3132] <=  8'h74;        memory[3133] <=  8'h79;        memory[3134] <=  8'h73;        memory[3135] <=  8'h6e;        memory[3136] <=  8'h63;        memory[3137] <=  8'h74;        memory[3138] <=  8'h61;        memory[3139] <=  8'h6e;        memory[3140] <=  8'h62;        memory[3141] <=  8'h61;        memory[3142] <=  8'h63;        memory[3143] <=  8'h72;        memory[3144] <=  8'h6e;        memory[3145] <=  8'h74;        memory[3146] <=  8'h61;        memory[3147] <=  8'h62;        memory[3148] <=  8'h74;        memory[3149] <=  8'h6e;        memory[3150] <=  8'h61;        memory[3151] <=  8'h72;        memory[3152] <=  8'h62;        memory[3153] <=  8'h78;        memory[3154] <=  8'h74;        memory[3155] <=  8'h61;        memory[3156] <=  8'h72;        memory[3157] <=  8'h5d;        memory[3158] <=  8'h5d;        memory[3159] <=  8'h65;        memory[3160] <=  8'h66;        memory[3161] <=  8'h77;        memory[3162] <=  8'h65;        memory[3163] <=  8'h5d;        memory[3164] <=  8'h65;        memory[3165] <=  8'h67;        memory[3166] <=  8'h73;        memory[3167] <=  8'h67;        memory[3168] <=  8'h66;        memory[3169] <=  8'h62;        memory[3170] <=  8'h61;        memory[3171] <=  8'h72;        memory[3172] <=  8'h74;        memory[3173] <=  8'h74;        memory[3174] <=  8'h62;        memory[3175] <=  8'h61;        memory[3176] <=  8'h72;        memory[3177] <=  8'h74;        memory[3178] <=  8'h78;        memory[3179] <=  8'h61;        memory[3180] <=  8'h74;        memory[3181] <=  8'h6b;        memory[3182] <=  8'h73;        memory[3183] <=  8'h68;        memory[3184] <=  8'h63;        memory[3185] <=  8'h66;        memory[3186] <=  8'h69;        memory[3187] <=  8'h77;        memory[3188] <=  8'h68;        memory[3189] <=  8'h61;        memory[3190] <=  8'h74;        memory[3191] <=  8'h61;        memory[3192] <=  8'h6e;        memory[3193] <=  8'h61;        memory[3194] <=  8'h62;        memory[3195] <=  8'h61;        memory[3196] <=  8'h63;        memory[3197] <=  8'h61;        memory[3198] <=  8'h74;        memory[3199] <=  8'h61;        memory[3200] <=  8'h62;        memory[3201] <=  8'h61;        memory[3202] <=  8'h72;        memory[3203] <=  8'h63;        memory[3204] <=  8'h61;        memory[3205] <=  8'h68;        memory[3206] <=  8'h64;        memory[3207] <=  8'h75;        memory[3208] <=  8'h63;        memory[3209] <=  8'h74;        memory[3210] <=  8'h61;        memory[3211] <=  8'h64;        memory[3212] <=  8'h61;        memory[3213] <=  8'h61;        memory[3214] <=  8'h63;        memory[3215] <=  8'h61;        memory[3216] <=  8'h72;        memory[3217] <=  8'h63;        memory[3218] <=  8'h74;        memory[3219] <=  8'h72;        memory[3220] <=  8'h63;        memory[3221] <=  8'h61;        memory[3222] <=  8'h74;        memory[3223] <=  8'h72;        memory[3224] <=  8'h63;        memory[3225] <=  8'h61;        memory[3226] <=  8'h74;        memory[3227] <=  8'h63;        memory[3228] <=  8'h62;        memory[3229] <=  8'h61;        memory[3230] <=  8'h74;        memory[3231] <=  8'h62;        memory[3232] <=  8'h72;        memory[3233] <=  8'h63;        memory[3234] <=  8'h61;        memory[3235] <=  8'h74;        memory[3236] <=  8'h72;        memory[3237] <=  8'h6e;        memory[3238] <=  8'h62;        memory[3239] <=  8'h61;        memory[3240] <=  8'h63;        memory[3241] <=  8'h61;        memory[3242] <=  8'h74;        memory[3243] <=  8'h79;        memory[3244] <=  8'h73;        memory[3245] <=  8'h6e;        memory[3246] <=  8'h63;        memory[3247] <=  8'h74;        memory[3248] <=  8'h61;        memory[3249] <=  8'h6e;        memory[3250] <=  8'h62;        memory[3251] <=  8'h61;        memory[3252] <=  8'h63;        memory[3253] <=  8'h72;        memory[3254] <=  8'h6e;        memory[3255] <=  8'h74;        memory[3256] <=  8'h61;        memory[3257] <=  8'h62;        memory[3258] <=  8'h74;        memory[3259] <=  8'h6e;        memory[3260] <=  8'h61;        memory[3261] <=  8'h72;        memory[3262] <=  8'h62;        memory[3263] <=  8'h78;        memory[3264] <=  8'h74;        memory[3265] <=  8'h61;        memory[3266] <=  8'h72;        memory[3267] <=  8'h62;        memory[3268] <=  8'h61;        memory[3269] <=  8'h72;        memory[3270] <=  8'h74;        memory[3271] <=  8'h74;        memory[3272] <=  8'h62;        memory[3273] <=  8'h61;        memory[3274] <=  8'h72;        memory[3275] <=  8'h74;        memory[3276] <=  8'h78;        memory[3277] <=  8'h61;        memory[3278] <=  8'h74;        memory[3279] <=  8'h6b;        memory[3280] <=  8'h73;        memory[3281] <=  8'h68;        memory[3282] <=  8'h63;        memory[3283] <=  8'h66;        memory[3284] <=  8'h69;        memory[3285] <=  8'h77;        memory[3286] <=  8'h68;        memory[3287] <=  8'h61;        memory[3288] <=  8'h74;        memory[3289] <=  8'h61;        memory[3290] <=  8'h6e;        memory[3291] <=  8'h61;        memory[3292] <=  8'h62;        memory[3293] <=  8'h61;        memory[3294] <=  8'h63;        memory[3295] <=  8'h61;        memory[3296] <=  8'h74;        memory[3297] <=  8'h61;        memory[3298] <=  8'h62;        memory[3299] <=  8'h61;        memory[3300] <=  8'h72;        memory[3301] <=  8'h63;        memory[3302] <=  8'h61;        memory[3303] <=  8'h68;        memory[3304] <=  8'h64;        memory[3305] <=  8'h75;        memory[3306] <=  8'h63;        memory[3307] <=  8'h74;        memory[3308] <=  8'h61;        memory[3309] <=  8'h64;        memory[3310] <=  8'h61;        memory[3311] <=  8'h61;        memory[3312] <=  8'h63;        memory[3313] <=  8'h61;        memory[3314] <=  8'h72;        memory[3315] <=  8'h63;        memory[3316] <=  8'h74;        memory[3317] <=  8'h72;        memory[3318] <=  8'h63;        memory[3319] <=  8'h61;        memory[3320] <=  8'h74;        memory[3321] <=  8'h72;        memory[3322] <=  8'h63;        memory[3323] <=  8'h61;        memory[3324] <=  8'h74;        memory[3325] <=  8'h63;        memory[3326] <=  8'h62;        memory[3327] <=  8'h61;        memory[3328] <=  8'h74;        memory[3329] <=  8'h62;        memory[3330] <=  8'h72;        memory[3331] <=  8'h63;        memory[3332] <=  8'h61;        memory[3333] <=  8'h74;        memory[3334] <=  8'h72;        memory[3335] <=  8'h6e;        memory[3336] <=  8'h62;        memory[3337] <=  8'h61;        memory[3338] <=  8'h63;        memory[3339] <=  8'h61;        memory[3340] <=  8'h74;        memory[3341] <=  8'h79;        memory[3342] <=  8'h73;        memory[3343] <=  8'h6e;        memory[3344] <=  8'h63;        memory[3345] <=  8'h74;        memory[3346] <=  8'h61;        memory[3347] <=  8'h6e;        memory[3348] <=  8'h62;        memory[3349] <=  8'h61;        memory[3350] <=  8'h63;        memory[3351] <=  8'h72;        memory[3352] <=  8'h6e;        memory[3353] <=  8'h74;        memory[3354] <=  8'h61;        memory[3355] <=  8'h62;        memory[3356] <=  8'h74;        memory[3357] <=  8'h6e;        memory[3358] <=  8'h61;        memory[3359] <=  8'h72;        memory[3360] <=  8'h62;        memory[3361] <=  8'h78;        memory[3362] <=  8'h74;        memory[3363] <=  8'h61;        memory[3364] <=  8'h72;        memory[3365] <=  8'h64;        memory[3366] <=  8'h66;        memory[3367] <=  8'h73;        memory[3368] <=  8'h67;        memory[3369] <=  8'h76;        memory[3370] <=  8'h68;        memory[3371] <=  8'h62;        memory[3372] <=  8'h6b;        memory[3373] <=  8'h6a;        memory[3374] <=  8'h6e;        memory[3375] <=  8'h6d;        memory[3376] <=  8'h62;        memory[3377] <=  8'h76;        memory[3378] <=  8'h78;        memory[3379] <=  8'h63;        memory[3380] <=  8'h73;        memory[3381] <=  8'h66;        memory[3382] <=  8'h72;        memory[3383] <=  8'h74;        memory[3384] <=  8'h79;        memory[3385] <=  8'h75;        memory[3386] <=  8'h6a;        memory[3387] <=  8'h6e;        memory[3388] <=  8'h62;        memory[3389] <=  8'h76;        memory[3390] <=  8'h63;        memory[3391] <=  8'h64;        memory[3392] <=  8'h74;        memory[3393] <=  8'h79;        memory[3394] <=  8'h75;        memory[3395] <=  8'h69;        memory[3396] <=  8'h6b;        memory[3397] <=  8'h6d;        memory[3398] <=  8'h6e;        memory[3399] <=  8'h62;        memory[3400] <=  8'h76;        memory[3401] <=  8'h63;        memory[3402] <=  8'h78;        memory[3403] <=  8'h73;        memory[3404] <=  8'h64;        memory[3405] <=  8'h72;        memory[3406] <=  8'h74;        memory[3407] <=  8'h79;        memory[3408] <=  8'h75;        memory[3409] <=  8'h69;        memory[3410] <=  8'h6b;        memory[3411] <=  8'h6d;        memory[3412] <=  8'h6e;        memory[3413] <=  8'h62;        memory[3414] <=  8'h76;        memory[3415] <=  8'h63;        memory[3416] <=  8'h73;        memory[3417] <=  8'h77;        memory[3418] <=  8'h33;        memory[3419] <=  8'h34;        memory[3420] <=  8'h35;        memory[3421] <=  8'h36;        memory[3422] <=  8'h37;        memory[3423] <=  8'h38;        memory[3424] <=  8'h69;        memory[3425] <=  8'h6b;        memory[3426] <=  8'h6d;        memory[3427] <=  8'h6e;        memory[3428] <=  8'h62;        memory[3429] <=  8'h76;        memory[3430] <=  8'h63;        memory[3431] <=  8'h64;        memory[3432] <=  8'h65;        memory[3433] <=  8'h72;        memory[3434] <=  8'h36;        memory[3435] <=  8'h37;        memory[3436] <=  8'h38;        memory[3437] <=  8'h69;        memory[3438] <=  8'h6f;        memory[3439] <=  8'h6b;        memory[3440] <=  8'h6a;        memory[3441] <=  8'h6e;        memory[3442] <=  8'h62;        memory[3443] <=  8'h76;        memory[3444] <=  8'h63;        memory[3445] <=  8'h64;        memory[3446] <=  8'h72;        memory[3447] <=  8'h74;        memory[3448] <=  8'h79;        memory[3449] <=  8'h75;        memory[3450] <=  8'h73;        memory[3451] <=  8'h6a;        memory[3452] <=  8'h63;        memory[3453] <=  8'h6e;        memory[3454] <=  8'h62;        memory[3455] <=  8'h64;        memory[3456] <=  8'h66;        memory[3457] <=  8'h73;        memory[3458] <=  8'h74;        memory[3459] <=  8'h79;        memory[3460] <=  8'h75;        memory[3461] <=  8'h61;        memory[3462] <=  8'h69;        memory[3463] <=  8'h6b;        memory[3464] <=  8'h78;        memory[3465] <=  8'h6d;        memory[3466] <=  8'h6e;        memory[3467] <=  8'h73;        memory[3468] <=  8'h6a;        memory[3469] <=  8'h6f;        memory[3470] <=  8'h64;        memory[3471] <=  8'h6c;        memory[3472] <=  8'h63;        memory[3473] <=  8'h78;        memory[3474] <=  8'h62;        memory[3475] <=  8'h61;        memory[3476] <=  8'h72;        memory[3477] <=  8'h74;        memory[3478] <=  8'h78;        memory[3479] <=  8'h61;        memory[3480] <=  8'h74;        memory[3481] <=  8'h6b;        memory[3482] <=  8'h73;        memory[3483] <=  8'h68;        memory[3484] <=  8'h63;        memory[3485] <=  8'h66;        memory[3486] <=  8'h69;        memory[3487] <=  8'h77;        memory[3488] <=  8'h68;        memory[3489] <=  8'h61;        memory[3490] <=  8'h74;        memory[3491] <=  8'h61;        memory[3492] <=  8'h6e;        memory[3493] <=  8'h61;        memory[3494] <=  8'h62;        memory[3495] <=  8'h61;        memory[3496] <=  8'h63;        memory[3497] <=  8'h61;        memory[3498] <=  8'h74;        memory[3499] <=  8'h61;        memory[3500] <=  8'h62;        memory[3501] <=  8'h61;        memory[3502] <=  8'h72;        memory[3503] <=  8'h63;        memory[3504] <=  8'h61;        memory[3505] <=  8'h68;        memory[3506] <=  8'h64;        memory[3507] <=  8'h75;        memory[3508] <=  8'h63;        memory[3509] <=  8'h74;        memory[3510] <=  8'h61;        memory[3511] <=  8'h64;        memory[3512] <=  8'h61;        memory[3513] <=  8'h61;        memory[3514] <=  8'h63;        memory[3515] <=  8'h61;        memory[3516] <=  8'h72;        memory[3517] <=  8'h62;        memory[3518] <=  8'h61;        memory[3519] <=  8'h72;        memory[3520] <=  8'h74;        memory[3521] <=  8'h78;        memory[3522] <=  8'h61;        memory[3523] <=  8'h74;        memory[3524] <=  8'h6b;        memory[3525] <=  8'h73;        memory[3526] <=  8'h68;        memory[3527] <=  8'h63;        memory[3528] <=  8'h66;        memory[3529] <=  8'h69;        memory[3530] <=  8'h77;        memory[3531] <=  8'h68;        memory[3532] <=  8'h61;        memory[3533] <=  8'h74;        memory[3534] <=  8'h61;        memory[3535] <=  8'h6e;        memory[3536] <=  8'h61;        memory[3537] <=  8'h62;        memory[3538] <=  8'h61;        memory[3539] <=  8'h63;        memory[3540] <=  8'h61;        memory[3541] <=  8'h74;        memory[3542] <=  8'h61;        memory[3543] <=  8'h62;        memory[3544] <=  8'h61;        memory[3545] <=  8'h72;        memory[3546] <=  8'h63;        memory[3547] <=  8'h61;        memory[3548] <=  8'h68;        memory[3549] <=  8'h64;        memory[3550] <=  8'h75;        memory[3551] <=  8'h63;        memory[3552] <=  8'h74;        memory[3553] <=  8'h61;        memory[3554] <=  8'h64;        memory[3555] <=  8'h61;        memory[3556] <=  8'h61;        memory[3557] <=  8'h63;        memory[3558] <=  8'h61;        memory[3559] <=  8'h72;        memory[3560] <=  8'h62;        memory[3561] <=  8'h61;        memory[3562] <=  8'h72;        memory[3563] <=  8'h74;        memory[3564] <=  8'h78;        memory[3565] <=  8'h61;        memory[3566] <=  8'h74;        memory[3567] <=  8'h6b;        memory[3568] <=  8'h73;        memory[3569] <=  8'h68;        memory[3570] <=  8'h63;        memory[3571] <=  8'h66;        memory[3572] <=  8'h69;        memory[3573] <=  8'h77;        memory[3574] <=  8'h68;        memory[3575] <=  8'h61;        memory[3576] <=  8'h74;        memory[3577] <=  8'h61;        memory[3578] <=  8'h6e;        memory[3579] <=  8'h61;        memory[3580] <=  8'h62;        memory[3581] <=  8'h61;        memory[3582] <=  8'h63;        memory[3583] <=  8'h61;        memory[3584] <=  8'h74;        memory[3585] <=  8'h61;        memory[3586] <=  8'h62;        memory[3587] <=  8'h61;        memory[3588] <=  8'h72;        memory[3589] <=  8'h63;        memory[3590] <=  8'h61;        memory[3591] <=  8'h68;        memory[3592] <=  8'h64;        memory[3593] <=  8'h75;        memory[3594] <=  8'h63;        memory[3595] <=  8'h74;        memory[3596] <=  8'h61;        memory[3597] <=  8'h64;        memory[3598] <=  8'h61;        memory[3599] <=  8'h61;        memory[3600] <=  8'h63;        memory[3601] <=  8'h61;        memory[3602] <=  8'h72;        memory[3603] <=  8'h62;        memory[3604] <=  8'h61;        memory[3605] <=  8'h72;        memory[3606] <=  8'h74;        memory[3607] <=  8'h78;        memory[3608] <=  8'h61;        memory[3609] <=  8'h74;        memory[3610] <=  8'h6b;        memory[3611] <=  8'h73;        memory[3612] <=  8'h68;        memory[3613] <=  8'h63;        memory[3614] <=  8'h66;        memory[3615] <=  8'h69;        memory[3616] <=  8'h77;        memory[3617] <=  8'h68;        memory[3618] <=  8'h61;        memory[3619] <=  8'h74;        memory[3620] <=  8'h61;        memory[3621] <=  8'h6e;        memory[3622] <=  8'h61;        memory[3623] <=  8'h62;        memory[3624] <=  8'h61;        memory[3625] <=  8'h63;        memory[3626] <=  8'h61;        memory[3627] <=  8'h74;        memory[3628] <=  8'h61;        memory[3629] <=  8'h62;        memory[3630] <=  8'h61;        memory[3631] <=  8'h72;        memory[3632] <=  8'h63;        memory[3633] <=  8'h61;        memory[3634] <=  8'h68;        memory[3635] <=  8'h64;        memory[3636] <=  8'h75;        memory[3637] <=  8'h63;        memory[3638] <=  8'h74;        memory[3639] <=  8'h61;        memory[3640] <=  8'h64;        memory[3641] <=  8'h61;        memory[3642] <=  8'h61;        memory[3643] <=  8'h63;        memory[3644] <=  8'h61;        memory[3645] <=  8'h72;        memory[3646] <=  8'h62;        memory[3647] <=  8'h61;        memory[3648] <=  8'h72;        memory[3649] <=  8'h74;        memory[3650] <=  8'h78;        memory[3651] <=  8'h61;        memory[3652] <=  8'h74;        memory[3653] <=  8'h6b;        memory[3654] <=  8'h73;        memory[3655] <=  8'h68;        memory[3656] <=  8'h63;        memory[3657] <=  8'h66;        memory[3658] <=  8'h69;        memory[3659] <=  8'h77;        memory[3660] <=  8'h68;        memory[3661] <=  8'h61;        memory[3662] <=  8'h74;        memory[3663] <=  8'h61;        memory[3664] <=  8'h6e;        memory[3665] <=  8'h61;        memory[3666] <=  8'h62;        memory[3667] <=  8'h61;        memory[3668] <=  8'h63;        memory[3669] <=  8'h61;        memory[3670] <=  8'h74;        memory[3671] <=  8'h61;        memory[3672] <=  8'h62;        memory[3673] <=  8'h61;        memory[3674] <=  8'h72;        memory[3675] <=  8'h63;        memory[3676] <=  8'h61;        memory[3677] <=  8'h68;        memory[3678] <=  8'h64;        memory[3679] <=  8'h75;        memory[3680] <=  8'h63;        memory[3681] <=  8'h74;        memory[3682] <=  8'h61;        memory[3683] <=  8'h64;        memory[3684] <=  8'h61;        memory[3685] <=  8'h61;        memory[3686] <=  8'h63;        memory[3687] <=  8'h61;        memory[3688] <=  8'h72;        memory[3689] <=  8'h62;        memory[3690] <=  8'h61;        memory[3691] <=  8'h72;        memory[3692] <=  8'h74;        memory[3693] <=  8'h78;        memory[3694] <=  8'h61;        memory[3695] <=  8'h74;        memory[3696] <=  8'h6b;        memory[3697] <=  8'h73;        memory[3698] <=  8'h68;        memory[3699] <=  8'h63;        memory[3700] <=  8'h66;        memory[3701] <=  8'h69;        memory[3702] <=  8'h77;        memory[3703] <=  8'h68;        memory[3704] <=  8'h61;        memory[3705] <=  8'h74;        memory[3706] <=  8'h61;        memory[3707] <=  8'h6e;        memory[3708] <=  8'h61;        memory[3709] <=  8'h62;        memory[3710] <=  8'h61;        memory[3711] <=  8'h63;        memory[3712] <=  8'h61;        memory[3713] <=  8'h74;        memory[3714] <=  8'h61;        memory[3715] <=  8'h62;        memory[3716] <=  8'h61;        memory[3717] <=  8'h72;        memory[3718] <=  8'h63;        memory[3719] <=  8'h61;        memory[3720] <=  8'h68;        memory[3721] <=  8'h64;        memory[3722] <=  8'h75;        memory[3723] <=  8'h63;        memory[3724] <=  8'h74;        memory[3725] <=  8'h61;        memory[3726] <=  8'h64;        memory[3727] <=  8'h61;        memory[3728] <=  8'h61;        memory[3729] <=  8'h63;        memory[3730] <=  8'h61;        memory[3731] <=  8'h72;        memory[3732] <=  8'h62;        memory[3733] <=  8'h61;        memory[3734] <=  8'h72;        memory[3735] <=  8'h74;        memory[3736] <=  8'h78;        memory[3737] <=  8'h61;        memory[3738] <=  8'h74;        memory[3739] <=  8'h6b;        memory[3740] <=  8'h73;        memory[3741] <=  8'h68;        memory[3742] <=  8'h63;        memory[3743] <=  8'h66;        memory[3744] <=  8'h69;        memory[3745] <=  8'h77;        memory[3746] <=  8'h68;        memory[3747] <=  8'h61;        memory[3748] <=  8'h74;        memory[3749] <=  8'h61;        memory[3750] <=  8'h6e;        memory[3751] <=  8'h61;        memory[3752] <=  8'h62;        memory[3753] <=  8'h61;        memory[3754] <=  8'h63;        memory[3755] <=  8'h61;        memory[3756] <=  8'h74;        memory[3757] <=  8'h61;        memory[3758] <=  8'h62;        memory[3759] <=  8'h61;        memory[3760] <=  8'h72;        memory[3761] <=  8'h63;        memory[3762] <=  8'h61;        memory[3763] <=  8'h68;        memory[3764] <=  8'h64;        memory[3765] <=  8'h75;        memory[3766] <=  8'h63;        memory[3767] <=  8'h74;        memory[3768] <=  8'h61;        memory[3769] <=  8'h64;        memory[3770] <=  8'h61;        memory[3771] <=  8'h61;        memory[3772] <=  8'h63;        memory[3773] <=  8'h61;        memory[3774] <=  8'h72;        memory[3775] <=  8'h62;        memory[3776] <=  8'h61;        memory[3777] <=  8'h72;        memory[3778] <=  8'h74;        memory[3779] <=  8'h78;        memory[3780] <=  8'h61;        memory[3781] <=  8'h74;        memory[3782] <=  8'h6b;        memory[3783] <=  8'h73;        memory[3784] <=  8'h68;        memory[3785] <=  8'h63;        memory[3786] <=  8'h66;        memory[3787] <=  8'h69;        memory[3788] <=  8'h77;        memory[3789] <=  8'h68;        memory[3790] <=  8'h61;        memory[3791] <=  8'h74;        memory[3792] <=  8'h61;        memory[3793] <=  8'h6e;        memory[3794] <=  8'h61;        memory[3795] <=  8'h62;        memory[3796] <=  8'h61;        memory[3797] <=  8'h63;        memory[3798] <=  8'h61;        memory[3799] <=  8'h74;        memory[3800] <=  8'h61;        memory[3801] <=  8'h62;        memory[3802] <=  8'h61;        memory[3803] <=  8'h72;        memory[3804] <=  8'h63;        memory[3805] <=  8'h61;        memory[3806] <=  8'h68;        memory[3807] <=  8'h64;        memory[3808] <=  8'h75;        memory[3809] <=  8'h63;        memory[3810] <=  8'h74;        memory[3811] <=  8'h61;        memory[3812] <=  8'h64;        memory[3813] <=  8'h61;        memory[3814] <=  8'h61;        memory[3815] <=  8'h63;        memory[3816] <=  8'h61;        memory[3817] <=  8'h72;        memory[3818] <=  8'h62;        memory[3819] <=  8'h61;        memory[3820] <=  8'h72;        memory[3821] <=  8'h74;        memory[3822] <=  8'h78;        memory[3823] <=  8'h61;        memory[3824] <=  8'h74;        memory[3825] <=  8'h6b;        memory[3826] <=  8'h73;        memory[3827] <=  8'h68;        memory[3828] <=  8'h63;        memory[3829] <=  8'h66;        memory[3830] <=  8'h69;        memory[3831] <=  8'h77;        memory[3832] <=  8'h68;        memory[3833] <=  8'h61;        memory[3834] <=  8'h74;        memory[3835] <=  8'h61;        memory[3836] <=  8'h6e;        memory[3837] <=  8'h61;        memory[3838] <=  8'h62;        memory[3839] <=  8'h61;        memory[3840] <=  8'h63;        memory[3841] <=  8'h61;        memory[3842] <=  8'h74;        memory[3843] <=  8'h61;        memory[3844] <=  8'h62;        memory[3845] <=  8'h61;        memory[3846] <=  8'h72;        memory[3847] <=  8'h63;        memory[3848] <=  8'h61;        memory[3849] <=  8'h68;        memory[3850] <=  8'h64;        memory[3851] <=  8'h75;        memory[3852] <=  8'h63;        memory[3853] <=  8'h74;        memory[3854] <=  8'h61;        memory[3855] <=  8'h64;        memory[3856] <=  8'h61;        memory[3857] <=  8'h61;        memory[3858] <=  8'h63;        memory[3859] <=  8'h61;        memory[3860] <=  8'h72;        memory[3861] <=  8'h62;        memory[3862] <=  8'h61;        memory[3863] <=  8'h72;        memory[3864] <=  8'h74;        memory[3865] <=  8'h74;        memory[3866] <=  8'h62;        memory[3867] <=  8'h61;        memory[3868] <=  8'h72;        memory[3869] <=  8'h74;        memory[3870] <=  8'h78;        memory[3871] <=  8'h61;        memory[3872] <=  8'h74;        memory[3873] <=  8'h6b;        memory[3874] <=  8'h73;        memory[3875] <=  8'h68;        memory[3876] <=  8'h63;        memory[3877] <=  8'h66;        memory[3878] <=  8'h69;        memory[3879] <=  8'h77;        memory[3880] <=  8'h68;        memory[3881] <=  8'h61;        memory[3882] <=  8'h74;        memory[3883] <=  8'h61;        memory[3884] <=  8'h6e;        memory[3885] <=  8'h61;        memory[3886] <=  8'h62;        memory[3887] <=  8'h61;        memory[3888] <=  8'h63;        memory[3889] <=  8'h61;        memory[3890] <=  8'h74;        memory[3891] <=  8'h61;        memory[3892] <=  8'h62;        memory[3893] <=  8'h61;        memory[3894] <=  8'h72;        memory[3895] <=  8'h63;        memory[3896] <=  8'h61;        memory[3897] <=  8'h68;        memory[3898] <=  8'h64;        memory[3899] <=  8'h75;        memory[3900] <=  8'h63;        memory[3901] <=  8'h74;        memory[3902] <=  8'h61;        memory[3903] <=  8'h64;        memory[3904] <=  8'h61;        memory[3905] <=  8'h61;        memory[3906] <=  8'h63;        memory[3907] <=  8'h61;        memory[3908] <=  8'h72;        memory[3909] <=  8'h63;        memory[3910] <=  8'h74;        memory[3911] <=  8'h72;        memory[3912] <=  8'h63;        memory[3913] <=  8'h61;        memory[3914] <=  8'h74;        memory[3915] <=  8'h72;        memory[3916] <=  8'h63;        memory[3917] <=  8'h61;        memory[3918] <=  8'h74;        memory[3919] <=  8'h63;        memory[3920] <=  8'h62;        memory[3921] <=  8'h61;        memory[3922] <=  8'h74;        memory[3923] <=  8'h62;        memory[3924] <=  8'h72;        memory[3925] <=  8'h63;        memory[3926] <=  8'h61;        memory[3927] <=  8'h72;        memory[3928] <=  8'h62;        memory[3929] <=  8'h78;        memory[3930] <=  8'h74;        memory[3931] <=  8'h61;        memory[3932] <=  8'h72;        memory[3933] <=  8'h64;        memory[3934] <=  8'h66;        memory[3935] <=  8'h73;        memory[3936] <=  8'h67;        memory[3937] <=  8'h76;        memory[3938] <=  8'h68;        memory[3939] <=  8'h62;        memory[3940] <=  8'h6b;        memory[3941] <=  8'h6a;        memory[3942] <=  8'h6e;        memory[3943] <=  8'h6d;        memory[3944] <=  8'h62;        memory[3945] <=  8'h76;        memory[3946] <=  8'h78;        memory[3947] <=  8'h63;        memory[3948] <=  8'h73;        memory[3949] <=  8'h66;        memory[3950] <=  8'h72;        memory[3951] <=  8'h74;        memory[3952] <=  8'h79;        memory[3953] <=  8'h75;        memory[3954] <=  8'h6a;        memory[3955] <=  8'h6e;        memory[3956] <=  8'h62;        memory[3957] <=  8'h76;        memory[3958] <=  8'h63;        memory[3959] <=  8'h64;        memory[3960] <=  8'h74;        memory[3961] <=  8'h79;        memory[3962] <=  8'h75;        memory[3963] <=  8'h69;        memory[3964] <=  8'h6b;        memory[3965] <=  8'h6d;        memory[3966] <=  8'h6e;        memory[3967] <=  8'h62;        memory[3968] <=  8'h76;        memory[3969] <=  8'h63;        memory[3970] <=  8'h78;        memory[3971] <=  8'h73;        memory[3972] <=  8'h64;        memory[3973] <=  8'h72;        memory[3974] <=  8'h74;        memory[3975] <=  8'h79;        memory[3976] <=  8'h75;        memory[3977] <=  8'h69;        memory[3978] <=  8'h6b;        memory[3979] <=  8'h6d;        memory[3980] <=  8'h6e;        memory[3981] <=  8'h62;        memory[3982] <=  8'h76;        memory[3983] <=  8'h63;        memory[3984] <=  8'h73;        memory[3985] <=  8'h77;        memory[3986] <=  8'h33;        memory[3987] <=  8'h34;        memory[3988] <=  8'h35;        memory[3989] <=  8'h36;        memory[3990] <=  8'h37;        memory[3991] <=  8'h38;        memory[3992] <=  8'h69;        memory[3993] <=  8'h6b;        memory[3994] <=  8'h6d;        memory[3995] <=  8'h6e;        memory[3996] <=  8'h62;        memory[3997] <=  8'h76;        memory[3998] <=  8'h63;        memory[3999] <=  8'h64;        memory[4000] <=  8'h65;        memory[4001] <=  8'h72;        memory[4002] <=  8'h36;        memory[4003] <=  8'h37;        memory[4004] <=  8'h38;        memory[4005] <=  8'h69;        memory[4006] <=  8'h6f;        memory[4007] <=  8'h6b;        memory[4008] <=  8'h6a;        memory[4009] <=  8'h6e;        memory[4010] <=  8'h62;        memory[4011] <=  8'h76;        memory[4012] <=  8'h63;        memory[4013] <=  8'h64;        memory[4014] <=  8'h72;        memory[4015] <=  8'h74;        memory[4016] <=  8'h79;        memory[4017] <=  8'h75;        memory[4018] <=  8'h73;        memory[4019] <=  8'h6a;        memory[4020] <=  8'h63;        memory[4021] <=  8'h6e;        memory[4022] <=  8'h62;        memory[4023] <=  8'h64;        memory[4024] <=  8'h66;        memory[4025] <=  8'h73;        memory[4026] <=  8'h74;        memory[4027] <=  8'h79;        memory[4028] <=  8'h75;        memory[4029] <=  8'h61;        memory[4030] <=  8'h69;        memory[4031] <=  8'h6b;        memory[4032] <=  8'h78;        memory[4033] <=  8'h6d;        memory[4034] <=  8'h6e;        memory[4035] <=  8'h73;        memory[4036] <=  8'h6a;        memory[4037] <=  8'h6f;        memory[4038] <=  8'h64;        memory[4039] <=  8'h6c;        memory[4040] <=  8'h63;        memory[4041] <=  8'h78;        memory[4042] <=  8'h2c;        memory[4043] <=  8'h6d;        memory[4044] <=  8'h73;        memory[4045] <=  8'h6b;        memory[4046] <=  8'h64;        memory[4047] <=  8'h6c;        memory[4048] <=  8'h70;        memory[4049] <=  8'h5b;        memory[4050] <=  8'h3b;        memory[4051] <=  8'h73;        memory[4052] <=  8'h6c;        memory[4053] <=  8'h64;        memory[4054] <=  8'h70;        memory[4055] <=  8'h76;        memory[4056] <=  8'h63;        memory[4057] <=  8'h5b;        memory[4058] <=  8'h78;        memory[4059] <=  8'h76;        memory[4060] <=  8'h63;        memory[4061] <=  8'h5b;        memory[4062] <=  8'h78;        memory[4063] <=  8'h70;        memory[4064] <=  8'h6f;        memory[4065] <=  8'h20;        memory[4066] <=  8'h62;        memory[4067] <=  8'h61;        memory[4068] <=  8'h72;        memory[4069] <=  8'h74;        memory[4070] <=  8'h74;        memory[4071] <=  8'h62;        memory[4072] <=  8'h61;        memory[4073] <=  8'h72;        memory[4074] <=  8'h74;        memory[4075] <=  8'h78;        memory[4076] <=  8'h61;        memory[4077] <=  8'h74;        memory[4078] <=  8'h6b;        memory[4079] <=  8'h73;        memory[4080] <=  8'h68;        memory[4081] <=  8'h63;        memory[4082] <=  8'h66;        memory[4083] <=  8'h69;        memory[4084] <=  8'h77;        memory[4085] <=  8'h68;        memory[4086] <=  8'h61;        memory[4087] <=  8'h69;        memory[4088] <=  8'h6a;        memory[4089] <=  8'h78;        memory[4090] <=  8'h5d;        memory[4091] <=  8'h65;        memory[4092] <=  8'h6b;        memory[4093] <=  8'h6f;        memory[4094] <=  8'h39;        memory[4095] <=  8'h64;        memory[4096] <=  8'h75;        memory[4097] <=  8'h38;        memory[4098] <=  8'h79;        memory[4099] <=  8'h20;        memory[4100] <=  8'h37;        memory[4101] <=  8'h63;        memory[4102] <=  8'h67;        memory[4103] <=  8'h78;        memory[4104] <=  8'h63;        memory[4105] <=  8'h75;        memory[4106] <=  8'h68;        memory[4107] <=  8'h69;        memory[4108] <=  8'h6a;        memory[4109] <=  8'h77;        memory[4110] <=  8'h69;        memory[4111] <=  8'h64;        memory[4112] <=  8'h66;        memory[4113] <=  8'h68;        memory[4114] <=  8'h75;        memory[4115] <=  8'h76;        memory[4116] <=  8'h64;        memory[4117] <=  8'h62;        memory[4118] <=  8'h66;        memory[4119] <=  8'h6a;        memory[4120] <=  8'h6e;        memory[4121] <=  8'h6b;        memory[4122] <=  8'h6a;        memory[4123] <=  8'h65;        memory[4124] <=  8'h38;        memory[4125] <=  8'h66;        memory[4126] <=  8'h37;        memory[4127] <=  8'h67;        memory[4128] <=  8'h79;        memory[4129] <=  8'h76;        memory[4130] <=  8'h63;        memory[4131] <=  8'h68;        memory[4132] <=  8'h69;        memory[4133] <=  8'h6a;        memory[4134] <=  8'h33;        memory[4135] <=  8'h65;        memory[4136] <=  8'h67;        memory[4137] <=  8'h79;        memory[4138] <=  8'h72;        memory[4139] <=  8'h64;        memory[4140] <=  8'h62;        memory[4141] <=  8'h6e;        memory[4142] <=  8'h63;        memory[4143] <=  8'h7a;        memory[4144] <=  8'h6a;        memory[4145] <=  8'h6f;        memory[4146] <=  8'h66;        memory[4147] <=  8'h78;        memory[4148] <=  8'h6a;        memory[4149] <=  8'h69;        memory[4150] <=  8'h63;        memory[4151] <=  8'h68;        memory[4152] <=  8'h62;        memory[4153] <=  8'h6e;        memory[4154] <=  8'h6d;        memory[4155] <=  8'h63;        memory[4156] <=  8'h73;        memory[4157] <=  8'h6c;        memory[4158] <=  8'h6b;        memory[4159] <=  8'h6a;        memory[4160] <=  8'h69;        memory[4161] <=  8'h68;        memory[4162] <=  8'h76;        memory[4163] <=  8'h75;        memory[4164] <=  8'h69;        memory[4165] <=  8'h64;        memory[4166] <=  8'h68;        memory[4167] <=  8'h75;        memory[4168] <=  8'h67;        memory[4169] <=  8'h79;        memory[4170] <=  8'h62;        memory[4171] <=  8'h68;        memory[4172] <=  8'h65;        memory[4173] <=  8'h6a;        memory[4174] <=  8'h72;        memory[4175] <=  8'h6b;        memory[4176] <=  8'h6a;        memory[4177] <=  8'h6f;        memory[4178] <=  8'h64;        memory[4179] <=  8'h67;        memory[4180] <=  8'h69;        memory[4181] <=  8'h75;        memory[4182] <=  8'h69;        memory[4183] <=  8'h67;        memory[4184] <=  8'h76;        memory[4185] <=  8'h79;        memory[4186] <=  8'h75;        memory[4187] <=  8'h67;        memory[4188] <=  8'h78;        memory[4189] <=  8'h68;        memory[4190] <=  8'h63;        memory[4191] <=  8'h20;        memory[4192] <=  8'h20;        memory[4193] <=  8'h20;        memory[4194] <=  8'h78;        memory[4195] <=  8'h76;        memory[4196] <=  8'h20;        memory[4197] <=  8'h63;        memory[4198] <=  8'h78;        memory[4199] <=  8'h67;        memory[4200] <=  8'h79;        memory[4201] <=  8'h63;        memory[4202] <=  8'h75;        memory[4203] <=  8'h68;        memory[4204] <=  8'h6a;        memory[4205] <=  8'h6b;        memory[4206] <=  8'h61;        memory[4207] <=  8'h6c;        memory[4208] <=  8'h78;        memory[4209] <=  8'h76;        memory[4210] <=  8'h70;        memory[4211] <=  8'h6f;        memory[4212] <=  8'h69;        memory[4213] <=  8'h6a;        memory[4214] <=  8'h69;        memory[4215] <=  8'h68;        memory[4216] <=  8'h6a;        memory[4217] <=  8'h62;        memory[4218] <=  8'h77;        memory[4219] <=  8'h65;        memory[4220] <=  8'h6e;        memory[4221] <=  8'h61;        memory[4222] <=  8'h66;        memory[4223] <=  8'h6d;        memory[4224] <=  8'h64;        memory[4225] <=  8'h6b;        memory[4226] <=  8'h6d;        memory[4227] <=  8'h76;        memory[4228] <=  8'h6c;        memory[4229] <=  8'h63;        memory[4230] <=  8'h6f;        memory[4231] <=  8'h64;        memory[4232] <=  8'h69;        memory[4233] <=  8'h75;        memory[4234] <=  8'h68;        memory[4235] <=  8'h73;        memory[4236] <=  8'h66;        memory[4237] <=  8'h65;        memory[4238] <=  8'h62;        memory[4239] <=  8'h6e;        memory[4240] <=  8'h64;        memory[4241] <=  8'h73;        memory[4242] <=  8'h63;        memory[4243] <=  8'h6b;        memory[4244] <=  8'h20;        memory[4245] <=  8'h78;        memory[4246] <=  8'h6a;        memory[4247] <=  8'h78;        memory[4248] <=  8'h63;        memory[4249] <=  8'h73;        memory[4250] <=  8'h64;        memory[4251] <=  8'h66;        memory[4252] <=  8'h6b;        memory[4253] <=  8'h64;        memory[4254] <=  8'h6e;        memory[4255] <=  8'h6d;        memory[4256] <=  8'h64;        memory[4257] <=  8'h73;        memory[4258] <=  8'h63;        memory[4259] <=  8'h6b;        memory[4260] <=  8'h78;        memory[4261] <=  8'h6c;        memory[4262] <=  8'h6f;        memory[4263] <=  8'h66;        memory[4264] <=  8'h6a;        memory[4265] <=  8'h69;        memory[4266] <=  8'h61;        memory[4267] <=  8'h62;        memory[4268] <=  8'h6e;        memory[4269] <=  8'h20;        memory[4270] <=  8'h78;        memory[4271] <=  8'h6b;        memory[4272] <=  8'h6d;        memory[4273] <=  8'h20;        memory[4274] <=  8'h6f;        memory[4275] <=  8'h63;        memory[4276] <=  8'h76;        memory[4277] <=  8'h73;        memory[4278] <=  8'h64;        memory[4279] <=  8'h69;        memory[4280] <=  8'h66;        memory[4281] <=  8'h68;        memory[4282] <=  8'h65;        memory[4283] <=  8'h71;        memory[4284] <=  8'h6a;        memory[4285] <=  8'h77;        memory[4286] <=  8'h62;        memory[4287] <=  8'h65;        memory[4288] <=  8'h6e;        memory[4289] <=  8'h20;        memory[4290] <=  8'h6d;        memory[4291] <=  8'h64;        memory[4292] <=  8'h73;        memory[4293] <=  8'h6c;        memory[4294] <=  8'h76;        memory[4295] <=  8'h6b;        memory[4296] <=  8'h63;        memory[4297] <=  8'h78;        memory[4298] <=  8'h20;        memory[4299] <=  8'h6f;        memory[4300] <=  8'h78;        memory[4301] <=  8'h69;        memory[4302] <=  8'h63;        memory[4303] <=  8'h6a;        memory[4304] <=  8'h76;        memory[4305] <=  8'h64;        memory[4306] <=  8'h66;        memory[4307] <=  8'h65;        memory[4308] <=  8'h71;        memory[4309] <=  8'h6e;        memory[4310] <=  8'h20;        memory[4311] <=  8'h64;        memory[4312] <=  8'h6d;        memory[4313] <=  8'h73;        memory[4314] <=  8'h6c;        memory[4315] <=  8'h63;        memory[4316] <=  8'h78;        memory[4317] <=  8'h6b;        memory[4318] <=  8'h20;        memory[4319] <=  8'h6f;        memory[4320] <=  8'h78;        memory[4321] <=  8'h63;        memory[4322] <=  8'h76;        memory[4323] <=  8'h6a;        memory[4324] <=  8'h64;        memory[4325] <=  8'h62;        memory[4326] <=  8'h71;        memory[4327] <=  8'h77;        memory[4328] <=  8'h65;        memory[4329] <=  8'h6e;        memory[4330] <=  8'h6d;        memory[4331] <=  8'h64;        memory[4332] <=  8'h6c;        memory[4333] <=  8'h73;        memory[4334] <=  8'h2c;        memory[4335] <=  8'h76;        memory[4336] <=  8'h63;        memory[4337] <=  8'h78;        memory[4338] <=  8'h20;        memory[4339] <=  8'h63;        memory[4340] <=  8'h6f;        memory[4341] <=  8'h69;        memory[4342] <=  8'h76;        memory[4343] <=  8'h68;        memory[4344] <=  8'h73;        memory[4345] <=  8'h64;        memory[4346] <=  8'h62;        memory[4347] <=  8'h71;        memory[4348] <=  8'h77;        memory[4349] <=  8'h65;        memory[4350] <=  8'h6e;        memory[4351] <=  8'h64;        memory[4352] <=  8'h6b;        memory[4353] <=  8'h73;        memory[4354] <=  8'h76;        memory[4355] <=  8'h6f;        memory[4356] <=  8'h63;        memory[4357] <=  8'h20;        memory[4358] <=  8'h76;        memory[4359] <=  8'h69;        memory[4360] <=  8'h75;        memory[4361] <=  8'h69;        memory[4362] <=  8'h68;        memory[4363] <=  8'h63;        memory[4364] <=  8'h78;        memory[4365] <=  8'h69;        memory[4366] <=  8'h6f;        memory[4367] <=  8'h76;        memory[4368] <=  8'h73;        memory[4369] <=  8'h64;        memory[4370] <=  8'h61;        memory[4371] <=  8'h64;        memory[4372] <=  8'h6e;        memory[4373] <=  8'h77;        memory[4374] <=  8'h71;        memory[4375] <=  8'h6b;        memory[4376] <=  8'h6c;        memory[4377] <=  8'h73;        memory[4378] <=  8'h76;        memory[4379] <=  8'h6e;        memory[4380] <=  8'h62;        memory[4381] <=  8'h20;        memory[4382] <=  8'h64;        memory[4383] <=  8'h66;        memory[4384] <=  8'h6a;        memory[4385] <=  8'h6b;        memory[4386] <=  8'h71;        memory[4387] <=  8'h64;        memory[4388] <=  8'h77;        memory[4389] <=  8'h65;        memory[4390] <=  8'h6e;        memory[4391] <=  8'h62;        memory[4392] <=  8'h20;        memory[4393] <=  8'h64;        memory[4394] <=  8'h73;        memory[4395] <=  8'h76;        memory[4396] <=  8'h68;        memory[4397] <=  8'h64;        memory[4398] <=  8'h61;        memory[4399] <=  8'h71;        memory[4400] <=  8'h77;        memory[4401] <=  8'h6a;        memory[4402] <=  8'h65;        memory[4403] <=  8'h6e;        memory[4404] <=  8'h64;        memory[4405] <=  8'h20;        memory[4406] <=  8'h61;        memory[4407] <=  8'h63;        memory[4408] <=  8'h62;        memory[4409] <=  8'h68;        memory[4410] <=  8'h64;        memory[4411] <=  8'h61;        memory[4412] <=  8'h77;        memory[4413] <=  8'h71;        memory[4414] <=  8'h6e;        memory[4415] <=  8'h20;        memory[4416] <=  8'h62;        memory[4417] <=  8'h73;        memory[4418] <=  8'h76;        memory[4419] <=  8'h61;        memory[4420] <=  8'h67;        memory[4421] <=  8'h76;        memory[4422] <=  8'h68;        memory[4423] <=  8'h67;        memory[4424] <=  8'h61;        memory[4425] <=  8'h73;        memory[4426] <=  8'h6a;        memory[4427] <=  8'h6b;        memory[4428] <=  8'h63;        memory[4429] <=  8'h78;        memory[4430] <=  8'h76;        memory[4431] <=  8'h6e;        memory[4432] <=  8'h73;        memory[4433] <=  8'h64;        memory[4434] <=  8'h20;        memory[4435] <=  8'h66;        memory[4436] <=  8'h62;        memory[4437] <=  8'h64;        memory[4438] <=  8'h61;        memory[4439] <=  8'h73;        memory[4440] <=  8'h76;        memory[4441] <=  8'h67;        memory[4442] <=  8'h63;        memory[4443] <=  8'h79;        memory[4444] <=  8'h7a;        memory[4445] <=  8'h78;        memory[4446] <=  8'h79;        memory[4447] <=  8'h75;        memory[4448] <=  8'h20;        memory[4449] <=  8'h69;        memory[4450] <=  8'h6a;        memory[4451] <=  8'h64;        memory[4452] <=  8'h66;        memory[4453] <=  8'h6b;        memory[4454] <=  8'h61;        memory[4455] <=  8'h64;        memory[4456] <=  8'h63;        memory[4457] <=  8'h78;        memory[4458] <=  8'h68;        memory[4459] <=  8'h20;        memory[4460] <=  8'h67;        memory[4461] <=  8'h61;        memory[4462] <=  8'h68;        memory[4463] <=  8'h75;        memory[4464] <=  8'h64;        memory[4465] <=  8'h73;        memory[4466] <=  8'h69;        memory[4467] <=  8'h6a;        memory[4468] <=  8'h61;        memory[4469] <=  8'h6b;        memory[4470] <=  8'h63;        memory[4471] <=  8'h62;        memory[4472] <=  8'h61;        memory[4473] <=  8'h72;        memory[4474] <=  8'h73;        memory[4475] <=  8'h68;        memory[4476] <=  8'h64;        memory[4477] <=  8'h66;        memory[4478] <=  8'h67;        memory[4479] <=  8'h73;        memory[4480] <=  8'h68;        memory[4481] <=  8'h64;        memory[4482] <=  8'h66;        memory[4483] <=  8'h68;        memory[4484] <=  8'h64;        memory[4485] <=  8'h6a;        memory[4486] <=  8'h68;        memory[4487] <=  8'h62;        memory[4488] <=  8'h67;        memory[4489] <=  8'h63;        memory[4490] <=  8'h61;        memory[4491] <=  8'h66;        memory[4492] <=  8'h73;        memory[4493] <=  8'h79;        memory[4494] <=  8'h67;        memory[4495] <=  8'h6b;        memory[4496] <=  8'h75;        memory[4497] <=  8'h64;        memory[4498] <=  8'h68;        memory[4499] <=  8'h62;        memory[4500] <=  8'h77;        memory[4501] <=  8'h76;        memory[4502] <=  8'h67;        memory[4503] <=  8'h61;        memory[4504] <=  8'h66;        memory[4505] <=  8'h64;        memory[4506] <=  8'h74;        memory[4507] <=  8'h75;        memory[4508] <=  8'h66;        memory[4509] <=  8'h79;        memory[4510] <=  8'h67;        memory[4511] <=  8'h69;        memory[4512] <=  8'h75;        memory[4513] <=  8'h68;        memory[4514] <=  8'h6c;        memory[4515] <=  8'h6a;        memory[4516] <=  8'h62;        memory[4517] <=  8'h6b;        memory[4518] <=  8'h68;        memory[4519] <=  8'h76;        memory[4520] <=  8'h67;        memory[4521] <=  8'h63;        memory[4522] <=  8'h66;        memory[4523] <=  8'h78;        memory[4524] <=  8'h64;        memory[4525] <=  8'h74;        memory[4526] <=  8'h75;        memory[4527] <=  8'h79;        memory[4528] <=  8'h69;        memory[4529] <=  8'h75;        memory[4530] <=  8'h68;        memory[4531] <=  8'h6c;        memory[4532] <=  8'h6a;        memory[4533] <=  8'h6b;        memory[4534] <=  8'h67;        memory[4535] <=  8'h6a;        memory[4536] <=  8'h63;        memory[4537] <=  8'h66;        memory[4538] <=  8'h68;        memory[4539] <=  8'h64;        memory[4540] <=  8'h67;        memory[4541] <=  8'h72;        memory[4542] <=  8'h79;        memory[4543] <=  8'h74;        memory[4544] <=  8'h66;        memory[4545] <=  8'h75;        memory[4546] <=  8'h79;        memory[4547] <=  8'h69;        memory[4548] <=  8'h68;        memory[4549] <=  8'h6c;        memory[4550] <=  8'h62;        memory[4551] <=  8'h6d;        memory[4552] <=  8'h76;        memory[4553] <=  8'h6e;        memory[4554] <=  8'h63;        memory[4555] <=  8'h66;        memory[4556] <=  8'h68;        memory[4557] <=  8'h64;        memory[4558] <=  8'h74;        memory[4559] <=  8'h75;        memory[4560] <=  8'h67;        memory[4561] <=  8'h79;        memory[4562] <=  8'h69;        memory[4563] <=  8'h68;        memory[4564] <=  8'h75;        memory[4565] <=  8'h6a;        memory[4566] <=  8'h6c;        memory[4567] <=  8'h62;        memory[4568] <=  8'h6d;        memory[4569] <=  8'h76;        memory[4570] <=  8'h6e;        memory[4571] <=  8'h63;        memory[4572] <=  8'h66;        memory[4573] <=  8'h68;        memory[4574] <=  8'h67;        memory[4575] <=  8'h79;        memory[4576] <=  8'h68;        memory[4577] <=  8'h75;        memory[4578] <=  8'h6a;        memory[4579] <=  8'h6e;        memory[4580] <=  8'h2c;        memory[4581] <=  8'h62;        memory[4582] <=  8'h6e;        memory[4583] <=  8'h6d;        memory[4584] <=  8'h76;        memory[4585] <=  8'h6e;        memory[4586] <=  8'h63;        memory[4587] <=  8'h66;        memory[4588] <=  8'h68;        memory[4589] <=  8'h74;        memory[4590] <=  8'h79;        memory[4591] <=  8'h69;        memory[4592] <=  8'h75;        memory[4593] <=  8'h6c;        memory[4594] <=  8'h6a;        memory[4595] <=  8'h62;        memory[4596] <=  8'h6d;        memory[4597] <=  8'h76;        memory[4598] <=  8'h6e;        memory[4599] <=  8'h63;        memory[4600] <=  8'h66;        memory[4601] <=  8'h74;        memory[4602] <=  8'h75;        memory[4603] <=  8'h79;        memory[4604] <=  8'h69;        memory[4605] <=  8'h68;        memory[4606] <=  8'h6b;        memory[4607] <=  8'h62;        memory[4608] <=  8'h76;        memory[4609] <=  8'h63;        memory[4610] <=  8'h66;        memory[4611] <=  8'h67;        memory[4612] <=  8'h74;        memory[4613] <=  8'h75;        memory[4614] <=  8'h79;        memory[4615] <=  8'h69;        memory[4616] <=  8'h75;        memory[4617] <=  8'h68;        memory[4618] <=  8'h6a;        memory[4619] <=  8'h6b;        memory[4620] <=  8'h62;        memory[4621] <=  8'h76;        memory[4622] <=  8'h63;        memory[4623] <=  8'h66;        memory[4624] <=  8'h74;        memory[4625] <=  8'h75;        memory[4626] <=  8'h79;        memory[4627] <=  8'h69;        memory[4628] <=  8'h75;        memory[4629] <=  8'h6a;        memory[4630] <=  8'h6b;        memory[4631] <=  8'h6e;        memory[4632] <=  8'h62;        memory[4633] <=  8'h76;        memory[4634] <=  8'h67;        memory[4635] <=  8'h66;        memory[4636] <=  8'h74;        memory[4637] <=  8'h79;        memory[4638] <=  8'h75;        memory[4639] <=  8'h75;        memory[4640] <=  8'h69;        memory[4641] <=  8'h6a;        memory[4642] <=  8'h6b;        memory[4643] <=  8'h68;        memory[4644] <=  8'h62;        memory[4645] <=  8'h6a;        memory[4646] <=  8'h67;        memory[4647] <=  8'h68;        memory[4648] <=  8'h66;        memory[4649] <=  8'h79;        memory[4650] <=  8'h74;        memory[4651] <=  8'h79;        memory[4652] <=  8'h69;        memory[4653] <=  8'h75;        memory[4654] <=  8'h64;        memory[4655] <=  8'h6a;        memory[4656] <=  8'h6b;        memory[4657] <=  8'h68;        memory[4658] <=  8'h63;        memory[4659] <=  8'h7a;        memory[4660] <=  8'h67;        memory[4661] <=  8'h68;        memory[4662] <=  8'h74;        memory[4663] <=  8'h75;        memory[4664] <=  8'h79;        memory[4665] <=  8'h69;        memory[4666] <=  8'h61;        memory[4667] <=  8'h73;        memory[4668] <=  8'h75;        memory[4669] <=  8'h6a;        memory[4670] <=  8'h6b;        memory[4671] <=  8'h62;        memory[4672] <=  8'h6e;        memory[4673] <=  8'h61;        memory[4674] <=  8'h76;        memory[4675] <=  8'h63;        memory[4676] <=  8'h66;        memory[4677] <=  8'h68;        memory[4678] <=  8'h75;        memory[4679] <=  8'h61;        memory[4680] <=  8'h73;        memory[4681] <=  8'h79;        memory[4682] <=  8'h64;        memory[4683] <=  8'h75;        memory[4684] <=  8'h69;        memory[4685] <=  8'h6a;        memory[4686] <=  8'h61;        memory[4687] <=  8'h6b;        memory[4688] <=  8'h62;        memory[4689] <=  8'h63;        memory[4690] <=  8'h78;        memory[4691] <=  8'h68;        memory[4692] <=  8'h67;        memory[4693] <=  8'h79;        memory[4694] <=  8'h75;        memory[4695] <=  8'h7a;        memory[4696] <=  8'h63;        memory[4697] <=  8'h61;        memory[4698] <=  8'h73;        memory[4699] <=  8'h69;        memory[4700] <=  8'h75;        memory[4701] <=  8'h6f;        memory[4702] <=  8'h69;        memory[4703] <=  8'h6a;        memory[4704] <=  8'h61;        memory[4705] <=  8'h6c;        memory[4706] <=  8'h63;        memory[4707] <=  8'h78;        memory[4708] <=  8'h62;        memory[4709] <=  8'h63;        memory[4710] <=  8'h20;        memory[4711] <=  8'h6e;        memory[4712] <=  8'h76;        memory[4713] <=  8'h63;        memory[4714] <=  8'h61;        memory[4715] <=  8'h64;        memory[4716] <=  8'h73;        memory[4717] <=  8'h67;        memory[4718] <=  8'h79;        memory[4719] <=  8'h68;        memory[4720] <=  8'h75;        memory[4721] <=  8'h61;        memory[4722] <=  8'h6a;        memory[4723] <=  8'h6b;        memory[4724] <=  8'h78;        memory[4725] <=  8'h62;        memory[4726] <=  8'h20;        memory[4727] <=  8'h6e;        memory[4728] <=  8'h76;        memory[4729] <=  8'h63;        memory[4730] <=  8'h61;        memory[4731] <=  8'h73;        memory[4732] <=  8'h67;        memory[4733] <=  8'h68;        memory[4734] <=  8'h75;        memory[4735] <=  8'h6a;        memory[4736] <=  8'h6c;        memory[4737] <=  8'h6b;        memory[4738] <=  8'h63;        memory[4739] <=  8'h78;        memory[4740] <=  8'h20;        memory[4741] <=  8'h6a;        memory[4742] <=  8'h6b;        memory[4743] <=  8'h68;        memory[4744] <=  8'h61;        memory[4745] <=  8'h73;        memory[4746] <=  8'h76;        memory[4747] <=  8'h64;        memory[4748] <=  8'h6e;        memory[4749] <=  8'h20;        memory[4750] <=  8'h62;        memory[4751] <=  8'h6e;        memory[4752] <=  8'h6d;        memory[4753] <=  8'h6b;        memory[4754] <=  8'h77;        memory[4755] <=  8'h64;        memory[4756] <=  8'h6f;        memory[4757] <=  8'h77;        memory[4758] <=  8'h69;        memory[4759] <=  8'h6f;        memory[4760] <=  8'h75;        memory[4761] <=  8'h69;        memory[4762] <=  8'h68;        memory[4763] <=  8'h62;        memory[4764] <=  8'h6e;        memory[4765] <=  8'h6b;        memory[4766] <=  8'h77;        memory[4767] <=  8'h69;        memory[4768] <=  8'h6f;        memory[4769] <=  8'h75;        memory[4770] <=  8'h71;        memory[4771] <=  8'h69;        memory[4772] <=  8'h79;        memory[4773] <=  8'h67;        memory[4774] <=  8'h6a;        memory[4775] <=  8'h64;        memory[4776] <=  8'h61;        memory[4777] <=  8'h76;        memory[4778] <=  8'h62;        memory[4779] <=  8'h6e;        memory[4780] <=  8'h6b;        memory[4781] <=  8'h6f;        memory[4782] <=  8'h70;        memory[4783] <=  8'h64;        memory[4784] <=  8'h76;        memory[4785] <=  8'h69;        memory[4786] <=  8'h6f;        memory[4787] <=  8'h75;        memory[4788] <=  8'h69;        memory[4789] <=  8'h48;        memory[4790] <=  8'h42;        memory[4791] <=  8'h6b;        memory[4792] <=  8'h64;        memory[4793] <=  8'h6e;        memory[4794] <=  8'h6c;        memory[4795] <=  8'h71;        memory[4796] <=  8'h6b;        memory[4797] <=  8'h6d;        memory[4798] <=  8'h6a;        memory[4799] <=  8'h70;        memory[4800] <=  8'h69;        memory[4801] <=  8'h6f;        memory[4802] <=  8'h68;        memory[4803] <=  8'h65;        memory[4804] <=  8'h66;        memory[4805] <=  8'h75;        memory[4806] <=  8'h67;        memory[4807] <=  8'h69;        memory[4808] <=  8'h73;        memory[4809] <=  8'h61;        memory[4810] <=  8'h62;        memory[4811] <=  8'h64;        memory[4812] <=  8'h6b;        memory[4813] <=  8'h6a;        memory[4814] <=  8'h6b;        memory[4815] <=  8'h6c;        memory[4816] <=  8'h6a;        memory[4817] <=  8'h69;        memory[4818] <=  8'h73;        memory[4819] <=  8'h6f;        memory[4820] <=  8'h71;        memory[4821] <=  8'h68;        memory[4822] <=  8'h77;        memory[4823] <=  8'h67;        memory[4824] <=  8'h69;        memory[4825] <=  8'h79;        memory[4826] <=  8'h6a;        memory[4827] <=  8'h64;        memory[4828] <=  8'h76;        memory[4829] <=  8'h62;        memory[4830] <=  8'h6e;        memory[4831] <=  8'h61;        memory[4832] <=  8'h73;        memory[4833] <=  8'h66;        memory[4834] <=  8'h6c;        memory[4835] <=  8'h6b;        memory[4836] <=  8'h64;        memory[4837] <=  8'h6a;        memory[4838] <=  8'h68;        memory[4839] <=  8'h63;        memory[4840] <=  8'h67;        memory[4841] <=  8'h6a;        memory[4842] <=  8'h76;        memory[4843] <=  8'h73;        memory[4844] <=  8'h64;        memory[4845] <=  8'h62;        memory[4846] <=  8'h62;        memory[4847] <=  8'h61;        memory[4848] <=  8'h72;        memory[4849] <=  8'h62;        memory[4850] <=  8'h62;        memory[4851] <=  8'h73;        memory[4852] <=  8'h62;        memory[4853] <=  8'h67;        memory[4854] <=  8'h73;        memory[4855] <=  8'h66;        memory[4856] <=  8'h67;        memory[4857] <=  8'h61;        memory[4858] <=  8'h68;        memory[4859] <=  8'h66;        memory[4860] <=  8'h73;        memory[4861] <=  8'h68;        memory[4862] <=  8'h61;        memory[4863] <=  8'h66;        memory[4864] <=  8'h73;        memory[4865] <=  8'h66;        memory[4866] <=  8'h68;        memory[4867] <=  8'h61;        memory[4868] <=  8'h69;        memory[4869] <=  8'h64;        memory[4870] <=  8'h75;        memory[4871] <=  8'h67;        memory[4872] <=  8'h64;        memory[4873] <=  8'h77;        memory[4874] <=  8'h62;        memory[4875] <=  8'h61;        memory[4876] <=  8'h62;        memory[4877] <=  8'h72;        memory[4878] <=  8'h62;        memory[4879] <=  8'h61;        memory[4880] <=  8'h62;        memory[4881] <=  8'h62;        memory[4882] <=  8'h74;        memory[4883] <=  8'h62;        memory[4884] <=  8'h62;        memory[4885] <=  8'h62;        memory[4886] <=  8'h62;        memory[4887] <=  8'h62;        memory[4888] <=  8'h62;        memory[4889] <=  8'h62;        memory[4890] <=  8'h62;        memory[4891] <=  8'h61;        memory[4892] <=  8'h62;        memory[4893] <=  8'h62;        memory[4894] <=  8'h72;        memory[4895] <=  8'h74;        memory[4896] <=  8'h62;        memory[4897] <=  8'h62;        memory[4898] <=  8'h61;        memory[4899] <=  8'h62;        memory[4900] <=  8'h72;        memory[4901] <=  8'h62;        memory[4902] <=  8'h74;        memory[4903] <=  8'h62;        memory[4904] <=  8'h62;        memory[4905] <=  8'h62;        memory[4906] <=  8'h63;        memory[4907] <=  8'h61;        memory[4908] <=  8'h72;        memory[4909] <=  8'h74;        memory[4910] <=  8'h73;        memory[4911] <=  8'h62;        memory[4912] <=  8'h61;        memory[4913] <=  8'h72;        memory[4914] <=  8'h74;        memory[4915] <=  8'h74;        memory[4916] <=  8'h62;        memory[4917] <=  8'h61;        memory[4918] <=  8'h72;        memory[4919] <=  8'h74;        memory[4920] <=  8'h78;        memory[4921] <=  8'h61;        memory[4922] <=  8'h74;        memory[4923] <=  8'h6b;        memory[4924] <=  8'h73;        memory[4925] <=  8'h68;        memory[4926] <=  8'h63;        memory[4927] <=  8'h66;        memory[4928] <=  8'h69;        memory[4929] <=  8'h77;        memory[4930] <=  8'h68;        memory[4931] <=  8'h61;        memory[4932] <=  8'h74;        memory[4933] <=  8'h61;        memory[4934] <=  8'h6e;        memory[4935] <=  8'h61;        memory[4936] <=  8'h62;        memory[4937] <=  8'h61;        memory[4938] <=  8'h63;        memory[4939] <=  8'h61;        memory[4940] <=  8'h74;        memory[4941] <=  8'h61;        memory[4942] <=  8'h62;        memory[4943] <=  8'h61;        memory[4944] <=  8'h72;        memory[4945] <=  8'h63;        memory[4946] <=  8'h61;        memory[4947] <=  8'h68;        memory[4948] <=  8'h64;        memory[4949] <=  8'h75;        memory[4950] <=  8'h63;        memory[4951] <=  8'h74;        memory[4952] <=  8'h61;        memory[4953] <=  8'h64;        memory[4954] <=  8'h61;        memory[4955] <=  8'h61;        memory[4956] <=  8'h63;        memory[4957] <=  8'h61;        memory[4958] <=  8'h72;        memory[4959] <=  8'h63;        memory[4960] <=  8'h74;        memory[4961] <=  8'h72;        memory[4962] <=  8'h63;        memory[4963] <=  8'h61;        memory[4964] <=  8'h74;        memory[4965] <=  8'h72;        memory[4966] <=  8'h63;        memory[4967] <=  8'h61;        memory[4968] <=  8'h74;        memory[4969] <=  8'h63;        memory[4970] <=  8'h62;        memory[4971] <=  8'h61;        memory[4972] <=  8'h74;        memory[4973] <=  8'h62;        memory[4974] <=  8'h72;        memory[4975] <=  8'h63;        memory[4976] <=  8'h61;        memory[4977] <=  8'h74;        memory[4978] <=  8'h72;        memory[4979] <=  8'h6e;        memory[4980] <=  8'h62;        memory[4981] <=  8'h61;        memory[4982] <=  8'h63;        memory[4983] <=  8'h61;        memory[4984] <=  8'h74;        memory[4985] <=  8'h79;        memory[4986] <=  8'h73;        memory[4987] <=  8'h6e;        memory[4988] <=  8'h63;        memory[4989] <=  8'h74;        memory[4990] <=  8'h61;        memory[4991] <=  8'h6e;        memory[4992] <=  8'h62;        memory[4993] <=  8'h61;        memory[4994] <=  8'h63;        memory[4995] <=  8'h72;        memory[4996] <=  8'h6e;        memory[4997] <=  8'h74;        memory[4998] <=  8'h61;        memory[4999] <=  8'h62;        memory[5000] <=  8'h74;        memory[5001] <=  8'h6e;        memory[5002] <=  8'h61;        memory[5003] <=  8'h72;        memory[5004] <=  8'h62;        memory[5005] <=  8'h78;        memory[5006] <=  8'h74;        memory[5007] <=  8'h61;        memory[5008] <=  8'h72;        memory[5009] <=  8'h62;        memory[5010] <=  8'h61;        memory[5011] <=  8'h72;        memory[5012] <=  8'h74;        memory[5013] <=  8'h74;        memory[5014] <=  8'h62;        memory[5015] <=  8'h61;        memory[5016] <=  8'h72;        memory[5017] <=  8'h74;        memory[5018] <=  8'h78;        memory[5019] <=  8'h61;        memory[5020] <=  8'h74;        memory[5021] <=  8'h6b;        memory[5022] <=  8'h73;        memory[5023] <=  8'h68;        memory[5024] <=  8'h63;        memory[5025] <=  8'h66;        memory[5026] <=  8'h69;        memory[5027] <=  8'h77;        memory[5028] <=  8'h68;        memory[5029] <=  8'h61;        memory[5030] <=  8'h74;        memory[5031] <=  8'h61;        memory[5032] <=  8'h6e;        memory[5033] <=  8'h61;        memory[5034] <=  8'h62;        memory[5035] <=  8'h61;        memory[5036] <=  8'h63;        memory[5037] <=  8'h61;        memory[5038] <=  8'h74;        memory[5039] <=  8'h61;        memory[5040] <=  8'h62;        memory[5041] <=  8'h61;        memory[5042] <=  8'h72;        memory[5043] <=  8'h63;        memory[5044] <=  8'h61;        memory[5045] <=  8'h68;        memory[5046] <=  8'h64;        memory[5047] <=  8'h75;        memory[5048] <=  8'h63;        memory[5049] <=  8'h74;        memory[5050] <=  8'h61;        memory[5051] <=  8'h64;        memory[5052] <=  8'h61;        memory[5053] <=  8'h61;        memory[5054] <=  8'h63;        memory[5055] <=  8'h61;        memory[5056] <=  8'h72;        memory[5057] <=  8'h63;        memory[5058] <=  8'h74;        memory[5059] <=  8'h72;        memory[5060] <=  8'h63;        memory[5061] <=  8'h61;        memory[5062] <=  8'h74;        memory[5063] <=  8'h72;        memory[5064] <=  8'h63;        memory[5065] <=  8'h61;        memory[5066] <=  8'h74;        memory[5067] <=  8'h63;        memory[5068] <=  8'h62;        memory[5069] <=  8'h61;        memory[5070] <=  8'h74;        memory[5071] <=  8'h62;        memory[5072] <=  8'h72;        memory[5073] <=  8'h63;        memory[5074] <=  8'h61;        memory[5075] <=  8'h74;        memory[5076] <=  8'h72;        memory[5077] <=  8'h6e;        memory[5078] <=  8'h62;        memory[5079] <=  8'h61;        memory[5080] <=  8'h63;        memory[5081] <=  8'h61;        memory[5082] <=  8'h74;        memory[5083] <=  8'h79;        memory[5084] <=  8'h73;        memory[5085] <=  8'h6e;        memory[5086] <=  8'h63;        memory[5087] <=  8'h74;        memory[5088] <=  8'h61;        memory[5089] <=  8'h6e;        memory[5090] <=  8'h62;        memory[5091] <=  8'h61;        memory[5092] <=  8'h63;        memory[5093] <=  8'h72;        memory[5094] <=  8'h6e;        memory[5095] <=  8'h74;        memory[5096] <=  8'h61;        memory[5097] <=  8'h62;        memory[5098] <=  8'h74;        memory[5099] <=  8'h6e;        memory[5100] <=  8'h61;        memory[5101] <=  8'h72;        memory[5102] <=  8'h62;        memory[5103] <=  8'h78;        memory[5104] <=  8'h74;        memory[5105] <=  8'h61;        memory[5106] <=  8'h72;        memory[5107] <=  8'h62;        memory[5108] <=  8'h61;        memory[5109] <=  8'h72;        memory[5110] <=  8'h74;        memory[5111] <=  8'h74;        memory[5112] <=  8'h62;        memory[5113] <=  8'h61;        memory[5114] <=  8'h72;        memory[5115] <=  8'h74;        memory[5116] <=  8'h78;        memory[5117] <=  8'h61;        memory[5118] <=  8'h74;        memory[5119] <=  8'h6b;        memory[5120] <=  8'h73;        memory[5121] <=  8'h68;        memory[5122] <=  8'h63;        memory[5123] <=  8'h66;        memory[5124] <=  8'h69;        memory[5125] <=  8'h77;        memory[5126] <=  8'h68;        memory[5127] <=  8'h61;        memory[5128] <=  8'h74;        memory[5129] <=  8'h61;        memory[5130] <=  8'h6e;        memory[5131] <=  8'h61;        memory[5132] <=  8'h62;        memory[5133] <=  8'h61;        memory[5134] <=  8'h63;        memory[5135] <=  8'h61;        memory[5136] <=  8'h74;        memory[5137] <=  8'h61;        memory[5138] <=  8'h62;        memory[5139] <=  8'h61;        memory[5140] <=  8'h72;        memory[5141] <=  8'h63;        memory[5142] <=  8'h61;        memory[5143] <=  8'h68;        memory[5144] <=  8'h64;        memory[5145] <=  8'h75;        memory[5146] <=  8'h63;        memory[5147] <=  8'h74;        memory[5148] <=  8'h61;        memory[5149] <=  8'h64;        memory[5150] <=  8'h61;        memory[5151] <=  8'h61;        memory[5152] <=  8'h63;        memory[5153] <=  8'h61;        memory[5154] <=  8'h72;        memory[5155] <=  8'h63;        memory[5156] <=  8'h74;        memory[5157] <=  8'h72;        memory[5158] <=  8'h63;        memory[5159] <=  8'h61;        memory[5160] <=  8'h74;        memory[5161] <=  8'h72;        memory[5162] <=  8'h63;        memory[5163] <=  8'h61;        memory[5164] <=  8'h74;        memory[5165] <=  8'h63;        memory[5166] <=  8'h62;        memory[5167] <=  8'h61;        memory[5168] <=  8'h74;        memory[5169] <=  8'h62;        memory[5170] <=  8'h72;        memory[5171] <=  8'h63;        memory[5172] <=  8'h61;        memory[5173] <=  8'h74;        memory[5174] <=  8'h72;        memory[5175] <=  8'h6e;        memory[5176] <=  8'h62;        memory[5177] <=  8'h61;        memory[5178] <=  8'h63;        memory[5179] <=  8'h61;        memory[5180] <=  8'h74;        memory[5181] <=  8'h79;        memory[5182] <=  8'h73;        memory[5183] <=  8'h6e;        memory[5184] <=  8'h63;        memory[5185] <=  8'h74;        memory[5186] <=  8'h61;        memory[5187] <=  8'h6e;        memory[5188] <=  8'h62;        memory[5189] <=  8'h61;        memory[5190] <=  8'h63;        memory[5191] <=  8'h72;        memory[5192] <=  8'h6e;        memory[5193] <=  8'h74;        memory[5194] <=  8'h61;        memory[5195] <=  8'h62;        memory[5196] <=  8'h74;        memory[5197] <=  8'h6e;        memory[5198] <=  8'h61;        memory[5199] <=  8'h72;        memory[5200] <=  8'h62;        memory[5201] <=  8'h78;        memory[5202] <=  8'h74;        memory[5203] <=  8'h61;        memory[5204] <=  8'h72;        memory[5205] <=  8'h5d;        memory[5206] <=  8'h5d;        memory[5207] <=  8'h65;        memory[5208] <=  8'h66;        memory[5209] <=  8'h77;        memory[5210] <=  8'h65;        memory[5211] <=  8'h5d;        memory[5212] <=  8'h65;        memory[5213] <=  8'h67;        memory[5214] <=  8'h73;        memory[5215] <=  8'h67;        memory[5216] <=  8'h66;        memory[5217] <=  8'h62;        memory[5218] <=  8'h61;        memory[5219] <=  8'h72;        memory[5220] <=  8'h74;        memory[5221] <=  8'h74;        memory[5222] <=  8'h62;        memory[5223] <=  8'h61;        memory[5224] <=  8'h72;        memory[5225] <=  8'h74;        memory[5226] <=  8'h78;        memory[5227] <=  8'h61;        memory[5228] <=  8'h74;        memory[5229] <=  8'h6b;        memory[5230] <=  8'h73;        memory[5231] <=  8'h68;        memory[5232] <=  8'h63;        memory[5233] <=  8'h66;        memory[5234] <=  8'h69;        memory[5235] <=  8'h77;        memory[5236] <=  8'h68;        memory[5237] <=  8'h61;        memory[5238] <=  8'h74;        memory[5239] <=  8'h61;        memory[5240] <=  8'h6e;        memory[5241] <=  8'h61;        memory[5242] <=  8'h62;        memory[5243] <=  8'h61;        memory[5244] <=  8'h63;        memory[5245] <=  8'h61;        memory[5246] <=  8'h74;        memory[5247] <=  8'h61;        memory[5248] <=  8'h62;        memory[5249] <=  8'h61;        memory[5250] <=  8'h72;        memory[5251] <=  8'h63;        memory[5252] <=  8'h61;        memory[5253] <=  8'h68;        memory[5254] <=  8'h64;        memory[5255] <=  8'h75;        memory[5256] <=  8'h63;        memory[5257] <=  8'h74;        memory[5258] <=  8'h61;        memory[5259] <=  8'h64;        memory[5260] <=  8'h61;        memory[5261] <=  8'h61;        memory[5262] <=  8'h63;        memory[5263] <=  8'h61;        memory[5264] <=  8'h72;        memory[5265] <=  8'h63;        memory[5266] <=  8'h74;        memory[5267] <=  8'h72;        memory[5268] <=  8'h63;        memory[5269] <=  8'h61;        memory[5270] <=  8'h74;        memory[5271] <=  8'h72;        memory[5272] <=  8'h63;        memory[5273] <=  8'h61;        memory[5274] <=  8'h74;        memory[5275] <=  8'h63;        memory[5276] <=  8'h62;        memory[5277] <=  8'h61;        memory[5278] <=  8'h74;        memory[5279] <=  8'h62;        memory[5280] <=  8'h72;        memory[5281] <=  8'h63;        memory[5282] <=  8'h61;        memory[5283] <=  8'h74;        memory[5284] <=  8'h72;        memory[5285] <=  8'h6e;        memory[5286] <=  8'h62;        memory[5287] <=  8'h61;        memory[5288] <=  8'h63;        memory[5289] <=  8'h61;        memory[5290] <=  8'h74;        memory[5291] <=  8'h79;        memory[5292] <=  8'h73;        memory[5293] <=  8'h6e;        memory[5294] <=  8'h63;        memory[5295] <=  8'h74;        memory[5296] <=  8'h61;        memory[5297] <=  8'h6e;        memory[5298] <=  8'h62;        memory[5299] <=  8'h61;        memory[5300] <=  8'h63;        memory[5301] <=  8'h72;        memory[5302] <=  8'h6e;        memory[5303] <=  8'h74;        memory[5304] <=  8'h61;        memory[5305] <=  8'h62;        memory[5306] <=  8'h74;        memory[5307] <=  8'h6e;        memory[5308] <=  8'h61;        memory[5309] <=  8'h72;        memory[5310] <=  8'h62;        memory[5311] <=  8'h78;        memory[5312] <=  8'h74;        memory[5313] <=  8'h61;        memory[5314] <=  8'h72;        memory[5315] <=  8'h62;        memory[5316] <=  8'h61;        memory[5317] <=  8'h72;        memory[5318] <=  8'h74;        memory[5319] <=  8'h74;        memory[5320] <=  8'h62;        memory[5321] <=  8'h61;        memory[5322] <=  8'h72;        memory[5323] <=  8'h74;        memory[5324] <=  8'h78;        memory[5325] <=  8'h61;        memory[5326] <=  8'h74;        memory[5327] <=  8'h6b;        memory[5328] <=  8'h73;        memory[5329] <=  8'h68;        memory[5330] <=  8'h63;        memory[5331] <=  8'h66;        memory[5332] <=  8'h69;        memory[5333] <=  8'h77;        memory[5334] <=  8'h68;        memory[5335] <=  8'h61;        memory[5336] <=  8'h74;        memory[5337] <=  8'h61;        memory[5338] <=  8'h6e;        memory[5339] <=  8'h61;        memory[5340] <=  8'h62;        memory[5341] <=  8'h61;        memory[5342] <=  8'h63;        memory[5343] <=  8'h61;        memory[5344] <=  8'h74;        memory[5345] <=  8'h61;        memory[5346] <=  8'h62;        memory[5347] <=  8'h61;        memory[5348] <=  8'h72;        memory[5349] <=  8'h63;        memory[5350] <=  8'h61;        memory[5351] <=  8'h68;        memory[5352] <=  8'h64;        memory[5353] <=  8'h75;        memory[5354] <=  8'h63;        memory[5355] <=  8'h74;        memory[5356] <=  8'h61;        memory[5357] <=  8'h64;        memory[5358] <=  8'h61;        memory[5359] <=  8'h61;        memory[5360] <=  8'h63;        memory[5361] <=  8'h61;        memory[5362] <=  8'h72;        memory[5363] <=  8'h63;        memory[5364] <=  8'h74;        memory[5365] <=  8'h72;        memory[5366] <=  8'h63;        memory[5367] <=  8'h61;        memory[5368] <=  8'h74;        memory[5369] <=  8'h72;        memory[5370] <=  8'h63;        memory[5371] <=  8'h61;        memory[5372] <=  8'h74;        memory[5373] <=  8'h63;        memory[5374] <=  8'h62;        memory[5375] <=  8'h61;        memory[5376] <=  8'h74;        memory[5377] <=  8'h62;        memory[5378] <=  8'h72;        memory[5379] <=  8'h63;        memory[5380] <=  8'h61;        memory[5381] <=  8'h74;        memory[5382] <=  8'h72;        memory[5383] <=  8'h6e;        memory[5384] <=  8'h62;        memory[5385] <=  8'h61;        memory[5386] <=  8'h63;        memory[5387] <=  8'h61;        memory[5388] <=  8'h74;        memory[5389] <=  8'h79;        memory[5390] <=  8'h73;        memory[5391] <=  8'h6e;        memory[5392] <=  8'h63;        memory[5393] <=  8'h74;        memory[5394] <=  8'h61;        memory[5395] <=  8'h6e;        memory[5396] <=  8'h62;        memory[5397] <=  8'h61;        memory[5398] <=  8'h63;        memory[5399] <=  8'h72;        memory[5400] <=  8'h6e;        memory[5401] <=  8'h74;        memory[5402] <=  8'h61;        memory[5403] <=  8'h62;        memory[5404] <=  8'h74;        memory[5405] <=  8'h6e;        memory[5406] <=  8'h61;        memory[5407] <=  8'h72;        memory[5408] <=  8'h62;        memory[5409] <=  8'h78;        memory[5410] <=  8'h74;        memory[5411] <=  8'h61;        memory[5412] <=  8'h72;        memory[5413] <=  8'h64;        memory[5414] <=  8'h66;        memory[5415] <=  8'h73;        memory[5416] <=  8'h67;        memory[5417] <=  8'h76;        memory[5418] <=  8'h68;        memory[5419] <=  8'h62;        memory[5420] <=  8'h6b;        memory[5421] <=  8'h6a;        memory[5422] <=  8'h6e;        memory[5423] <=  8'h6d;        memory[5424] <=  8'h62;        memory[5425] <=  8'h76;        memory[5426] <=  8'h78;        memory[5427] <=  8'h63;        memory[5428] <=  8'h73;        memory[5429] <=  8'h66;        memory[5430] <=  8'h72;        memory[5431] <=  8'h74;        memory[5432] <=  8'h79;        memory[5433] <=  8'h75;        memory[5434] <=  8'h6a;        memory[5435] <=  8'h6e;        memory[5436] <=  8'h62;        memory[5437] <=  8'h76;        memory[5438] <=  8'h63;        memory[5439] <=  8'h64;        memory[5440] <=  8'h74;        memory[5441] <=  8'h79;        memory[5442] <=  8'h75;        memory[5443] <=  8'h69;        memory[5444] <=  8'h6b;        memory[5445] <=  8'h6d;        memory[5446] <=  8'h6e;        memory[5447] <=  8'h62;        memory[5448] <=  8'h76;        memory[5449] <=  8'h63;        memory[5450] <=  8'h78;        memory[5451] <=  8'h73;        memory[5452] <=  8'h64;        memory[5453] <=  8'h72;        memory[5454] <=  8'h74;        memory[5455] <=  8'h79;        memory[5456] <=  8'h75;        memory[5457] <=  8'h69;        memory[5458] <=  8'h6b;        memory[5459] <=  8'h6d;        memory[5460] <=  8'h6e;        memory[5461] <=  8'h62;        memory[5462] <=  8'h76;        memory[5463] <=  8'h63;        memory[5464] <=  8'h73;        memory[5465] <=  8'h77;        memory[5466] <=  8'h33;        memory[5467] <=  8'h34;        memory[5468] <=  8'h35;        memory[5469] <=  8'h36;        memory[5470] <=  8'h37;        memory[5471] <=  8'h38;        memory[5472] <=  8'h69;        memory[5473] <=  8'h6b;        memory[5474] <=  8'h6d;        memory[5475] <=  8'h6e;        memory[5476] <=  8'h62;        memory[5477] <=  8'h76;        memory[5478] <=  8'h63;        memory[5479] <=  8'h64;        memory[5480] <=  8'h65;        memory[5481] <=  8'h72;        memory[5482] <=  8'h36;        memory[5483] <=  8'h37;        memory[5484] <=  8'h38;        memory[5485] <=  8'h69;        memory[5486] <=  8'h6f;        memory[5487] <=  8'h6b;        memory[5488] <=  8'h6a;        memory[5489] <=  8'h6e;        memory[5490] <=  8'h62;        memory[5491] <=  8'h76;        memory[5492] <=  8'h63;        memory[5493] <=  8'h64;        memory[5494] <=  8'h72;        memory[5495] <=  8'h74;        memory[5496] <=  8'h79;        memory[5497] <=  8'h75;        memory[5498] <=  8'h73;        memory[5499] <=  8'h6a;        memory[5500] <=  8'h63;        memory[5501] <=  8'h6e;        memory[5502] <=  8'h62;        memory[5503] <=  8'h64;        memory[5504] <=  8'h66;        memory[5505] <=  8'h73;        memory[5506] <=  8'h74;        memory[5507] <=  8'h79;        memory[5508] <=  8'h75;        memory[5509] <=  8'h61;        memory[5510] <=  8'h69;        memory[5511] <=  8'h6b;        memory[5512] <=  8'h78;        memory[5513] <=  8'h6d;        memory[5514] <=  8'h6e;        memory[5515] <=  8'h73;        memory[5516] <=  8'h6a;        memory[5517] <=  8'h6f;        memory[5518] <=  8'h64;        memory[5519] <=  8'h6c;        memory[5520] <=  8'h63;        memory[5521] <=  8'h78;        memory[5522] <=  8'h62;        memory[5523] <=  8'h61;        memory[5524] <=  8'h72;        memory[5525] <=  8'h74;        memory[5526] <=  8'h78;        memory[5527] <=  8'h61;        memory[5528] <=  8'h74;        memory[5529] <=  8'h6b;        memory[5530] <=  8'h73;        memory[5531] <=  8'h68;        memory[5532] <=  8'h63;        memory[5533] <=  8'h66;        memory[5534] <=  8'h69;        memory[5535] <=  8'h77;        memory[5536] <=  8'h68;        memory[5537] <=  8'h61;        memory[5538] <=  8'h74;        memory[5539] <=  8'h61;        memory[5540] <=  8'h6e;        memory[5541] <=  8'h61;        memory[5542] <=  8'h62;        memory[5543] <=  8'h61;        memory[5544] <=  8'h63;        memory[5545] <=  8'h61;        memory[5546] <=  8'h74;        memory[5547] <=  8'h61;        memory[5548] <=  8'h62;        memory[5549] <=  8'h61;        memory[5550] <=  8'h72;        memory[5551] <=  8'h63;        memory[5552] <=  8'h61;        memory[5553] <=  8'h68;        memory[5554] <=  8'h64;        memory[5555] <=  8'h75;        memory[5556] <=  8'h63;        memory[5557] <=  8'h74;        memory[5558] <=  8'h61;        memory[5559] <=  8'h64;        memory[5560] <=  8'h61;        memory[5561] <=  8'h61;        memory[5562] <=  8'h63;        memory[5563] <=  8'h61;        memory[5564] <=  8'h72;        memory[5565] <=  8'h62;        memory[5566] <=  8'h61;        memory[5567] <=  8'h72;        memory[5568] <=  8'h74;        memory[5569] <=  8'h78;        memory[5570] <=  8'h61;        memory[5571] <=  8'h74;        memory[5572] <=  8'h6b;        memory[5573] <=  8'h73;        memory[5574] <=  8'h68;        memory[5575] <=  8'h63;        memory[5576] <=  8'h66;        memory[5577] <=  8'h69;        memory[5578] <=  8'h77;        memory[5579] <=  8'h68;        memory[5580] <=  8'h61;        memory[5581] <=  8'h74;        memory[5582] <=  8'h61;        memory[5583] <=  8'h6e;        memory[5584] <=  8'h61;        memory[5585] <=  8'h62;        memory[5586] <=  8'h61;        memory[5587] <=  8'h63;        memory[5588] <=  8'h61;        memory[5589] <=  8'h74;        memory[5590] <=  8'h61;        memory[5591] <=  8'h62;        memory[5592] <=  8'h61;        memory[5593] <=  8'h72;        memory[5594] <=  8'h63;        memory[5595] <=  8'h61;        memory[5596] <=  8'h68;        memory[5597] <=  8'h64;        memory[5598] <=  8'h75;        memory[5599] <=  8'h63;        memory[5600] <=  8'h74;        memory[5601] <=  8'h61;        memory[5602] <=  8'h64;        memory[5603] <=  8'h61;        memory[5604] <=  8'h61;        memory[5605] <=  8'h63;        memory[5606] <=  8'h61;        memory[5607] <=  8'h72;        memory[5608] <=  8'h62;        memory[5609] <=  8'h61;        memory[5610] <=  8'h72;        memory[5611] <=  8'h74;        memory[5612] <=  8'h78;        memory[5613] <=  8'h61;        memory[5614] <=  8'h74;        memory[5615] <=  8'h6b;        memory[5616] <=  8'h73;        memory[5617] <=  8'h68;        memory[5618] <=  8'h63;        memory[5619] <=  8'h66;        memory[5620] <=  8'h69;        memory[5621] <=  8'h77;        memory[5622] <=  8'h68;        memory[5623] <=  8'h61;        memory[5624] <=  8'h74;        memory[5625] <=  8'h61;        memory[5626] <=  8'h6e;        memory[5627] <=  8'h61;        memory[5628] <=  8'h62;        memory[5629] <=  8'h61;        memory[5630] <=  8'h63;        memory[5631] <=  8'h61;        memory[5632] <=  8'h74;        memory[5633] <=  8'h61;        memory[5634] <=  8'h62;        memory[5635] <=  8'h61;        memory[5636] <=  8'h72;        memory[5637] <=  8'h63;        memory[5638] <=  8'h61;        memory[5639] <=  8'h68;        memory[5640] <=  8'h64;        memory[5641] <=  8'h75;        memory[5642] <=  8'h63;        memory[5643] <=  8'h74;        memory[5644] <=  8'h61;        memory[5645] <=  8'h64;        memory[5646] <=  8'h61;        memory[5647] <=  8'h61;        memory[5648] <=  8'h63;        memory[5649] <=  8'h61;        memory[5650] <=  8'h72;        memory[5651] <=  8'h62;        memory[5652] <=  8'h61;        memory[5653] <=  8'h72;        memory[5654] <=  8'h74;        memory[5655] <=  8'h78;        memory[5656] <=  8'h61;        memory[5657] <=  8'h74;        memory[5658] <=  8'h6b;        memory[5659] <=  8'h73;        memory[5660] <=  8'h68;        memory[5661] <=  8'h63;        memory[5662] <=  8'h66;        memory[5663] <=  8'h69;        memory[5664] <=  8'h77;        memory[5665] <=  8'h68;        memory[5666] <=  8'h61;        memory[5667] <=  8'h74;        memory[5668] <=  8'h61;        memory[5669] <=  8'h6e;        memory[5670] <=  8'h61;        memory[5671] <=  8'h62;        memory[5672] <=  8'h61;        memory[5673] <=  8'h63;        memory[5674] <=  8'h61;        memory[5675] <=  8'h74;        memory[5676] <=  8'h61;        memory[5677] <=  8'h62;        memory[5678] <=  8'h61;        memory[5679] <=  8'h72;        memory[5680] <=  8'h63;        memory[5681] <=  8'h61;        memory[5682] <=  8'h68;        memory[5683] <=  8'h64;        memory[5684] <=  8'h75;        memory[5685] <=  8'h63;        memory[5686] <=  8'h74;        memory[5687] <=  8'h61;        memory[5688] <=  8'h64;        memory[5689] <=  8'h61;        memory[5690] <=  8'h61;        memory[5691] <=  8'h63;        memory[5692] <=  8'h61;        memory[5693] <=  8'h72;        memory[5694] <=  8'h62;        memory[5695] <=  8'h61;        memory[5696] <=  8'h72;        memory[5697] <=  8'h74;        memory[5698] <=  8'h78;        memory[5699] <=  8'h61;        memory[5700] <=  8'h74;        memory[5701] <=  8'h6b;        memory[5702] <=  8'h73;        memory[5703] <=  8'h68;        memory[5704] <=  8'h63;        memory[5705] <=  8'h66;        memory[5706] <=  8'h69;        memory[5707] <=  8'h77;        memory[5708] <=  8'h68;        memory[5709] <=  8'h61;        memory[5710] <=  8'h74;        memory[5711] <=  8'h61;        memory[5712] <=  8'h6e;        memory[5713] <=  8'h61;        memory[5714] <=  8'h62;        memory[5715] <=  8'h61;        memory[5716] <=  8'h63;        memory[5717] <=  8'h61;        memory[5718] <=  8'h74;        memory[5719] <=  8'h61;        memory[5720] <=  8'h62;        memory[5721] <=  8'h61;        memory[5722] <=  8'h72;        memory[5723] <=  8'h63;        memory[5724] <=  8'h61;        memory[5725] <=  8'h68;        memory[5726] <=  8'h64;        memory[5727] <=  8'h75;        memory[5728] <=  8'h63;        memory[5729] <=  8'h74;        memory[5730] <=  8'h61;        memory[5731] <=  8'h64;        memory[5732] <=  8'h61;        memory[5733] <=  8'h61;        memory[5734] <=  8'h63;        memory[5735] <=  8'h61;        memory[5736] <=  8'h72;        memory[5737] <=  8'h62;        memory[5738] <=  8'h61;        memory[5739] <=  8'h72;        memory[5740] <=  8'h74;        memory[5741] <=  8'h78;        memory[5742] <=  8'h61;        memory[5743] <=  8'h74;        memory[5744] <=  8'h6b;        memory[5745] <=  8'h73;        memory[5746] <=  8'h68;        memory[5747] <=  8'h63;        memory[5748] <=  8'h66;        memory[5749] <=  8'h69;        memory[5750] <=  8'h77;        memory[5751] <=  8'h68;        memory[5752] <=  8'h61;        memory[5753] <=  8'h74;        memory[5754] <=  8'h61;        memory[5755] <=  8'h6e;        memory[5756] <=  8'h61;        memory[5757] <=  8'h62;        memory[5758] <=  8'h61;        memory[5759] <=  8'h63;        memory[5760] <=  8'h61;        memory[5761] <=  8'h74;        memory[5762] <=  8'h61;        memory[5763] <=  8'h62;        memory[5764] <=  8'h61;        memory[5765] <=  8'h72;        memory[5766] <=  8'h63;        memory[5767] <=  8'h61;        memory[5768] <=  8'h68;        memory[5769] <=  8'h64;        memory[5770] <=  8'h75;        memory[5771] <=  8'h63;        memory[5772] <=  8'h74;        memory[5773] <=  8'h61;        memory[5774] <=  8'h64;        memory[5775] <=  8'h61;        memory[5776] <=  8'h61;        memory[5777] <=  8'h63;        memory[5778] <=  8'h61;        memory[5779] <=  8'h72;        memory[5780] <=  8'h62;        memory[5781] <=  8'h61;        memory[5782] <=  8'h72;        memory[5783] <=  8'h74;        memory[5784] <=  8'h78;        memory[5785] <=  8'h61;        memory[5786] <=  8'h74;        memory[5787] <=  8'h6b;        memory[5788] <=  8'h73;        memory[5789] <=  8'h68;        memory[5790] <=  8'h63;        memory[5791] <=  8'h66;        memory[5792] <=  8'h69;        memory[5793] <=  8'h77;        memory[5794] <=  8'h68;        memory[5795] <=  8'h61;        memory[5796] <=  8'h74;        memory[5797] <=  8'h61;        memory[5798] <=  8'h6e;        memory[5799] <=  8'h61;        memory[5800] <=  8'h62;        memory[5801] <=  8'h61;        memory[5802] <=  8'h63;        memory[5803] <=  8'h61;        memory[5804] <=  8'h74;        memory[5805] <=  8'h61;        memory[5806] <=  8'h62;        memory[5807] <=  8'h61;        memory[5808] <=  8'h72;        memory[5809] <=  8'h63;        memory[5810] <=  8'h61;        memory[5811] <=  8'h68;        memory[5812] <=  8'h64;        memory[5813] <=  8'h75;        memory[5814] <=  8'h63;        memory[5815] <=  8'h74;        memory[5816] <=  8'h61;        memory[5817] <=  8'h64;        memory[5818] <=  8'h61;        memory[5819] <=  8'h61;        memory[5820] <=  8'h63;        memory[5821] <=  8'h61;        memory[5822] <=  8'h72;        memory[5823] <=  8'h62;        memory[5824] <=  8'h61;        memory[5825] <=  8'h72;        memory[5826] <=  8'h74;        memory[5827] <=  8'h78;        memory[5828] <=  8'h61;        memory[5829] <=  8'h74;        memory[5830] <=  8'h6b;        memory[5831] <=  8'h73;        memory[5832] <=  8'h68;        memory[5833] <=  8'h63;        memory[5834] <=  8'h66;        memory[5835] <=  8'h69;        memory[5836] <=  8'h77;        memory[5837] <=  8'h68;        memory[5838] <=  8'h61;        memory[5839] <=  8'h74;        memory[5840] <=  8'h61;        memory[5841] <=  8'h6e;        memory[5842] <=  8'h61;        memory[5843] <=  8'h62;        memory[5844] <=  8'h61;        memory[5845] <=  8'h63;        memory[5846] <=  8'h61;        memory[5847] <=  8'h74;        memory[5848] <=  8'h61;        memory[5849] <=  8'h62;        memory[5850] <=  8'h61;        memory[5851] <=  8'h72;        memory[5852] <=  8'h63;        memory[5853] <=  8'h61;        memory[5854] <=  8'h68;        memory[5855] <=  8'h64;        memory[5856] <=  8'h75;        memory[5857] <=  8'h63;        memory[5858] <=  8'h74;        memory[5859] <=  8'h61;        memory[5860] <=  8'h64;        memory[5861] <=  8'h61;        memory[5862] <=  8'h61;        memory[5863] <=  8'h63;        memory[5864] <=  8'h61;        memory[5865] <=  8'h72;        memory[5866] <=  8'h62;        memory[5867] <=  8'h61;        memory[5868] <=  8'h72;        memory[5869] <=  8'h74;        memory[5870] <=  8'h78;        memory[5871] <=  8'h61;        memory[5872] <=  8'h74;        memory[5873] <=  8'h6b;        memory[5874] <=  8'h73;        memory[5875] <=  8'h68;        memory[5876] <=  8'h63;        memory[5877] <=  8'h66;        memory[5878] <=  8'h69;        memory[5879] <=  8'h77;        memory[5880] <=  8'h68;        memory[5881] <=  8'h61;        memory[5882] <=  8'h74;        memory[5883] <=  8'h61;        memory[5884] <=  8'h6e;        memory[5885] <=  8'h61;        memory[5886] <=  8'h62;        memory[5887] <=  8'h61;        memory[5888] <=  8'h63;        memory[5889] <=  8'h61;        memory[5890] <=  8'h74;        memory[5891] <=  8'h61;        memory[5892] <=  8'h62;        memory[5893] <=  8'h61;        memory[5894] <=  8'h72;        memory[5895] <=  8'h63;        memory[5896] <=  8'h61;        memory[5897] <=  8'h68;        memory[5898] <=  8'h64;        memory[5899] <=  8'h75;        memory[5900] <=  8'h63;        memory[5901] <=  8'h74;        memory[5902] <=  8'h61;        memory[5903] <=  8'h64;        memory[5904] <=  8'h61;        memory[5905] <=  8'h61;        memory[5906] <=  8'h63;        memory[5907] <=  8'h61;        memory[5908] <=  8'h72;        memory[5909] <=  8'h62;        memory[5910] <=  8'h61;        memory[5911] <=  8'h72;        memory[5912] <=  8'h74;        memory[5913] <=  8'h74;        memory[5914] <=  8'h62;        memory[5915] <=  8'h61;        memory[5916] <=  8'h72;        memory[5917] <=  8'h74;        memory[5918] <=  8'h78;        memory[5919] <=  8'h61;        memory[5920] <=  8'h74;        memory[5921] <=  8'h6b;        memory[5922] <=  8'h73;        memory[5923] <=  8'h68;        memory[5924] <=  8'h63;        memory[5925] <=  8'h66;        memory[5926] <=  8'h69;        memory[5927] <=  8'h77;        memory[5928] <=  8'h68;        memory[5929] <=  8'h61;        memory[5930] <=  8'h74;        memory[5931] <=  8'h61;        memory[5932] <=  8'h6e;        memory[5933] <=  8'h61;        memory[5934] <=  8'h62;        memory[5935] <=  8'h61;        memory[5936] <=  8'h63;        memory[5937] <=  8'h61;        memory[5938] <=  8'h74;        memory[5939] <=  8'h61;        memory[5940] <=  8'h62;        memory[5941] <=  8'h61;        memory[5942] <=  8'h72;        memory[5943] <=  8'h63;        memory[5944] <=  8'h61;        memory[5945] <=  8'h68;        memory[5946] <=  8'h64;        memory[5947] <=  8'h75;        memory[5948] <=  8'h63;        memory[5949] <=  8'h74;        memory[5950] <=  8'h61;        memory[5951] <=  8'h64;        memory[5952] <=  8'h61;        memory[5953] <=  8'h61;        memory[5954] <=  8'h63;        memory[5955] <=  8'h61;        memory[5956] <=  8'h72;        memory[5957] <=  8'h63;        memory[5958] <=  8'h74;        memory[5959] <=  8'h72;        memory[5960] <=  8'h63;        memory[5961] <=  8'h61;        memory[5962] <=  8'h74;        memory[5963] <=  8'h72;        memory[5964] <=  8'h63;        memory[5965] <=  8'h61;        memory[5966] <=  8'h74;        memory[5967] <=  8'h63;        memory[5968] <=  8'h62;        memory[5969] <=  8'h61;        memory[5970] <=  8'h74;        memory[5971] <=  8'h62;        memory[5972] <=  8'h72;        memory[5973] <=  8'h63;        memory[5974] <=  8'h61;        memory[5975] <=  8'h72;        memory[5976] <=  8'h62;        memory[5977] <=  8'h78;        memory[5978] <=  8'h74;        memory[5979] <=  8'h61;        memory[5980] <=  8'h72;        memory[5981] <=  8'h64;        memory[5982] <=  8'h66;        memory[5983] <=  8'h73;        memory[5984] <=  8'h67;        memory[5985] <=  8'h76;        memory[5986] <=  8'h68;        memory[5987] <=  8'h62;        memory[5988] <=  8'h6b;        memory[5989] <=  8'h6a;        memory[5990] <=  8'h6e;        memory[5991] <=  8'h6d;        memory[5992] <=  8'h62;        memory[5993] <=  8'h76;        memory[5994] <=  8'h78;        memory[5995] <=  8'h63;        memory[5996] <=  8'h73;        memory[5997] <=  8'h66;        memory[5998] <=  8'h72;        memory[5999] <=  8'h74;        memory[6000] <=  8'h79;        memory[6001] <=  8'h75;        memory[6002] <=  8'h6a;        memory[6003] <=  8'h6e;        memory[6004] <=  8'h62;        memory[6005] <=  8'h76;        memory[6006] <=  8'h63;        memory[6007] <=  8'h64;        memory[6008] <=  8'h74;        memory[6009] <=  8'h79;        memory[6010] <=  8'h75;        memory[6011] <=  8'h69;        memory[6012] <=  8'h6b;        memory[6013] <=  8'h6d;        memory[6014] <=  8'h6e;        memory[6015] <=  8'h62;        memory[6016] <=  8'h76;        memory[6017] <=  8'h63;        memory[6018] <=  8'h78;        memory[6019] <=  8'h73;        memory[6020] <=  8'h64;        memory[6021] <=  8'h72;        memory[6022] <=  8'h74;        memory[6023] <=  8'h79;        memory[6024] <=  8'h75;        memory[6025] <=  8'h69;        memory[6026] <=  8'h6b;        memory[6027] <=  8'h6d;        memory[6028] <=  8'h6e;        memory[6029] <=  8'h62;        memory[6030] <=  8'h76;        memory[6031] <=  8'h63;        memory[6032] <=  8'h73;        memory[6033] <=  8'h77;        memory[6034] <=  8'h33;        memory[6035] <=  8'h34;        memory[6036] <=  8'h35;        memory[6037] <=  8'h36;        memory[6038] <=  8'h37;        memory[6039] <=  8'h38;        memory[6040] <=  8'h69;        memory[6041] <=  8'h6b;        memory[6042] <=  8'h6d;        memory[6043] <=  8'h6e;        memory[6044] <=  8'h62;        memory[6045] <=  8'h76;        memory[6046] <=  8'h63;        memory[6047] <=  8'h64;        memory[6048] <=  8'h65;        memory[6049] <=  8'h72;        memory[6050] <=  8'h36;        memory[6051] <=  8'h37;        memory[6052] <=  8'h38;        memory[6053] <=  8'h69;        memory[6054] <=  8'h6f;        memory[6055] <=  8'h6b;        memory[6056] <=  8'h6a;        memory[6057] <=  8'h6e;        memory[6058] <=  8'h62;        memory[6059] <=  8'h76;        memory[6060] <=  8'h63;        memory[6061] <=  8'h64;        memory[6062] <=  8'h72;        memory[6063] <=  8'h74;        memory[6064] <=  8'h79;        memory[6065] <=  8'h75;        memory[6066] <=  8'h73;        memory[6067] <=  8'h6a;        memory[6068] <=  8'h63;        memory[6069] <=  8'h6e;        memory[6070] <=  8'h62;        memory[6071] <=  8'h64;        memory[6072] <=  8'h66;        memory[6073] <=  8'h73;        memory[6074] <=  8'h74;        memory[6075] <=  8'h79;        memory[6076] <=  8'h75;        memory[6077] <=  8'h61;        memory[6078] <=  8'h69;        memory[6079] <=  8'h6b;        memory[6080] <=  8'h78;        memory[6081] <=  8'h6d;        memory[6082] <=  8'h6e;        memory[6083] <=  8'h73;        memory[6084] <=  8'h6a;        memory[6085] <=  8'h6f;        memory[6086] <=  8'h64;        memory[6087] <=  8'h6c;        memory[6088] <=  8'h63;        memory[6089] <=  8'h78;        memory[6090] <=  8'h2c;        memory[6091] <=  8'h6d;        memory[6092] <=  8'h73;        memory[6093] <=  8'h6b;        memory[6094] <=  8'h64;        memory[6095] <=  8'h6c;        memory[6096] <=  8'h70;        memory[6097] <=  8'h5b;        memory[6098] <=  8'h3b;        memory[6099] <=  8'h73;        memory[6100] <=  8'h6c;        memory[6101] <=  8'h64;        memory[6102] <=  8'h70;        memory[6103] <=  8'h76;        memory[6104] <=  8'h63;        memory[6105] <=  8'h5b;        memory[6106] <=  8'h78;        memory[6107] <=  8'h76;        memory[6108] <=  8'h63;        memory[6109] <=  8'h5b;        memory[6110] <=  8'h78;        memory[6111] <=  8'h70;        memory[6112] <=  8'h6f;        memory[6113] <=  8'h20;        memory[6114] <=  8'h62;        memory[6115] <=  8'h61;        memory[6116] <=  8'h72;        memory[6117] <=  8'h74;        memory[6118] <=  8'h74;        memory[6119] <=  8'h62;        memory[6120] <=  8'h61;        memory[6121] <=  8'h72;        memory[6122] <=  8'h74;        memory[6123] <=  8'h78;        memory[6124] <=  8'h61;        memory[6125] <=  8'h74;        memory[6126] <=  8'h6b;        memory[6127] <=  8'h73;        memory[6128] <=  8'h68;        memory[6129] <=  8'h63;        memory[6130] <=  8'h66;        memory[6131] <=  8'h69;        memory[6132] <=  8'h77;        memory[6133] <=  8'h68;        memory[6134] <=  8'h61;        memory[6135] <=  8'h69;        memory[6136] <=  8'h6a;        memory[6137] <=  8'h78;        memory[6138] <=  8'h5d;        memory[6139] <=  8'h65;        memory[6140] <=  8'h6b;        memory[6141] <=  8'h6f;        memory[6142] <=  8'h39;        memory[6143] <=  8'h64;        memory[6144] <=  8'h75;        memory[6145] <=  8'h38;        memory[6146] <=  8'h79;        memory[6147] <=  8'h20;        memory[6148] <=  8'h37;        memory[6149] <=  8'h63;        memory[6150] <=  8'h67;        memory[6151] <=  8'h78;        memory[6152] <=  8'h63;        memory[6153] <=  8'h75;        memory[6154] <=  8'h68;        memory[6155] <=  8'h69;        memory[6156] <=  8'h6a;        memory[6157] <=  8'h77;        memory[6158] <=  8'h69;        memory[6159] <=  8'h64;        memory[6160] <=  8'h66;        memory[6161] <=  8'h68;        memory[6162] <=  8'h75;        memory[6163] <=  8'h76;        memory[6164] <=  8'h64;        memory[6165] <=  8'h62;        memory[6166] <=  8'h66;        memory[6167] <=  8'h6a;        memory[6168] <=  8'h6e;        memory[6169] <=  8'h6b;        memory[6170] <=  8'h6a;        memory[6171] <=  8'h65;        memory[6172] <=  8'h38;        memory[6173] <=  8'h66;        memory[6174] <=  8'h37;        memory[6175] <=  8'h67;        memory[6176] <=  8'h79;        memory[6177] <=  8'h76;        memory[6178] <=  8'h63;        memory[6179] <=  8'h68;        memory[6180] <=  8'h69;        memory[6181] <=  8'h6a;        memory[6182] <=  8'h33;        memory[6183] <=  8'h65;        memory[6184] <=  8'h67;        memory[6185] <=  8'h79;        memory[6186] <=  8'h72;        memory[6187] <=  8'h64;        memory[6188] <=  8'h62;        memory[6189] <=  8'h6e;        memory[6190] <=  8'h63;        memory[6191] <=  8'h7a;        memory[6192] <=  8'h6a;        memory[6193] <=  8'h6f;        memory[6194] <=  8'h66;        memory[6195] <=  8'h78;        memory[6196] <=  8'h6a;        memory[6197] <=  8'h69;        memory[6198] <=  8'h63;        memory[6199] <=  8'h68;        memory[6200] <=  8'h62;        memory[6201] <=  8'h6e;        memory[6202] <=  8'h6d;        memory[6203] <=  8'h63;        memory[6204] <=  8'h73;        memory[6205] <=  8'h6c;        memory[6206] <=  8'h6b;        memory[6207] <=  8'h6a;        memory[6208] <=  8'h69;        memory[6209] <=  8'h68;        memory[6210] <=  8'h76;        memory[6211] <=  8'h75;        memory[6212] <=  8'h69;        memory[6213] <=  8'h64;        memory[6214] <=  8'h68;        memory[6215] <=  8'h75;        memory[6216] <=  8'h67;        memory[6217] <=  8'h79;        memory[6218] <=  8'h62;        memory[6219] <=  8'h68;        memory[6220] <=  8'h65;        memory[6221] <=  8'h6a;        memory[6222] <=  8'h72;        memory[6223] <=  8'h6b;        memory[6224] <=  8'h6a;        memory[6225] <=  8'h6f;        memory[6226] <=  8'h64;        memory[6227] <=  8'h67;        memory[6228] <=  8'h69;        memory[6229] <=  8'h75;        memory[6230] <=  8'h69;        memory[6231] <=  8'h67;        memory[6232] <=  8'h76;        memory[6233] <=  8'h79;        memory[6234] <=  8'h75;        memory[6235] <=  8'h67;        memory[6236] <=  8'h78;        memory[6237] <=  8'h68;        memory[6238] <=  8'h63;        memory[6239] <=  8'h20;        memory[6240] <=  8'h20;        memory[6241] <=  8'h20;        memory[6242] <=  8'h78;        memory[6243] <=  8'h76;        memory[6244] <=  8'h20;        memory[6245] <=  8'h63;        memory[6246] <=  8'h78;        memory[6247] <=  8'h67;        memory[6248] <=  8'h79;        memory[6249] <=  8'h63;        memory[6250] <=  8'h75;        memory[6251] <=  8'h68;        memory[6252] <=  8'h6a;        memory[6253] <=  8'h6b;        memory[6254] <=  8'h61;        memory[6255] <=  8'h6c;        memory[6256] <=  8'h78;        memory[6257] <=  8'h76;        memory[6258] <=  8'h70;        memory[6259] <=  8'h6f;        memory[6260] <=  8'h69;        memory[6261] <=  8'h6a;        memory[6262] <=  8'h69;        memory[6263] <=  8'h68;        memory[6264] <=  8'h6a;        memory[6265] <=  8'h62;        memory[6266] <=  8'h77;        memory[6267] <=  8'h65;        memory[6268] <=  8'h6e;        memory[6269] <=  8'h61;        memory[6270] <=  8'h66;        memory[6271] <=  8'h6d;        memory[6272] <=  8'h64;        memory[6273] <=  8'h6b;        memory[6274] <=  8'h6d;        memory[6275] <=  8'h76;        memory[6276] <=  8'h6c;        memory[6277] <=  8'h63;        memory[6278] <=  8'h6f;        memory[6279] <=  8'h64;        memory[6280] <=  8'h69;        memory[6281] <=  8'h75;        memory[6282] <=  8'h68;        memory[6283] <=  8'h73;        memory[6284] <=  8'h66;        memory[6285] <=  8'h65;        memory[6286] <=  8'h62;        memory[6287] <=  8'h6e;        memory[6288] <=  8'h64;        memory[6289] <=  8'h73;        memory[6290] <=  8'h63;        memory[6291] <=  8'h6b;        memory[6292] <=  8'h20;        memory[6293] <=  8'h78;        memory[6294] <=  8'h6a;        memory[6295] <=  8'h78;        memory[6296] <=  8'h63;        memory[6297] <=  8'h73;        memory[6298] <=  8'h64;        memory[6299] <=  8'h66;        memory[6300] <=  8'h6b;        memory[6301] <=  8'h64;        memory[6302] <=  8'h6e;        memory[6303] <=  8'h6d;        memory[6304] <=  8'h64;        memory[6305] <=  8'h73;        memory[6306] <=  8'h63;        memory[6307] <=  8'h6b;        memory[6308] <=  8'h78;        memory[6309] <=  8'h6c;        memory[6310] <=  8'h6f;        memory[6311] <=  8'h66;        memory[6312] <=  8'h6a;        memory[6313] <=  8'h69;        memory[6314] <=  8'h61;        memory[6315] <=  8'h62;        memory[6316] <=  8'h6e;        memory[6317] <=  8'h20;        memory[6318] <=  8'h78;        memory[6319] <=  8'h6b;        memory[6320] <=  8'h6d;        memory[6321] <=  8'h20;        memory[6322] <=  8'h6f;        memory[6323] <=  8'h63;        memory[6324] <=  8'h76;        memory[6325] <=  8'h73;        memory[6326] <=  8'h64;        memory[6327] <=  8'h69;        memory[6328] <=  8'h66;        memory[6329] <=  8'h68;        memory[6330] <=  8'h65;        memory[6331] <=  8'h71;        memory[6332] <=  8'h6a;        memory[6333] <=  8'h77;        memory[6334] <=  8'h62;        memory[6335] <=  8'h65;        memory[6336] <=  8'h6e;        memory[6337] <=  8'h20;        memory[6338] <=  8'h6d;        memory[6339] <=  8'h64;        memory[6340] <=  8'h73;        memory[6341] <=  8'h6c;        memory[6342] <=  8'h76;        memory[6343] <=  8'h6b;        memory[6344] <=  8'h63;        memory[6345] <=  8'h78;        memory[6346] <=  8'h20;        memory[6347] <=  8'h6f;        memory[6348] <=  8'h78;        memory[6349] <=  8'h69;        memory[6350] <=  8'h63;        memory[6351] <=  8'h6a;        memory[6352] <=  8'h76;        memory[6353] <=  8'h64;        memory[6354] <=  8'h66;        memory[6355] <=  8'h65;        memory[6356] <=  8'h71;        memory[6357] <=  8'h6e;        memory[6358] <=  8'h20;        memory[6359] <=  8'h64;        memory[6360] <=  8'h6d;        memory[6361] <=  8'h73;        memory[6362] <=  8'h6c;        memory[6363] <=  8'h63;        memory[6364] <=  8'h78;        memory[6365] <=  8'h6b;        memory[6366] <=  8'h20;        memory[6367] <=  8'h6f;        memory[6368] <=  8'h78;        memory[6369] <=  8'h63;        memory[6370] <=  8'h76;        memory[6371] <=  8'h6a;        memory[6372] <=  8'h64;        memory[6373] <=  8'h62;        memory[6374] <=  8'h71;        memory[6375] <=  8'h77;        memory[6376] <=  8'h65;        memory[6377] <=  8'h6e;        memory[6378] <=  8'h6d;        memory[6379] <=  8'h64;        memory[6380] <=  8'h6c;        memory[6381] <=  8'h73;        memory[6382] <=  8'h2c;        memory[6383] <=  8'h76;        memory[6384] <=  8'h63;        memory[6385] <=  8'h78;        memory[6386] <=  8'h20;        memory[6387] <=  8'h63;        memory[6388] <=  8'h6f;        memory[6389] <=  8'h69;        memory[6390] <=  8'h76;        memory[6391] <=  8'h68;        memory[6392] <=  8'h73;        memory[6393] <=  8'h64;        memory[6394] <=  8'h62;        memory[6395] <=  8'h71;        memory[6396] <=  8'h77;        memory[6397] <=  8'h65;        memory[6398] <=  8'h6e;        memory[6399] <=  8'h64;        memory[6400] <=  8'h6b;        memory[6401] <=  8'h73;        memory[6402] <=  8'h76;        memory[6403] <=  8'h6f;        memory[6404] <=  8'h63;        memory[6405] <=  8'h20;        memory[6406] <=  8'h76;        memory[6407] <=  8'h69;        memory[6408] <=  8'h75;        memory[6409] <=  8'h69;        memory[6410] <=  8'h68;        memory[6411] <=  8'h63;        memory[6412] <=  8'h78;        memory[6413] <=  8'h69;        memory[6414] <=  8'h6f;        memory[6415] <=  8'h76;        memory[6416] <=  8'h73;        memory[6417] <=  8'h64;        memory[6418] <=  8'h61;        memory[6419] <=  8'h64;        memory[6420] <=  8'h6e;        memory[6421] <=  8'h77;        memory[6422] <=  8'h71;        memory[6423] <=  8'h6b;        memory[6424] <=  8'h6c;        memory[6425] <=  8'h73;        memory[6426] <=  8'h76;        memory[6427] <=  8'h6e;        memory[6428] <=  8'h62;        memory[6429] <=  8'h20;        memory[6430] <=  8'h64;        memory[6431] <=  8'h66;        memory[6432] <=  8'h6a;        memory[6433] <=  8'h6b;        memory[6434] <=  8'h71;        memory[6435] <=  8'h64;        memory[6436] <=  8'h77;        memory[6437] <=  8'h65;        memory[6438] <=  8'h6e;        memory[6439] <=  8'h62;        memory[6440] <=  8'h20;        memory[6441] <=  8'h64;        memory[6442] <=  8'h73;        memory[6443] <=  8'h76;        memory[6444] <=  8'h68;        memory[6445] <=  8'h64;        memory[6446] <=  8'h61;        memory[6447] <=  8'h71;        memory[6448] <=  8'h77;        memory[6449] <=  8'h6a;        memory[6450] <=  8'h65;        memory[6451] <=  8'h6e;        memory[6452] <=  8'h64;        memory[6453] <=  8'h20;        memory[6454] <=  8'h61;        memory[6455] <=  8'h63;        memory[6456] <=  8'h62;        memory[6457] <=  8'h68;        memory[6458] <=  8'h64;        memory[6459] <=  8'h61;        memory[6460] <=  8'h77;        memory[6461] <=  8'h71;        memory[6462] <=  8'h6e;        memory[6463] <=  8'h20;        memory[6464] <=  8'h62;        memory[6465] <=  8'h73;        memory[6466] <=  8'h76;        memory[6467] <=  8'h61;        memory[6468] <=  8'h67;        memory[6469] <=  8'h76;        memory[6470] <=  8'h68;        memory[6471] <=  8'h67;        memory[6472] <=  8'h61;        memory[6473] <=  8'h73;        memory[6474] <=  8'h6a;        memory[6475] <=  8'h6b;        memory[6476] <=  8'h63;        memory[6477] <=  8'h78;        memory[6478] <=  8'h76;        memory[6479] <=  8'h6e;        memory[6480] <=  8'h73;        memory[6481] <=  8'h64;        memory[6482] <=  8'h20;        memory[6483] <=  8'h66;        memory[6484] <=  8'h62;        memory[6485] <=  8'h64;        memory[6486] <=  8'h61;        memory[6487] <=  8'h73;        memory[6488] <=  8'h76;        memory[6489] <=  8'h67;        memory[6490] <=  8'h63;        memory[6491] <=  8'h79;        memory[6492] <=  8'h7a;        memory[6493] <=  8'h78;        memory[6494] <=  8'h79;        memory[6495] <=  8'h75;        memory[6496] <=  8'h20;        memory[6497] <=  8'h69;        memory[6498] <=  8'h6a;        memory[6499] <=  8'h64;        memory[6500] <=  8'h66;        memory[6501] <=  8'h6b;        memory[6502] <=  8'h61;        memory[6503] <=  8'h64;        memory[6504] <=  8'h63;        memory[6505] <=  8'h78;        memory[6506] <=  8'h68;        memory[6507] <=  8'h20;        memory[6508] <=  8'h67;        memory[6509] <=  8'h61;        memory[6510] <=  8'h68;        memory[6511] <=  8'h75;        memory[6512] <=  8'h64;        memory[6513] <=  8'h73;        memory[6514] <=  8'h69;        memory[6515] <=  8'h6a;        memory[6516] <=  8'h61;        memory[6517] <=  8'h6b;        memory[6518] <=  8'h63;        memory[6519] <=  8'h62;        memory[6520] <=  8'h61;        memory[6521] <=  8'h72;        memory[6522] <=  8'h73;        memory[6523] <=  8'h68;        memory[6524] <=  8'h64;        memory[6525] <=  8'h66;        memory[6526] <=  8'h67;        memory[6527] <=  8'h73;        memory[6528] <=  8'h68;        memory[6529] <=  8'h64;        memory[6530] <=  8'h66;        memory[6531] <=  8'h68;        memory[6532] <=  8'h64;        memory[6533] <=  8'h6a;        memory[6534] <=  8'h68;        memory[6535] <=  8'h62;        memory[6536] <=  8'h67;        memory[6537] <=  8'h63;        memory[6538] <=  8'h61;        memory[6539] <=  8'h66;        memory[6540] <=  8'h73;        memory[6541] <=  8'h79;        memory[6542] <=  8'h67;        memory[6543] <=  8'h6b;        memory[6544] <=  8'h75;        memory[6545] <=  8'h64;        memory[6546] <=  8'h68;        memory[6547] <=  8'h62;        memory[6548] <=  8'h77;        memory[6549] <=  8'h76;        memory[6550] <=  8'h67;        memory[6551] <=  8'h61;        memory[6552] <=  8'h66;        memory[6553] <=  8'h64;        memory[6554] <=  8'h74;        memory[6555] <=  8'h75;        memory[6556] <=  8'h66;        memory[6557] <=  8'h79;        memory[6558] <=  8'h67;        memory[6559] <=  8'h69;        memory[6560] <=  8'h75;        memory[6561] <=  8'h68;        memory[6562] <=  8'h6c;        memory[6563] <=  8'h6a;        memory[6564] <=  8'h62;        memory[6565] <=  8'h6b;        memory[6566] <=  8'h68;        memory[6567] <=  8'h76;        memory[6568] <=  8'h67;        memory[6569] <=  8'h63;        memory[6570] <=  8'h66;        memory[6571] <=  8'h78;        memory[6572] <=  8'h64;        memory[6573] <=  8'h74;        memory[6574] <=  8'h75;        memory[6575] <=  8'h79;        memory[6576] <=  8'h69;        memory[6577] <=  8'h75;        memory[6578] <=  8'h68;        memory[6579] <=  8'h6c;        memory[6580] <=  8'h6a;        memory[6581] <=  8'h6b;        memory[6582] <=  8'h67;        memory[6583] <=  8'h6a;        memory[6584] <=  8'h63;        memory[6585] <=  8'h66;        memory[6586] <=  8'h68;        memory[6587] <=  8'h64;        memory[6588] <=  8'h67;        memory[6589] <=  8'h72;        memory[6590] <=  8'h79;        memory[6591] <=  8'h74;        memory[6592] <=  8'h66;        memory[6593] <=  8'h75;        memory[6594] <=  8'h79;        memory[6595] <=  8'h69;        memory[6596] <=  8'h68;        memory[6597] <=  8'h6c;        memory[6598] <=  8'h62;        memory[6599] <=  8'h6d;        memory[6600] <=  8'h76;        memory[6601] <=  8'h6e;        memory[6602] <=  8'h63;        memory[6603] <=  8'h66;        memory[6604] <=  8'h68;        memory[6605] <=  8'h64;        memory[6606] <=  8'h74;        memory[6607] <=  8'h75;        memory[6608] <=  8'h67;        memory[6609] <=  8'h79;        memory[6610] <=  8'h69;        memory[6611] <=  8'h68;        memory[6612] <=  8'h75;        memory[6613] <=  8'h6a;        memory[6614] <=  8'h6c;        memory[6615] <=  8'h62;        memory[6616] <=  8'h6d;        memory[6617] <=  8'h76;        memory[6618] <=  8'h6e;        memory[6619] <=  8'h63;        memory[6620] <=  8'h66;        memory[6621] <=  8'h68;        memory[6622] <=  8'h67;        memory[6623] <=  8'h79;        memory[6624] <=  8'h68;        memory[6625] <=  8'h75;        memory[6626] <=  8'h6a;        memory[6627] <=  8'h6e;        memory[6628] <=  8'h2c;        memory[6629] <=  8'h62;        memory[6630] <=  8'h6e;        memory[6631] <=  8'h6d;        memory[6632] <=  8'h76;        memory[6633] <=  8'h6e;        memory[6634] <=  8'h63;        memory[6635] <=  8'h66;        memory[6636] <=  8'h68;        memory[6637] <=  8'h74;        memory[6638] <=  8'h79;        memory[6639] <=  8'h69;        memory[6640] <=  8'h75;        memory[6641] <=  8'h6c;        memory[6642] <=  8'h6a;        memory[6643] <=  8'h62;        memory[6644] <=  8'h6d;        memory[6645] <=  8'h76;        memory[6646] <=  8'h6e;        memory[6647] <=  8'h63;        memory[6648] <=  8'h66;        memory[6649] <=  8'h74;        memory[6650] <=  8'h75;        memory[6651] <=  8'h79;        memory[6652] <=  8'h69;        memory[6653] <=  8'h68;        memory[6654] <=  8'h6b;        memory[6655] <=  8'h62;        memory[6656] <=  8'h76;        memory[6657] <=  8'h63;        memory[6658] <=  8'h66;        memory[6659] <=  8'h67;        memory[6660] <=  8'h74;        memory[6661] <=  8'h75;        memory[6662] <=  8'h79;        memory[6663] <=  8'h69;        memory[6664] <=  8'h75;        memory[6665] <=  8'h68;        memory[6666] <=  8'h6a;        memory[6667] <=  8'h6b;        memory[6668] <=  8'h62;        memory[6669] <=  8'h76;        memory[6670] <=  8'h63;        memory[6671] <=  8'h66;        memory[6672] <=  8'h74;        memory[6673] <=  8'h75;        memory[6674] <=  8'h79;        memory[6675] <=  8'h69;        memory[6676] <=  8'h75;        memory[6677] <=  8'h6a;        memory[6678] <=  8'h6b;        memory[6679] <=  8'h6e;        memory[6680] <=  8'h62;        memory[6681] <=  8'h76;        memory[6682] <=  8'h67;        memory[6683] <=  8'h66;        memory[6684] <=  8'h74;        memory[6685] <=  8'h79;        memory[6686] <=  8'h75;        memory[6687] <=  8'h75;        memory[6688] <=  8'h69;        memory[6689] <=  8'h6a;        memory[6690] <=  8'h6b;        memory[6691] <=  8'h68;        memory[6692] <=  8'h62;        memory[6693] <=  8'h6a;        memory[6694] <=  8'h67;        memory[6695] <=  8'h68;        memory[6696] <=  8'h66;        memory[6697] <=  8'h79;        memory[6698] <=  8'h74;        memory[6699] <=  8'h79;        memory[6700] <=  8'h69;        memory[6701] <=  8'h75;        memory[6702] <=  8'h64;        memory[6703] <=  8'h6a;        memory[6704] <=  8'h6b;        memory[6705] <=  8'h68;        memory[6706] <=  8'h63;        memory[6707] <=  8'h7a;        memory[6708] <=  8'h67;        memory[6709] <=  8'h68;        memory[6710] <=  8'h74;        memory[6711] <=  8'h75;        memory[6712] <=  8'h79;        memory[6713] <=  8'h69;        memory[6714] <=  8'h61;        memory[6715] <=  8'h73;        memory[6716] <=  8'h75;        memory[6717] <=  8'h6a;        memory[6718] <=  8'h6b;        memory[6719] <=  8'h62;        memory[6720] <=  8'h6e;        memory[6721] <=  8'h61;        memory[6722] <=  8'h76;        memory[6723] <=  8'h63;        memory[6724] <=  8'h66;        memory[6725] <=  8'h68;        memory[6726] <=  8'h75;        memory[6727] <=  8'h61;        memory[6728] <=  8'h73;        memory[6729] <=  8'h79;        memory[6730] <=  8'h64;        memory[6731] <=  8'h75;        memory[6732] <=  8'h69;        memory[6733] <=  8'h6a;        memory[6734] <=  8'h61;        memory[6735] <=  8'h6b;        memory[6736] <=  8'h62;        memory[6737] <=  8'h63;        memory[6738] <=  8'h78;        memory[6739] <=  8'h68;        memory[6740] <=  8'h67;        memory[6741] <=  8'h79;        memory[6742] <=  8'h75;        memory[6743] <=  8'h7a;        memory[6744] <=  8'h63;        memory[6745] <=  8'h61;        memory[6746] <=  8'h73;        memory[6747] <=  8'h69;        memory[6748] <=  8'h75;        memory[6749] <=  8'h6f;        memory[6750] <=  8'h69;        memory[6751] <=  8'h6a;        memory[6752] <=  8'h61;        memory[6753] <=  8'h6c;        memory[6754] <=  8'h63;        memory[6755] <=  8'h78;        memory[6756] <=  8'h62;        memory[6757] <=  8'h63;        memory[6758] <=  8'h20;        memory[6759] <=  8'h6e;        memory[6760] <=  8'h76;        memory[6761] <=  8'h63;        memory[6762] <=  8'h61;        memory[6763] <=  8'h64;        memory[6764] <=  8'h73;        memory[6765] <=  8'h67;        memory[6766] <=  8'h79;        memory[6767] <=  8'h68;        memory[6768] <=  8'h75;        memory[6769] <=  8'h61;        memory[6770] <=  8'h6a;        memory[6771] <=  8'h6b;        memory[6772] <=  8'h78;        memory[6773] <=  8'h62;        memory[6774] <=  8'h20;        memory[6775] <=  8'h6e;        memory[6776] <=  8'h76;        memory[6777] <=  8'h63;        memory[6778] <=  8'h61;        memory[6779] <=  8'h73;        memory[6780] <=  8'h67;        memory[6781] <=  8'h68;        memory[6782] <=  8'h75;        memory[6783] <=  8'h6a;        memory[6784] <=  8'h6c;        memory[6785] <=  8'h6b;        memory[6786] <=  8'h63;        memory[6787] <=  8'h78;        memory[6788] <=  8'h20;        memory[6789] <=  8'h6a;        memory[6790] <=  8'h6b;        memory[6791] <=  8'h68;        memory[6792] <=  8'h61;        memory[6793] <=  8'h73;        memory[6794] <=  8'h76;        memory[6795] <=  8'h64;        memory[6796] <=  8'h6e;        memory[6797] <=  8'h20;        memory[6798] <=  8'h62;        memory[6799] <=  8'h6e;        memory[6800] <=  8'h6d;        memory[6801] <=  8'h6b;        memory[6802] <=  8'h77;        memory[6803] <=  8'h64;        memory[6804] <=  8'h6f;        memory[6805] <=  8'h77;        memory[6806] <=  8'h69;        memory[6807] <=  8'h6f;        memory[6808] <=  8'h75;        memory[6809] <=  8'h69;        memory[6810] <=  8'h68;        memory[6811] <=  8'h62;        memory[6812] <=  8'h6e;        memory[6813] <=  8'h6b;        memory[6814] <=  8'h77;        memory[6815] <=  8'h69;        memory[6816] <=  8'h6f;        memory[6817] <=  8'h75;        memory[6818] <=  8'h71;        memory[6819] <=  8'h69;        memory[6820] <=  8'h79;        memory[6821] <=  8'h67;        memory[6822] <=  8'h6a;        memory[6823] <=  8'h64;        memory[6824] <=  8'h61;        memory[6825] <=  8'h76;        memory[6826] <=  8'h62;        memory[6827] <=  8'h6e;        memory[6828] <=  8'h6b;        memory[6829] <=  8'h6f;        memory[6830] <=  8'h70;        memory[6831] <=  8'h64;        memory[6832] <=  8'h76;        memory[6833] <=  8'h69;        memory[6834] <=  8'h6f;        memory[6835] <=  8'h75;        memory[6836] <=  8'h69;        memory[6837] <=  8'h48;        memory[6838] <=  8'h42;        memory[6839] <=  8'h6b;        memory[6840] <=  8'h64;        memory[6841] <=  8'h6e;        memory[6842] <=  8'h6c;        memory[6843] <=  8'h71;        memory[6844] <=  8'h6b;        memory[6845] <=  8'h6d;        memory[6846] <=  8'h6a;        memory[6847] <=  8'h70;        memory[6848] <=  8'h69;        memory[6849] <=  8'h6f;        memory[6850] <=  8'h68;        memory[6851] <=  8'h65;        memory[6852] <=  8'h66;        memory[6853] <=  8'h75;        memory[6854] <=  8'h67;        memory[6855] <=  8'h69;        memory[6856] <=  8'h73;        memory[6857] <=  8'h61;        memory[6858] <=  8'h62;        memory[6859] <=  8'h64;        memory[6860] <=  8'h6b;        memory[6861] <=  8'h6a;        memory[6862] <=  8'h6b;        memory[6863] <=  8'h6c;        memory[6864] <=  8'h6a;        memory[6865] <=  8'h69;        memory[6866] <=  8'h73;        memory[6867] <=  8'h6f;        memory[6868] <=  8'h71;        memory[6869] <=  8'h68;        memory[6870] <=  8'h77;        memory[6871] <=  8'h67;        memory[6872] <=  8'h69;        memory[6873] <=  8'h79;        memory[6874] <=  8'h6a;        memory[6875] <=  8'h64;        memory[6876] <=  8'h76;        memory[6877] <=  8'h62;        memory[6878] <=  8'h6e;        memory[6879] <=  8'h61;        memory[6880] <=  8'h73;        memory[6881] <=  8'h66;        memory[6882] <=  8'h6c;        memory[6883] <=  8'h6b;        memory[6884] <=  8'h64;        memory[6885] <=  8'h6a;        memory[6886] <=  8'h68;        memory[6887] <=  8'h63;        memory[6888] <=  8'h67;        memory[6889] <=  8'h6a;        memory[6890] <=  8'h76;        memory[6891] <=  8'h73;        memory[6892] <=  8'h64;        memory[6893] <=  8'h62;        memory[6894] <=  8'h62;        memory[6895] <=  8'h61;        memory[6896] <=  8'h72;        memory[6897] <=  8'h62;        memory[6898] <=  8'h62;        memory[6899] <=  8'h73;        memory[6900] <=  8'h62;        memory[6901] <=  8'h67;        memory[6902] <=  8'h73;        memory[6903] <=  8'h66;        memory[6904] <=  8'h67;        memory[6905] <=  8'h61;        memory[6906] <=  8'h68;        memory[6907] <=  8'h66;        memory[6908] <=  8'h73;        memory[6909] <=  8'h68;        memory[6910] <=  8'h61;        memory[6911] <=  8'h66;        memory[6912] <=  8'h73;        memory[6913] <=  8'h66;        memory[6914] <=  8'h68;        memory[6915] <=  8'h61;        memory[6916] <=  8'h69;        memory[6917] <=  8'h64;        memory[6918] <=  8'h75;        memory[6919] <=  8'h67;        memory[6920] <=  8'h64;        memory[6921] <=  8'h77;        memory[6922] <=  8'h62;        memory[6923] <=  8'h61;        memory[6924] <=  8'h62;        memory[6925] <=  8'h72;        memory[6926] <=  8'h62;        memory[6927] <=  8'h61;        memory[6928] <=  8'h62;        memory[6929] <=  8'h62;        memory[6930] <=  8'h74;        memory[6931] <=  8'h62;        memory[6932] <=  8'h62;        memory[6933] <=  8'h62;        memory[6934] <=  8'h62;        memory[6935] <=  8'h62;        memory[6936] <=  8'h62;        memory[6937] <=  8'h62;        memory[6938] <=  8'h62;        memory[6939] <=  8'h61;        memory[6940] <=  8'h62;        memory[6941] <=  8'h62;        memory[6942] <=  8'h72;        memory[6943] <=  8'h74;        memory[6944] <=  8'h62;        memory[6945] <=  8'h62;        memory[6946] <=  8'h61;        memory[6947] <=  8'h62;        memory[6948] <=  8'h72;        memory[6949] <=  8'h62;        memory[6950] <=  8'h74;        memory[6951] <=  8'h62;        memory[6952] <=  8'h62;        memory[6953] <=  8'h62;        memory[6954] <=  8'h63;        memory[6955] <=  8'h61;        memory[6956] <=  8'h72;        memory[6957] <=  8'h74;        memory[6958] <=  8'h73;        memory[6959] <=  8'h62;        memory[6960] <=  8'h61;        memory[6961] <=  8'h72;        memory[6962] <=  8'h74;        memory[6963] <=  8'h74;        memory[6964] <=  8'h62;        memory[6965] <=  8'h61;        memory[6966] <=  8'h72;        memory[6967] <=  8'h74;        memory[6968] <=  8'h78;        memory[6969] <=  8'h61;        memory[6970] <=  8'h74;        memory[6971] <=  8'h6b;        memory[6972] <=  8'h73;        memory[6973] <=  8'h68;        memory[6974] <=  8'h63;        memory[6975] <=  8'h66;        memory[6976] <=  8'h69;        memory[6977] <=  8'h77;        memory[6978] <=  8'h68;        memory[6979] <=  8'h61;        memory[6980] <=  8'h74;        memory[6981] <=  8'h61;        memory[6982] <=  8'h6e;        memory[6983] <=  8'h61;        memory[6984] <=  8'h62;        memory[6985] <=  8'h61;        memory[6986] <=  8'h63;        memory[6987] <=  8'h61;        memory[6988] <=  8'h74;        memory[6989] <=  8'h61;        memory[6990] <=  8'h62;        memory[6991] <=  8'h61;        memory[6992] <=  8'h72;        memory[6993] <=  8'h63;        memory[6994] <=  8'h61;        memory[6995] <=  8'h68;        memory[6996] <=  8'h64;        memory[6997] <=  8'h75;        memory[6998] <=  8'h63;        memory[6999] <=  8'h74;        memory[7000] <=  8'h61;        memory[7001] <=  8'h64;        memory[7002] <=  8'h61;        memory[7003] <=  8'h61;        memory[7004] <=  8'h63;        memory[7005] <=  8'h61;        memory[7006] <=  8'h72;        memory[7007] <=  8'h63;        memory[7008] <=  8'h74;        memory[7009] <=  8'h72;        memory[7010] <=  8'h63;        memory[7011] <=  8'h61;        memory[7012] <=  8'h74;        memory[7013] <=  8'h72;        memory[7014] <=  8'h63;        memory[7015] <=  8'h61;        memory[7016] <=  8'h74;        memory[7017] <=  8'h63;        memory[7018] <=  8'h62;        memory[7019] <=  8'h61;        memory[7020] <=  8'h74;        memory[7021] <=  8'h62;        memory[7022] <=  8'h72;        memory[7023] <=  8'h63;        memory[7024] <=  8'h61;        memory[7025] <=  8'h74;        memory[7026] <=  8'h72;        memory[7027] <=  8'h6e;        memory[7028] <=  8'h62;        memory[7029] <=  8'h61;        memory[7030] <=  8'h63;        memory[7031] <=  8'h61;        memory[7032] <=  8'h74;        memory[7033] <=  8'h79;        memory[7034] <=  8'h73;        memory[7035] <=  8'h6e;        memory[7036] <=  8'h63;        memory[7037] <=  8'h74;        memory[7038] <=  8'h61;        memory[7039] <=  8'h6e;        memory[7040] <=  8'h62;        memory[7041] <=  8'h61;        memory[7042] <=  8'h63;        memory[7043] <=  8'h72;        memory[7044] <=  8'h6e;        memory[7045] <=  8'h74;        memory[7046] <=  8'h61;        memory[7047] <=  8'h62;        memory[7048] <=  8'h74;        memory[7049] <=  8'h6e;        memory[7050] <=  8'h61;        memory[7051] <=  8'h72;        memory[7052] <=  8'h62;        memory[7053] <=  8'h78;        memory[7054] <=  8'h74;        memory[7055] <=  8'h61;        memory[7056] <=  8'h72;        memory[7057] <=  8'h62;        memory[7058] <=  8'h61;        memory[7059] <=  8'h72;        memory[7060] <=  8'h74;        memory[7061] <=  8'h74;        memory[7062] <=  8'h62;        memory[7063] <=  8'h61;        memory[7064] <=  8'h72;        memory[7065] <=  8'h74;        memory[7066] <=  8'h78;        memory[7067] <=  8'h61;        memory[7068] <=  8'h74;        memory[7069] <=  8'h6b;        memory[7070] <=  8'h73;        memory[7071] <=  8'h68;        memory[7072] <=  8'h63;        memory[7073] <=  8'h66;        memory[7074] <=  8'h69;        memory[7075] <=  8'h77;        memory[7076] <=  8'h68;        memory[7077] <=  8'h61;        memory[7078] <=  8'h74;        memory[7079] <=  8'h61;        memory[7080] <=  8'h6e;        memory[7081] <=  8'h61;        memory[7082] <=  8'h62;        memory[7083] <=  8'h61;        memory[7084] <=  8'h63;        memory[7085] <=  8'h61;        memory[7086] <=  8'h74;        memory[7087] <=  8'h61;        memory[7088] <=  8'h62;        memory[7089] <=  8'h61;        memory[7090] <=  8'h72;        memory[7091] <=  8'h63;        memory[7092] <=  8'h61;        memory[7093] <=  8'h68;        memory[7094] <=  8'h64;        memory[7095] <=  8'h75;        memory[7096] <=  8'h63;        memory[7097] <=  8'h74;        memory[7098] <=  8'h61;        memory[7099] <=  8'h64;        memory[7100] <=  8'h61;        memory[7101] <=  8'h61;        memory[7102] <=  8'h63;        memory[7103] <=  8'h61;        memory[7104] <=  8'h72;        memory[7105] <=  8'h63;        memory[7106] <=  8'h74;        memory[7107] <=  8'h72;        memory[7108] <=  8'h63;        memory[7109] <=  8'h61;        memory[7110] <=  8'h74;        memory[7111] <=  8'h72;        memory[7112] <=  8'h63;        memory[7113] <=  8'h61;        memory[7114] <=  8'h74;        memory[7115] <=  8'h63;        memory[7116] <=  8'h62;        memory[7117] <=  8'h61;        memory[7118] <=  8'h74;        memory[7119] <=  8'h62;        memory[7120] <=  8'h72;        memory[7121] <=  8'h63;        memory[7122] <=  8'h61;        memory[7123] <=  8'h74;        memory[7124] <=  8'h72;        memory[7125] <=  8'h6e;        memory[7126] <=  8'h62;        memory[7127] <=  8'h61;        memory[7128] <=  8'h63;        memory[7129] <=  8'h61;        memory[7130] <=  8'h74;        memory[7131] <=  8'h79;        memory[7132] <=  8'h73;        memory[7133] <=  8'h6e;        memory[7134] <=  8'h63;        memory[7135] <=  8'h74;        memory[7136] <=  8'h61;        memory[7137] <=  8'h6e;        memory[7138] <=  8'h62;        memory[7139] <=  8'h61;        memory[7140] <=  8'h63;        memory[7141] <=  8'h72;        memory[7142] <=  8'h6e;        memory[7143] <=  8'h74;        memory[7144] <=  8'h61;        memory[7145] <=  8'h62;        memory[7146] <=  8'h74;        memory[7147] <=  8'h6e;        memory[7148] <=  8'h61;        memory[7149] <=  8'h72;        memory[7150] <=  8'h62;        memory[7151] <=  8'h78;        memory[7152] <=  8'h74;        memory[7153] <=  8'h61;        memory[7154] <=  8'h72;        memory[7155] <=  8'h62;        memory[7156] <=  8'h61;        memory[7157] <=  8'h72;        memory[7158] <=  8'h74;        memory[7159] <=  8'h74;        memory[7160] <=  8'h62;        memory[7161] <=  8'h61;        memory[7162] <=  8'h72;        memory[7163] <=  8'h74;        memory[7164] <=  8'h78;        memory[7165] <=  8'h61;        memory[7166] <=  8'h74;        memory[7167] <=  8'h6b;        memory[7168] <=  8'h73;        memory[7169] <=  8'h68;        memory[7170] <=  8'h63;        memory[7171] <=  8'h66;        memory[7172] <=  8'h69;        memory[7173] <=  8'h77;        memory[7174] <=  8'h68;        memory[7175] <=  8'h61;        memory[7176] <=  8'h74;        memory[7177] <=  8'h61;        memory[7178] <=  8'h6e;        memory[7179] <=  8'h61;        memory[7180] <=  8'h62;        memory[7181] <=  8'h61;        memory[7182] <=  8'h63;        memory[7183] <=  8'h61;        memory[7184] <=  8'h74;        memory[7185] <=  8'h61;        memory[7186] <=  8'h62;        memory[7187] <=  8'h61;        memory[7188] <=  8'h72;        memory[7189] <=  8'h63;        memory[7190] <=  8'h61;        memory[7191] <=  8'h68;        memory[7192] <=  8'h64;        memory[7193] <=  8'h75;        memory[7194] <=  8'h63;        memory[7195] <=  8'h74;        memory[7196] <=  8'h61;        memory[7197] <=  8'h64;        memory[7198] <=  8'h61;        memory[7199] <=  8'h61;        memory[7200] <=  8'h63;        memory[7201] <=  8'h61;        memory[7202] <=  8'h72;        memory[7203] <=  8'h63;        memory[7204] <=  8'h74;        memory[7205] <=  8'h72;        memory[7206] <=  8'h63;        memory[7207] <=  8'h61;        memory[7208] <=  8'h74;        memory[7209] <=  8'h72;        memory[7210] <=  8'h63;        memory[7211] <=  8'h61;        memory[7212] <=  8'h74;        memory[7213] <=  8'h63;        memory[7214] <=  8'h62;        memory[7215] <=  8'h61;        memory[7216] <=  8'h74;        memory[7217] <=  8'h62;        memory[7218] <=  8'h72;        memory[7219] <=  8'h63;        memory[7220] <=  8'h61;        memory[7221] <=  8'h74;        memory[7222] <=  8'h72;        memory[7223] <=  8'h6e;        memory[7224] <=  8'h62;        memory[7225] <=  8'h61;        memory[7226] <=  8'h63;        memory[7227] <=  8'h61;        memory[7228] <=  8'h74;        memory[7229] <=  8'h79;        memory[7230] <=  8'h73;        memory[7231] <=  8'h6e;        memory[7232] <=  8'h63;        memory[7233] <=  8'h74;        memory[7234] <=  8'h61;        memory[7235] <=  8'h6e;        memory[7236] <=  8'h62;        memory[7237] <=  8'h61;        memory[7238] <=  8'h63;        memory[7239] <=  8'h72;        memory[7240] <=  8'h6e;        memory[7241] <=  8'h74;        memory[7242] <=  8'h61;        memory[7243] <=  8'h62;        memory[7244] <=  8'h74;        memory[7245] <=  8'h6e;        memory[7246] <=  8'h61;        memory[7247] <=  8'h72;        memory[7248] <=  8'h62;        memory[7249] <=  8'h78;        memory[7250] <=  8'h74;        memory[7251] <=  8'h61;        memory[7252] <=  8'h72;        memory[7253] <=  8'h5d;        memory[7254] <=  8'h5d;        memory[7255] <=  8'h65;        memory[7256] <=  8'h66;        memory[7257] <=  8'h77;        memory[7258] <=  8'h65;        memory[7259] <=  8'h5d;        memory[7260] <=  8'h65;        memory[7261] <=  8'h67;        memory[7262] <=  8'h73;        memory[7263] <=  8'h67;        memory[7264] <=  8'h66;        memory[7265] <=  8'h62;        memory[7266] <=  8'h61;        memory[7267] <=  8'h72;        memory[7268] <=  8'h74;        memory[7269] <=  8'h74;        memory[7270] <=  8'h62;        memory[7271] <=  8'h61;        memory[7272] <=  8'h72;        memory[7273] <=  8'h74;        memory[7274] <=  8'h78;        memory[7275] <=  8'h61;        memory[7276] <=  8'h74;        memory[7277] <=  8'h6b;        memory[7278] <=  8'h73;        memory[7279] <=  8'h68;        memory[7280] <=  8'h63;        memory[7281] <=  8'h66;        memory[7282] <=  8'h69;        memory[7283] <=  8'h77;        memory[7284] <=  8'h68;        memory[7285] <=  8'h61;        memory[7286] <=  8'h74;        memory[7287] <=  8'h61;        memory[7288] <=  8'h6e;        memory[7289] <=  8'h61;        memory[7290] <=  8'h62;        memory[7291] <=  8'h61;        memory[7292] <=  8'h63;        memory[7293] <=  8'h61;        memory[7294] <=  8'h74;        memory[7295] <=  8'h61;        memory[7296] <=  8'h62;        memory[7297] <=  8'h61;        memory[7298] <=  8'h72;        memory[7299] <=  8'h63;        memory[7300] <=  8'h61;        memory[7301] <=  8'h68;        memory[7302] <=  8'h64;        memory[7303] <=  8'h75;        memory[7304] <=  8'h63;        memory[7305] <=  8'h74;        memory[7306] <=  8'h61;        memory[7307] <=  8'h64;        memory[7308] <=  8'h61;        memory[7309] <=  8'h61;        memory[7310] <=  8'h63;        memory[7311] <=  8'h61;        memory[7312] <=  8'h72;        memory[7313] <=  8'h63;        memory[7314] <=  8'h74;        memory[7315] <=  8'h72;        memory[7316] <=  8'h63;        memory[7317] <=  8'h61;        memory[7318] <=  8'h74;        memory[7319] <=  8'h72;        memory[7320] <=  8'h63;        memory[7321] <=  8'h61;        memory[7322] <=  8'h74;        memory[7323] <=  8'h63;        memory[7324] <=  8'h62;        memory[7325] <=  8'h61;        memory[7326] <=  8'h74;        memory[7327] <=  8'h62;        memory[7328] <=  8'h72;        memory[7329] <=  8'h63;        memory[7330] <=  8'h61;        memory[7331] <=  8'h74;        memory[7332] <=  8'h72;        memory[7333] <=  8'h6e;        memory[7334] <=  8'h62;        memory[7335] <=  8'h61;        memory[7336] <=  8'h63;        memory[7337] <=  8'h61;        memory[7338] <=  8'h74;        memory[7339] <=  8'h79;        memory[7340] <=  8'h73;        memory[7341] <=  8'h6e;        memory[7342] <=  8'h63;        memory[7343] <=  8'h74;        memory[7344] <=  8'h61;        memory[7345] <=  8'h6e;        memory[7346] <=  8'h62;        memory[7347] <=  8'h61;        memory[7348] <=  8'h63;        memory[7349] <=  8'h72;        memory[7350] <=  8'h6e;        memory[7351] <=  8'h74;        memory[7352] <=  8'h61;        memory[7353] <=  8'h62;        memory[7354] <=  8'h74;        memory[7355] <=  8'h6e;        memory[7356] <=  8'h61;        memory[7357] <=  8'h72;        memory[7358] <=  8'h62;        memory[7359] <=  8'h78;        memory[7360] <=  8'h74;        memory[7361] <=  8'h61;        memory[7362] <=  8'h72;        memory[7363] <=  8'h62;        memory[7364] <=  8'h61;        memory[7365] <=  8'h72;        memory[7366] <=  8'h74;        memory[7367] <=  8'h74;        memory[7368] <=  8'h62;        memory[7369] <=  8'h61;        memory[7370] <=  8'h72;        memory[7371] <=  8'h74;        memory[7372] <=  8'h78;        memory[7373] <=  8'h61;        memory[7374] <=  8'h74;        memory[7375] <=  8'h6b;        memory[7376] <=  8'h73;        memory[7377] <=  8'h68;        memory[7378] <=  8'h63;        memory[7379] <=  8'h66;        memory[7380] <=  8'h69;        memory[7381] <=  8'h77;        memory[7382] <=  8'h68;        memory[7383] <=  8'h61;        memory[7384] <=  8'h74;        memory[7385] <=  8'h61;        memory[7386] <=  8'h6e;        memory[7387] <=  8'h61;        memory[7388] <=  8'h62;        memory[7389] <=  8'h61;        memory[7390] <=  8'h63;        memory[7391] <=  8'h61;        memory[7392] <=  8'h74;        memory[7393] <=  8'h61;        memory[7394] <=  8'h62;        memory[7395] <=  8'h61;        memory[7396] <=  8'h72;        memory[7397] <=  8'h63;        memory[7398] <=  8'h61;        memory[7399] <=  8'h68;        memory[7400] <=  8'h64;        memory[7401] <=  8'h75;        memory[7402] <=  8'h63;        memory[7403] <=  8'h74;        memory[7404] <=  8'h61;        memory[7405] <=  8'h64;        memory[7406] <=  8'h61;        memory[7407] <=  8'h61;        memory[7408] <=  8'h63;        memory[7409] <=  8'h61;        memory[7410] <=  8'h72;        memory[7411] <=  8'h63;        memory[7412] <=  8'h74;        memory[7413] <=  8'h72;        memory[7414] <=  8'h63;        memory[7415] <=  8'h61;        memory[7416] <=  8'h74;        memory[7417] <=  8'h72;        memory[7418] <=  8'h63;        memory[7419] <=  8'h61;        memory[7420] <=  8'h74;        memory[7421] <=  8'h63;        memory[7422] <=  8'h62;        memory[7423] <=  8'h61;        memory[7424] <=  8'h74;        memory[7425] <=  8'h62;        memory[7426] <=  8'h72;        memory[7427] <=  8'h63;        memory[7428] <=  8'h61;        memory[7429] <=  8'h74;        memory[7430] <=  8'h72;        memory[7431] <=  8'h6e;        memory[7432] <=  8'h62;        memory[7433] <=  8'h61;        memory[7434] <=  8'h63;        memory[7435] <=  8'h61;        memory[7436] <=  8'h74;        memory[7437] <=  8'h79;        memory[7438] <=  8'h73;        memory[7439] <=  8'h6e;        memory[7440] <=  8'h63;        memory[7441] <=  8'h74;        memory[7442] <=  8'h61;        memory[7443] <=  8'h6e;        memory[7444] <=  8'h62;        memory[7445] <=  8'h61;        memory[7446] <=  8'h63;        memory[7447] <=  8'h72;        memory[7448] <=  8'h6e;        memory[7449] <=  8'h74;        memory[7450] <=  8'h61;        memory[7451] <=  8'h62;        memory[7452] <=  8'h74;        memory[7453] <=  8'h6e;        memory[7454] <=  8'h61;        memory[7455] <=  8'h72;        memory[7456] <=  8'h62;        memory[7457] <=  8'h78;        memory[7458] <=  8'h74;        memory[7459] <=  8'h61;        memory[7460] <=  8'h72;        memory[7461] <=  8'h64;        memory[7462] <=  8'h66;        memory[7463] <=  8'h73;        memory[7464] <=  8'h67;        memory[7465] <=  8'h76;        memory[7466] <=  8'h68;        memory[7467] <=  8'h62;        memory[7468] <=  8'h6b;        memory[7469] <=  8'h6a;        memory[7470] <=  8'h6e;        memory[7471] <=  8'h6d;        memory[7472] <=  8'h62;        memory[7473] <=  8'h76;        memory[7474] <=  8'h78;        memory[7475] <=  8'h63;        memory[7476] <=  8'h73;        memory[7477] <=  8'h66;        memory[7478] <=  8'h72;        memory[7479] <=  8'h74;        memory[7480] <=  8'h79;        memory[7481] <=  8'h75;        memory[7482] <=  8'h6a;        memory[7483] <=  8'h6e;        memory[7484] <=  8'h62;        memory[7485] <=  8'h76;        memory[7486] <=  8'h63;        memory[7487] <=  8'h64;        memory[7488] <=  8'h74;        memory[7489] <=  8'h79;        memory[7490] <=  8'h75;        memory[7491] <=  8'h69;        memory[7492] <=  8'h6b;        memory[7493] <=  8'h6d;        memory[7494] <=  8'h6e;        memory[7495] <=  8'h62;        memory[7496] <=  8'h76;        memory[7497] <=  8'h63;        memory[7498] <=  8'h78;        memory[7499] <=  8'h73;        memory[7500] <=  8'h64;        memory[7501] <=  8'h72;        memory[7502] <=  8'h74;        memory[7503] <=  8'h79;        memory[7504] <=  8'h75;        memory[7505] <=  8'h69;        memory[7506] <=  8'h6b;        memory[7507] <=  8'h6d;        memory[7508] <=  8'h6e;        memory[7509] <=  8'h62;        memory[7510] <=  8'h76;        memory[7511] <=  8'h63;        memory[7512] <=  8'h73;        memory[7513] <=  8'h77;        memory[7514] <=  8'h33;        memory[7515] <=  8'h34;        memory[7516] <=  8'h35;        memory[7517] <=  8'h36;        memory[7518] <=  8'h37;        memory[7519] <=  8'h38;        memory[7520] <=  8'h69;        memory[7521] <=  8'h6b;        memory[7522] <=  8'h6d;        memory[7523] <=  8'h6e;        memory[7524] <=  8'h62;        memory[7525] <=  8'h76;        memory[7526] <=  8'h63;        memory[7527] <=  8'h64;        memory[7528] <=  8'h65;        memory[7529] <=  8'h72;        memory[7530] <=  8'h36;        memory[7531] <=  8'h37;        memory[7532] <=  8'h38;        memory[7533] <=  8'h69;        memory[7534] <=  8'h6f;        memory[7535] <=  8'h6b;        memory[7536] <=  8'h6a;        memory[7537] <=  8'h6e;        memory[7538] <=  8'h62;        memory[7539] <=  8'h76;        memory[7540] <=  8'h63;        memory[7541] <=  8'h64;        memory[7542] <=  8'h72;        memory[7543] <=  8'h74;        memory[7544] <=  8'h79;        memory[7545] <=  8'h75;        memory[7546] <=  8'h73;        memory[7547] <=  8'h6a;        memory[7548] <=  8'h63;        memory[7549] <=  8'h6e;        memory[7550] <=  8'h62;        memory[7551] <=  8'h64;        memory[7552] <=  8'h66;        memory[7553] <=  8'h73;        memory[7554] <=  8'h74;        memory[7555] <=  8'h79;        memory[7556] <=  8'h75;        memory[7557] <=  8'h61;        memory[7558] <=  8'h69;        memory[7559] <=  8'h6b;        memory[7560] <=  8'h78;        memory[7561] <=  8'h6d;        memory[7562] <=  8'h6e;        memory[7563] <=  8'h73;        memory[7564] <=  8'h6a;        memory[7565] <=  8'h6f;        memory[7566] <=  8'h64;        memory[7567] <=  8'h6c;        memory[7568] <=  8'h63;        memory[7569] <=  8'h78;        memory[7570] <=  8'h62;        memory[7571] <=  8'h61;        memory[7572] <=  8'h72;        memory[7573] <=  8'h74;        memory[7574] <=  8'h78;        memory[7575] <=  8'h61;        memory[7576] <=  8'h74;        memory[7577] <=  8'h6b;        memory[7578] <=  8'h73;        memory[7579] <=  8'h68;        memory[7580] <=  8'h63;        memory[7581] <=  8'h66;        memory[7582] <=  8'h69;        memory[7583] <=  8'h77;        memory[7584] <=  8'h68;        memory[7585] <=  8'h61;        memory[7586] <=  8'h74;        memory[7587] <=  8'h61;        memory[7588] <=  8'h6e;        memory[7589] <=  8'h61;        memory[7590] <=  8'h62;        memory[7591] <=  8'h61;        memory[7592] <=  8'h63;        memory[7593] <=  8'h61;        memory[7594] <=  8'h74;        memory[7595] <=  8'h61;        memory[7596] <=  8'h62;        memory[7597] <=  8'h61;        memory[7598] <=  8'h72;        memory[7599] <=  8'h63;        memory[7600] <=  8'h61;        memory[7601] <=  8'h68;        memory[7602] <=  8'h64;        memory[7603] <=  8'h75;        memory[7604] <=  8'h63;        memory[7605] <=  8'h74;        memory[7606] <=  8'h61;        memory[7607] <=  8'h64;        memory[7608] <=  8'h61;        memory[7609] <=  8'h61;        memory[7610] <=  8'h63;        memory[7611] <=  8'h61;        memory[7612] <=  8'h72;        memory[7613] <=  8'h62;        memory[7614] <=  8'h61;        memory[7615] <=  8'h72;        memory[7616] <=  8'h74;        memory[7617] <=  8'h78;        memory[7618] <=  8'h61;        memory[7619] <=  8'h74;        memory[7620] <=  8'h6b;        memory[7621] <=  8'h73;        memory[7622] <=  8'h68;        memory[7623] <=  8'h63;        memory[7624] <=  8'h66;        memory[7625] <=  8'h69;        memory[7626] <=  8'h77;        memory[7627] <=  8'h68;        memory[7628] <=  8'h61;        memory[7629] <=  8'h74;        memory[7630] <=  8'h61;        memory[7631] <=  8'h6e;        memory[7632] <=  8'h61;        memory[7633] <=  8'h62;        memory[7634] <=  8'h61;        memory[7635] <=  8'h63;        memory[7636] <=  8'h61;        memory[7637] <=  8'h74;        memory[7638] <=  8'h61;        memory[7639] <=  8'h62;        memory[7640] <=  8'h61;        memory[7641] <=  8'h72;        memory[7642] <=  8'h63;        memory[7643] <=  8'h61;        memory[7644] <=  8'h68;        memory[7645] <=  8'h64;        memory[7646] <=  8'h75;        memory[7647] <=  8'h63;        memory[7648] <=  8'h74;        memory[7649] <=  8'h61;        memory[7650] <=  8'h64;        memory[7651] <=  8'h61;        memory[7652] <=  8'h61;        memory[7653] <=  8'h63;        memory[7654] <=  8'h61;        memory[7655] <=  8'h72;        memory[7656] <=  8'h62;        memory[7657] <=  8'h61;        memory[7658] <=  8'h72;        memory[7659] <=  8'h74;        memory[7660] <=  8'h78;        memory[7661] <=  8'h61;        memory[7662] <=  8'h74;        memory[7663] <=  8'h6b;        memory[7664] <=  8'h73;        memory[7665] <=  8'h68;        memory[7666] <=  8'h63;        memory[7667] <=  8'h66;        memory[7668] <=  8'h69;        memory[7669] <=  8'h77;        memory[7670] <=  8'h68;        memory[7671] <=  8'h61;        memory[7672] <=  8'h74;        memory[7673] <=  8'h61;        memory[7674] <=  8'h6e;        memory[7675] <=  8'h61;        memory[7676] <=  8'h62;        memory[7677] <=  8'h61;        memory[7678] <=  8'h63;        memory[7679] <=  8'h61;        memory[7680] <=  8'h74;        memory[7681] <=  8'h61;        memory[7682] <=  8'h62;        memory[7683] <=  8'h61;        memory[7684] <=  8'h72;        memory[7685] <=  8'h63;        memory[7686] <=  8'h61;        memory[7687] <=  8'h68;        memory[7688] <=  8'h64;        memory[7689] <=  8'h75;        memory[7690] <=  8'h63;        memory[7691] <=  8'h74;        memory[7692] <=  8'h61;        memory[7693] <=  8'h64;        memory[7694] <=  8'h61;        memory[7695] <=  8'h61;        memory[7696] <=  8'h63;        memory[7697] <=  8'h61;        memory[7698] <=  8'h72;        memory[7699] <=  8'h62;        memory[7700] <=  8'h61;        memory[7701] <=  8'h72;        memory[7702] <=  8'h74;        memory[7703] <=  8'h78;        memory[7704] <=  8'h61;        memory[7705] <=  8'h74;        memory[7706] <=  8'h6b;        memory[7707] <=  8'h73;        memory[7708] <=  8'h68;        memory[7709] <=  8'h63;        memory[7710] <=  8'h66;        memory[7711] <=  8'h69;        memory[7712] <=  8'h77;        memory[7713] <=  8'h68;        memory[7714] <=  8'h61;        memory[7715] <=  8'h74;        memory[7716] <=  8'h61;        memory[7717] <=  8'h6e;        memory[7718] <=  8'h61;        memory[7719] <=  8'h62;        memory[7720] <=  8'h61;        memory[7721] <=  8'h63;        memory[7722] <=  8'h61;        memory[7723] <=  8'h74;        memory[7724] <=  8'h61;        memory[7725] <=  8'h62;        memory[7726] <=  8'h61;        memory[7727] <=  8'h72;        memory[7728] <=  8'h63;        memory[7729] <=  8'h61;        memory[7730] <=  8'h68;        memory[7731] <=  8'h64;        memory[7732] <=  8'h75;        memory[7733] <=  8'h63;        memory[7734] <=  8'h74;        memory[7735] <=  8'h61;        memory[7736] <=  8'h64;        memory[7737] <=  8'h61;        memory[7738] <=  8'h61;        memory[7739] <=  8'h63;        memory[7740] <=  8'h61;        memory[7741] <=  8'h72;        memory[7742] <=  8'h62;        memory[7743] <=  8'h61;        memory[7744] <=  8'h72;        memory[7745] <=  8'h74;        memory[7746] <=  8'h78;        memory[7747] <=  8'h61;        memory[7748] <=  8'h74;        memory[7749] <=  8'h6b;        memory[7750] <=  8'h73;        memory[7751] <=  8'h68;        memory[7752] <=  8'h63;        memory[7753] <=  8'h66;        memory[7754] <=  8'h69;        memory[7755] <=  8'h77;        memory[7756] <=  8'h68;        memory[7757] <=  8'h61;        memory[7758] <=  8'h74;        memory[7759] <=  8'h61;        memory[7760] <=  8'h6e;        memory[7761] <=  8'h61;        memory[7762] <=  8'h62;        memory[7763] <=  8'h61;        memory[7764] <=  8'h63;        memory[7765] <=  8'h61;        memory[7766] <=  8'h74;        memory[7767] <=  8'h61;        memory[7768] <=  8'h62;        memory[7769] <=  8'h61;        memory[7770] <=  8'h72;        memory[7771] <=  8'h63;        memory[7772] <=  8'h61;        memory[7773] <=  8'h68;        memory[7774] <=  8'h64;        memory[7775] <=  8'h75;        memory[7776] <=  8'h63;        memory[7777] <=  8'h74;        memory[7778] <=  8'h61;        memory[7779] <=  8'h64;        memory[7780] <=  8'h61;        memory[7781] <=  8'h61;        memory[7782] <=  8'h63;        memory[7783] <=  8'h61;        memory[7784] <=  8'h72;        memory[7785] <=  8'h62;        memory[7786] <=  8'h61;        memory[7787] <=  8'h72;        memory[7788] <=  8'h74;        memory[7789] <=  8'h78;        memory[7790] <=  8'h61;        memory[7791] <=  8'h74;        memory[7792] <=  8'h6b;        memory[7793] <=  8'h73;        memory[7794] <=  8'h68;        memory[7795] <=  8'h63;        memory[7796] <=  8'h66;        memory[7797] <=  8'h69;        memory[7798] <=  8'h77;        memory[7799] <=  8'h68;        memory[7800] <=  8'h61;        memory[7801] <=  8'h74;        memory[7802] <=  8'h61;        memory[7803] <=  8'h6e;        memory[7804] <=  8'h61;        memory[7805] <=  8'h62;        memory[7806] <=  8'h61;        memory[7807] <=  8'h63;        memory[7808] <=  8'h61;        memory[7809] <=  8'h74;        memory[7810] <=  8'h61;        memory[7811] <=  8'h62;        memory[7812] <=  8'h61;        memory[7813] <=  8'h72;        memory[7814] <=  8'h63;        memory[7815] <=  8'h61;        memory[7816] <=  8'h68;        memory[7817] <=  8'h64;        memory[7818] <=  8'h75;        memory[7819] <=  8'h63;        memory[7820] <=  8'h74;        memory[7821] <=  8'h61;        memory[7822] <=  8'h64;        memory[7823] <=  8'h61;        memory[7824] <=  8'h61;        memory[7825] <=  8'h63;        memory[7826] <=  8'h61;        memory[7827] <=  8'h72;        memory[7828] <=  8'h62;        memory[7829] <=  8'h61;        memory[7830] <=  8'h72;        memory[7831] <=  8'h74;        memory[7832] <=  8'h78;        memory[7833] <=  8'h61;        memory[7834] <=  8'h74;        memory[7835] <=  8'h6b;        memory[7836] <=  8'h73;        memory[7837] <=  8'h68;        memory[7838] <=  8'h63;        memory[7839] <=  8'h66;        memory[7840] <=  8'h69;        memory[7841] <=  8'h77;        memory[7842] <=  8'h68;        memory[7843] <=  8'h61;        memory[7844] <=  8'h74;        memory[7845] <=  8'h61;        memory[7846] <=  8'h6e;        memory[7847] <=  8'h61;        memory[7848] <=  8'h62;        memory[7849] <=  8'h61;        memory[7850] <=  8'h63;        memory[7851] <=  8'h61;        memory[7852] <=  8'h74;        memory[7853] <=  8'h61;        memory[7854] <=  8'h62;        memory[7855] <=  8'h61;        memory[7856] <=  8'h72;        memory[7857] <=  8'h63;        memory[7858] <=  8'h61;        memory[7859] <=  8'h68;        memory[7860] <=  8'h64;        memory[7861] <=  8'h75;        memory[7862] <=  8'h63;        memory[7863] <=  8'h74;        memory[7864] <=  8'h61;        memory[7865] <=  8'h64;        memory[7866] <=  8'h61;        memory[7867] <=  8'h61;        memory[7868] <=  8'h63;        memory[7869] <=  8'h61;        memory[7870] <=  8'h72;        memory[7871] <=  8'h62;        memory[7872] <=  8'h61;        memory[7873] <=  8'h72;        memory[7874] <=  8'h74;        memory[7875] <=  8'h78;        memory[7876] <=  8'h61;        memory[7877] <=  8'h74;        memory[7878] <=  8'h6b;        memory[7879] <=  8'h73;        memory[7880] <=  8'h68;        memory[7881] <=  8'h63;        memory[7882] <=  8'h66;        memory[7883] <=  8'h69;        memory[7884] <=  8'h77;        memory[7885] <=  8'h68;        memory[7886] <=  8'h61;        memory[7887] <=  8'h74;        memory[7888] <=  8'h61;        memory[7889] <=  8'h6e;        memory[7890] <=  8'h61;        memory[7891] <=  8'h62;        memory[7892] <=  8'h61;        memory[7893] <=  8'h63;        memory[7894] <=  8'h61;        memory[7895] <=  8'h74;        memory[7896] <=  8'h61;        memory[7897] <=  8'h62;        memory[7898] <=  8'h61;        memory[7899] <=  8'h72;        memory[7900] <=  8'h63;        memory[7901] <=  8'h61;        memory[7902] <=  8'h68;        memory[7903] <=  8'h64;        memory[7904] <=  8'h75;        memory[7905] <=  8'h63;        memory[7906] <=  8'h74;        memory[7907] <=  8'h61;        memory[7908] <=  8'h64;        memory[7909] <=  8'h61;        memory[7910] <=  8'h61;        memory[7911] <=  8'h63;        memory[7912] <=  8'h61;        memory[7913] <=  8'h72;        memory[7914] <=  8'h62;        memory[7915] <=  8'h61;        memory[7916] <=  8'h72;        memory[7917] <=  8'h74;        memory[7918] <=  8'h78;        memory[7919] <=  8'h61;        memory[7920] <=  8'h74;        memory[7921] <=  8'h6b;        memory[7922] <=  8'h73;        memory[7923] <=  8'h68;        memory[7924] <=  8'h63;        memory[7925] <=  8'h66;        memory[7926] <=  8'h69;        memory[7927] <=  8'h77;        memory[7928] <=  8'h68;        memory[7929] <=  8'h61;        memory[7930] <=  8'h74;        memory[7931] <=  8'h61;        memory[7932] <=  8'h6e;        memory[7933] <=  8'h61;        memory[7934] <=  8'h62;        memory[7935] <=  8'h61;        memory[7936] <=  8'h63;        memory[7937] <=  8'h61;        memory[7938] <=  8'h74;        memory[7939] <=  8'h61;        memory[7940] <=  8'h62;        memory[7941] <=  8'h61;        memory[7942] <=  8'h72;        memory[7943] <=  8'h63;        memory[7944] <=  8'h61;        memory[7945] <=  8'h68;        memory[7946] <=  8'h64;        memory[7947] <=  8'h75;        memory[7948] <=  8'h63;        memory[7949] <=  8'h74;        memory[7950] <=  8'h61;        memory[7951] <=  8'h64;        memory[7952] <=  8'h61;        memory[7953] <=  8'h61;        memory[7954] <=  8'h63;        memory[7955] <=  8'h61;        memory[7956] <=  8'h72;        memory[7957] <=  8'h62;        memory[7958] <=  8'h61;        memory[7959] <=  8'h72;        memory[7960] <=  8'h74;        memory[7961] <=  8'h74;        memory[7962] <=  8'h62;        memory[7963] <=  8'h61;        memory[7964] <=  8'h72;        memory[7965] <=  8'h74;        memory[7966] <=  8'h78;        memory[7967] <=  8'h61;        memory[7968] <=  8'h74;        memory[7969] <=  8'h6b;        memory[7970] <=  8'h73;        memory[7971] <=  8'h68;        memory[7972] <=  8'h63;        memory[7973] <=  8'h66;        memory[7974] <=  8'h69;        memory[7975] <=  8'h77;        memory[7976] <=  8'h68;        memory[7977] <=  8'h61;        memory[7978] <=  8'h74;        memory[7979] <=  8'h61;        memory[7980] <=  8'h6e;        memory[7981] <=  8'h61;        memory[7982] <=  8'h62;        memory[7983] <=  8'h61;        memory[7984] <=  8'h63;        memory[7985] <=  8'h61;        memory[7986] <=  8'h74;        memory[7987] <=  8'h61;        memory[7988] <=  8'h62;        memory[7989] <=  8'h61;        memory[7990] <=  8'h72;        memory[7991] <=  8'h63;        memory[7992] <=  8'h61;        memory[7993] <=  8'h68;        memory[7994] <=  8'h64;        memory[7995] <=  8'h75;        memory[7996] <=  8'h63;        memory[7997] <=  8'h74;        memory[7998] <=  8'h61;        memory[7999] <=  8'h64;        memory[8000] <=  8'h61;        memory[8001] <=  8'h61;        memory[8002] <=  8'h63;        memory[8003] <=  8'h61;        memory[8004] <=  8'h72;        memory[8005] <=  8'h63;        memory[8006] <=  8'h74;        memory[8007] <=  8'h72;        memory[8008] <=  8'h63;        memory[8009] <=  8'h61;        memory[8010] <=  8'h74;        memory[8011] <=  8'h72;        memory[8012] <=  8'h63;        memory[8013] <=  8'h61;        memory[8014] <=  8'h74;        memory[8015] <=  8'h63;        memory[8016] <=  8'h62;        memory[8017] <=  8'h61;        memory[8018] <=  8'h74;        memory[8019] <=  8'h62;        memory[8020] <=  8'h72;        memory[8021] <=  8'h63;        memory[8022] <=  8'h61;        memory[8023] <=  8'h72;        memory[8024] <=  8'h62;        memory[8025] <=  8'h78;        memory[8026] <=  8'h74;        memory[8027] <=  8'h61;        memory[8028] <=  8'h72;        memory[8029] <=  8'h64;        memory[8030] <=  8'h66;        memory[8031] <=  8'h73;        memory[8032] <=  8'h67;        memory[8033] <=  8'h76;        memory[8034] <=  8'h68;        memory[8035] <=  8'h62;        memory[8036] <=  8'h6b;        memory[8037] <=  8'h6a;        memory[8038] <=  8'h6e;        memory[8039] <=  8'h6d;        memory[8040] <=  8'h62;        memory[8041] <=  8'h76;        memory[8042] <=  8'h78;        memory[8043] <=  8'h63;        memory[8044] <=  8'h73;        memory[8045] <=  8'h66;        memory[8046] <=  8'h72;        memory[8047] <=  8'h74;        memory[8048] <=  8'h79;        memory[8049] <=  8'h75;        memory[8050] <=  8'h6a;        memory[8051] <=  8'h6e;        memory[8052] <=  8'h62;        memory[8053] <=  8'h76;        memory[8054] <=  8'h63;        memory[8055] <=  8'h64;        memory[8056] <=  8'h74;        memory[8057] <=  8'h79;        memory[8058] <=  8'h75;        memory[8059] <=  8'h69;        memory[8060] <=  8'h6b;        memory[8061] <=  8'h6d;        memory[8062] <=  8'h6e;        memory[8063] <=  8'h62;        memory[8064] <=  8'h76;        memory[8065] <=  8'h63;        memory[8066] <=  8'h78;        memory[8067] <=  8'h73;        memory[8068] <=  8'h64;        memory[8069] <=  8'h72;        memory[8070] <=  8'h74;        memory[8071] <=  8'h79;        memory[8072] <=  8'h75;        memory[8073] <=  8'h69;        memory[8074] <=  8'h6b;        memory[8075] <=  8'h6d;        memory[8076] <=  8'h6e;        memory[8077] <=  8'h62;        memory[8078] <=  8'h76;        memory[8079] <=  8'h63;        memory[8080] <=  8'h73;        memory[8081] <=  8'h77;        memory[8082] <=  8'h33;        memory[8083] <=  8'h34;        memory[8084] <=  8'h35;        memory[8085] <=  8'h36;        memory[8086] <=  8'h37;        memory[8087] <=  8'h38;        memory[8088] <=  8'h69;        memory[8089] <=  8'h6b;        memory[8090] <=  8'h6d;        memory[8091] <=  8'h6e;        memory[8092] <=  8'h62;        memory[8093] <=  8'h76;        memory[8094] <=  8'h63;        memory[8095] <=  8'h64;        memory[8096] <=  8'h65;        memory[8097] <=  8'h72;        memory[8098] <=  8'h36;        memory[8099] <=  8'h37;        memory[8100] <=  8'h38;        memory[8101] <=  8'h69;        memory[8102] <=  8'h6f;        memory[8103] <=  8'h6b;        memory[8104] <=  8'h6a;        memory[8105] <=  8'h6e;        memory[8106] <=  8'h62;        memory[8107] <=  8'h76;        memory[8108] <=  8'h63;        memory[8109] <=  8'h64;        memory[8110] <=  8'h72;        memory[8111] <=  8'h74;        memory[8112] <=  8'h79;        memory[8113] <=  8'h75;        memory[8114] <=  8'h73;        memory[8115] <=  8'h6a;        memory[8116] <=  8'h63;        memory[8117] <=  8'h6e;        memory[8118] <=  8'h62;        memory[8119] <=  8'h64;        memory[8120] <=  8'h66;        memory[8121] <=  8'h73;        memory[8122] <=  8'h74;        memory[8123] <=  8'h79;        memory[8124] <=  8'h75;        memory[8125] <=  8'h61;        memory[8126] <=  8'h69;        memory[8127] <=  8'h6b;        memory[8128] <=  8'h78;        memory[8129] <=  8'h6d;        memory[8130] <=  8'h6e;        memory[8131] <=  8'h73;        memory[8132] <=  8'h6a;        memory[8133] <=  8'h6f;        memory[8134] <=  8'h64;        memory[8135] <=  8'h6c;        memory[8136] <=  8'h63;        memory[8137] <=  8'h78;        memory[8138] <=  8'h2c;        memory[8139] <=  8'h6d;        memory[8140] <=  8'h73;        memory[8141] <=  8'h6b;        memory[8142] <=  8'h64;        memory[8143] <=  8'h6c;        memory[8144] <=  8'h70;        memory[8145] <=  8'h5b;        memory[8146] <=  8'h3b;        memory[8147] <=  8'h73;        memory[8148] <=  8'h6c;        memory[8149] <=  8'h64;        memory[8150] <=  8'h70;        memory[8151] <=  8'h76;        memory[8152] <=  8'h63;        memory[8153] <=  8'h5b;        memory[8154] <=  8'h78;        memory[8155] <=  8'h76;        memory[8156] <=  8'h63;        memory[8157] <=  8'h5b;        memory[8158] <=  8'h78;        memory[8159] <=  8'h70;        memory[8160] <=  8'h6f;        memory[8161] <=  8'h20;        memory[8162] <=  8'h62;        memory[8163] <=  8'h61;        memory[8164] <=  8'h72;        memory[8165] <=  8'h74;        memory[8166] <=  8'h74;        memory[8167] <=  8'h62;        memory[8168] <=  8'h61;        memory[8169] <=  8'h72;        memory[8170] <=  8'h74;        memory[8171] <=  8'h78;        memory[8172] <=  8'h61;        memory[8173] <=  8'h74;        memory[8174] <=  8'h6b;        memory[8175] <=  8'h73;        memory[8176] <=  8'h68;        memory[8177] <=  8'h63;        memory[8178] <=  8'h66;        memory[8179] <=  8'h69;        memory[8180] <=  8'h77;        memory[8181] <=  8'h68;        memory[8182] <=  8'h61;        memory[8183] <=  8'h69;        memory[8184] <=  8'h6a;        memory[8185] <=  8'h78;        memory[8186] <=  8'h5d;        memory[8187] <=  8'h65;        memory[8188] <=  8'h6b;        memory[8189] <=  8'h6f;        memory[8190] <=  8'h39;        memory[8191] <=  8'h64;        memory[8192] <=  8'h75;        memory[8193] <=  8'h38;        memory[8194] <=  8'h79;        memory[8195] <=  8'h20;        memory[8196] <=  8'h37;        memory[8197] <=  8'h63;        memory[8198] <=  8'h67;        memory[8199] <=  8'h78;        memory[8200] <=  8'h63;        memory[8201] <=  8'h75;        memory[8202] <=  8'h68;        memory[8203] <=  8'h69;        memory[8204] <=  8'h6a;        memory[8205] <=  8'h77;        memory[8206] <=  8'h69;        memory[8207] <=  8'h64;        memory[8208] <=  8'h66;        memory[8209] <=  8'h68;        memory[8210] <=  8'h75;        memory[8211] <=  8'h76;        memory[8212] <=  8'h64;        memory[8213] <=  8'h62;        memory[8214] <=  8'h66;        memory[8215] <=  8'h6a;        memory[8216] <=  8'h6e;        memory[8217] <=  8'h6b;        memory[8218] <=  8'h6a;        memory[8219] <=  8'h65;        memory[8220] <=  8'h38;        memory[8221] <=  8'h66;        memory[8222] <=  8'h37;        memory[8223] <=  8'h67;        memory[8224] <=  8'h79;        memory[8225] <=  8'h76;        memory[8226] <=  8'h63;        memory[8227] <=  8'h68;        memory[8228] <=  8'h69;        memory[8229] <=  8'h6a;        memory[8230] <=  8'h33;        memory[8231] <=  8'h65;        memory[8232] <=  8'h67;        memory[8233] <=  8'h79;        memory[8234] <=  8'h72;        memory[8235] <=  8'h64;        memory[8236] <=  8'h62;        memory[8237] <=  8'h6e;        memory[8238] <=  8'h63;        memory[8239] <=  8'h7a;        memory[8240] <=  8'h6a;        memory[8241] <=  8'h6f;        memory[8242] <=  8'h66;        memory[8243] <=  8'h78;        memory[8244] <=  8'h6a;        memory[8245] <=  8'h69;        memory[8246] <=  8'h63;        memory[8247] <=  8'h68;        memory[8248] <=  8'h62;        memory[8249] <=  8'h6e;        memory[8250] <=  8'h6d;        memory[8251] <=  8'h63;        memory[8252] <=  8'h73;        memory[8253] <=  8'h6c;        memory[8254] <=  8'h6b;        memory[8255] <=  8'h6a;        memory[8256] <=  8'h69;        memory[8257] <=  8'h68;        memory[8258] <=  8'h76;        memory[8259] <=  8'h75;        memory[8260] <=  8'h69;        memory[8261] <=  8'h64;        memory[8262] <=  8'h68;        memory[8263] <=  8'h75;        memory[8264] <=  8'h67;        memory[8265] <=  8'h79;        memory[8266] <=  8'h62;        memory[8267] <=  8'h68;        memory[8268] <=  8'h65;        memory[8269] <=  8'h6a;        memory[8270] <=  8'h72;        memory[8271] <=  8'h6b;        memory[8272] <=  8'h6a;        memory[8273] <=  8'h6f;        memory[8274] <=  8'h64;        memory[8275] <=  8'h67;        memory[8276] <=  8'h69;        memory[8277] <=  8'h75;        memory[8278] <=  8'h69;        memory[8279] <=  8'h67;        memory[8280] <=  8'h76;        memory[8281] <=  8'h79;        memory[8282] <=  8'h75;        memory[8283] <=  8'h67;        memory[8284] <=  8'h78;        memory[8285] <=  8'h68;        memory[8286] <=  8'h63;        memory[8287] <=  8'h20;        memory[8288] <=  8'h20;        memory[8289] <=  8'h20;        memory[8290] <=  8'h78;        memory[8291] <=  8'h76;        memory[8292] <=  8'h20;        memory[8293] <=  8'h63;        memory[8294] <=  8'h78;        memory[8295] <=  8'h67;        memory[8296] <=  8'h79;        memory[8297] <=  8'h63;        memory[8298] <=  8'h75;        memory[8299] <=  8'h68;        memory[8300] <=  8'h6a;        memory[8301] <=  8'h6b;        memory[8302] <=  8'h61;        memory[8303] <=  8'h6c;        memory[8304] <=  8'h78;        memory[8305] <=  8'h76;        memory[8306] <=  8'h70;        memory[8307] <=  8'h6f;        memory[8308] <=  8'h69;        memory[8309] <=  8'h6a;        memory[8310] <=  8'h69;        memory[8311] <=  8'h68;        memory[8312] <=  8'h6a;        memory[8313] <=  8'h62;        memory[8314] <=  8'h77;        memory[8315] <=  8'h65;        memory[8316] <=  8'h6e;        memory[8317] <=  8'h61;        memory[8318] <=  8'h66;        memory[8319] <=  8'h6d;        memory[8320] <=  8'h64;        memory[8321] <=  8'h6b;        memory[8322] <=  8'h6d;        memory[8323] <=  8'h76;        memory[8324] <=  8'h6c;        memory[8325] <=  8'h63;        memory[8326] <=  8'h6f;        memory[8327] <=  8'h64;        memory[8328] <=  8'h69;        memory[8329] <=  8'h75;        memory[8330] <=  8'h68;        memory[8331] <=  8'h73;        memory[8332] <=  8'h66;        memory[8333] <=  8'h65;        memory[8334] <=  8'h62;        memory[8335] <=  8'h6e;        memory[8336] <=  8'h64;        memory[8337] <=  8'h73;        memory[8338] <=  8'h63;        memory[8339] <=  8'h6b;        memory[8340] <=  8'h20;        memory[8341] <=  8'h78;        memory[8342] <=  8'h6a;        memory[8343] <=  8'h78;        memory[8344] <=  8'h63;        memory[8345] <=  8'h73;        memory[8346] <=  8'h64;        memory[8347] <=  8'h66;        memory[8348] <=  8'h6b;        memory[8349] <=  8'h64;        memory[8350] <=  8'h6e;        memory[8351] <=  8'h6d;        memory[8352] <=  8'h64;        memory[8353] <=  8'h73;        memory[8354] <=  8'h63;        memory[8355] <=  8'h6b;        memory[8356] <=  8'h78;        memory[8357] <=  8'h6c;        memory[8358] <=  8'h6f;        memory[8359] <=  8'h66;        memory[8360] <=  8'h6a;        memory[8361] <=  8'h69;        memory[8362] <=  8'h61;        memory[8363] <=  8'h62;        memory[8364] <=  8'h6e;        memory[8365] <=  8'h20;        memory[8366] <=  8'h78;        memory[8367] <=  8'h6b;        memory[8368] <=  8'h6d;        memory[8369] <=  8'h20;        memory[8370] <=  8'h6f;        memory[8371] <=  8'h63;        memory[8372] <=  8'h76;        memory[8373] <=  8'h73;        memory[8374] <=  8'h64;        memory[8375] <=  8'h69;        memory[8376] <=  8'h66;        memory[8377] <=  8'h68;        memory[8378] <=  8'h65;        memory[8379] <=  8'h71;        memory[8380] <=  8'h6a;        memory[8381] <=  8'h77;        memory[8382] <=  8'h62;        memory[8383] <=  8'h65;        memory[8384] <=  8'h6e;        memory[8385] <=  8'h20;        memory[8386] <=  8'h6d;        memory[8387] <=  8'h64;        memory[8388] <=  8'h73;        memory[8389] <=  8'h6c;        memory[8390] <=  8'h76;        memory[8391] <=  8'h6b;        memory[8392] <=  8'h63;        memory[8393] <=  8'h78;        memory[8394] <=  8'h20;        memory[8395] <=  8'h6f;        memory[8396] <=  8'h78;        memory[8397] <=  8'h69;        memory[8398] <=  8'h63;        memory[8399] <=  8'h6a;        memory[8400] <=  8'h76;        memory[8401] <=  8'h64;        memory[8402] <=  8'h66;        memory[8403] <=  8'h65;        memory[8404] <=  8'h71;        memory[8405] <=  8'h6e;        memory[8406] <=  8'h20;        memory[8407] <=  8'h64;        memory[8408] <=  8'h6d;        memory[8409] <=  8'h73;        memory[8410] <=  8'h6c;        memory[8411] <=  8'h63;        memory[8412] <=  8'h78;        memory[8413] <=  8'h6b;        memory[8414] <=  8'h20;        memory[8415] <=  8'h6f;        memory[8416] <=  8'h78;        memory[8417] <=  8'h63;        memory[8418] <=  8'h76;        memory[8419] <=  8'h6a;        memory[8420] <=  8'h64;        memory[8421] <=  8'h62;        memory[8422] <=  8'h71;        memory[8423] <=  8'h77;        memory[8424] <=  8'h65;        memory[8425] <=  8'h6e;        memory[8426] <=  8'h6d;        memory[8427] <=  8'h64;        memory[8428] <=  8'h6c;        memory[8429] <=  8'h73;        memory[8430] <=  8'h2c;        memory[8431] <=  8'h76;        memory[8432] <=  8'h63;        memory[8433] <=  8'h78;        memory[8434] <=  8'h20;        memory[8435] <=  8'h63;        memory[8436] <=  8'h6f;        memory[8437] <=  8'h69;        memory[8438] <=  8'h76;        memory[8439] <=  8'h68;        memory[8440] <=  8'h73;        memory[8441] <=  8'h64;        memory[8442] <=  8'h62;        memory[8443] <=  8'h71;        memory[8444] <=  8'h77;        memory[8445] <=  8'h65;        memory[8446] <=  8'h6e;        memory[8447] <=  8'h64;        memory[8448] <=  8'h6b;        memory[8449] <=  8'h73;        memory[8450] <=  8'h76;        memory[8451] <=  8'h6f;        memory[8452] <=  8'h63;        memory[8453] <=  8'h20;        memory[8454] <=  8'h76;        memory[8455] <=  8'h69;        memory[8456] <=  8'h75;        memory[8457] <=  8'h69;        memory[8458] <=  8'h68;        memory[8459] <=  8'h63;        memory[8460] <=  8'h78;        memory[8461] <=  8'h69;        memory[8462] <=  8'h6f;        memory[8463] <=  8'h76;        memory[8464] <=  8'h73;        memory[8465] <=  8'h64;        memory[8466] <=  8'h61;        memory[8467] <=  8'h64;        memory[8468] <=  8'h6e;        memory[8469] <=  8'h77;        memory[8470] <=  8'h71;        memory[8471] <=  8'h6b;        memory[8472] <=  8'h6c;        memory[8473] <=  8'h73;        memory[8474] <=  8'h76;        memory[8475] <=  8'h6e;        memory[8476] <=  8'h62;        memory[8477] <=  8'h20;        memory[8478] <=  8'h64;        memory[8479] <=  8'h66;        memory[8480] <=  8'h6a;        memory[8481] <=  8'h6b;        memory[8482] <=  8'h71;        memory[8483] <=  8'h64;        memory[8484] <=  8'h77;        memory[8485] <=  8'h65;        memory[8486] <=  8'h6e;        memory[8487] <=  8'h62;        memory[8488] <=  8'h20;        memory[8489] <=  8'h64;        memory[8490] <=  8'h73;        memory[8491] <=  8'h76;        memory[8492] <=  8'h68;        memory[8493] <=  8'h64;        memory[8494] <=  8'h61;        memory[8495] <=  8'h71;        memory[8496] <=  8'h77;        memory[8497] <=  8'h6a;        memory[8498] <=  8'h65;        memory[8499] <=  8'h6e;        memory[8500] <=  8'h64;        memory[8501] <=  8'h20;        memory[8502] <=  8'h61;        memory[8503] <=  8'h63;        memory[8504] <=  8'h62;        memory[8505] <=  8'h68;        memory[8506] <=  8'h64;        memory[8507] <=  8'h61;        memory[8508] <=  8'h77;        memory[8509] <=  8'h71;        memory[8510] <=  8'h6e;        memory[8511] <=  8'h20;        memory[8512] <=  8'h62;        memory[8513] <=  8'h73;        memory[8514] <=  8'h76;        memory[8515] <=  8'h61;        memory[8516] <=  8'h67;        memory[8517] <=  8'h76;        memory[8518] <=  8'h68;        memory[8519] <=  8'h67;        memory[8520] <=  8'h61;        memory[8521] <=  8'h73;        memory[8522] <=  8'h6a;        memory[8523] <=  8'h6b;        memory[8524] <=  8'h63;        memory[8525] <=  8'h78;        memory[8526] <=  8'h76;        memory[8527] <=  8'h6e;        memory[8528] <=  8'h73;        memory[8529] <=  8'h64;        memory[8530] <=  8'h20;        memory[8531] <=  8'h66;        memory[8532] <=  8'h62;        memory[8533] <=  8'h64;        memory[8534] <=  8'h61;        memory[8535] <=  8'h73;        memory[8536] <=  8'h76;        memory[8537] <=  8'h67;        memory[8538] <=  8'h63;        memory[8539] <=  8'h79;        memory[8540] <=  8'h7a;        memory[8541] <=  8'h78;        memory[8542] <=  8'h79;        memory[8543] <=  8'h75;        memory[8544] <=  8'h20;        memory[8545] <=  8'h69;        memory[8546] <=  8'h6a;        memory[8547] <=  8'h64;        memory[8548] <=  8'h66;        memory[8549] <=  8'h6b;        memory[8550] <=  8'h61;        memory[8551] <=  8'h64;        memory[8552] <=  8'h63;        memory[8553] <=  8'h78;        memory[8554] <=  8'h68;        memory[8555] <=  8'h20;        memory[8556] <=  8'h67;        memory[8557] <=  8'h61;        memory[8558] <=  8'h68;        memory[8559] <=  8'h75;        memory[8560] <=  8'h64;        memory[8561] <=  8'h73;        memory[8562] <=  8'h69;        memory[8563] <=  8'h6a;        memory[8564] <=  8'h61;        memory[8565] <=  8'h6b;        memory[8566] <=  8'h63;        memory[8567] <=  8'h62;        memory[8568] <=  8'h61;        memory[8569] <=  8'h72;        memory[8570] <=  8'h73;        memory[8571] <=  8'h68;        memory[8572] <=  8'h64;        memory[8573] <=  8'h66;        memory[8574] <=  8'h67;        memory[8575] <=  8'h73;        memory[8576] <=  8'h68;        memory[8577] <=  8'h64;        memory[8578] <=  8'h66;        memory[8579] <=  8'h68;        memory[8580] <=  8'h64;        memory[8581] <=  8'h6a;        memory[8582] <=  8'h68;        memory[8583] <=  8'h62;        memory[8584] <=  8'h67;        memory[8585] <=  8'h63;        memory[8586] <=  8'h61;        memory[8587] <=  8'h66;        memory[8588] <=  8'h73;        memory[8589] <=  8'h79;        memory[8590] <=  8'h67;        memory[8591] <=  8'h6b;        memory[8592] <=  8'h75;        memory[8593] <=  8'h64;        memory[8594] <=  8'h68;        memory[8595] <=  8'h62;        memory[8596] <=  8'h77;        memory[8597] <=  8'h76;        memory[8598] <=  8'h67;        memory[8599] <=  8'h61;        memory[8600] <=  8'h66;        memory[8601] <=  8'h64;        memory[8602] <=  8'h74;        memory[8603] <=  8'h75;        memory[8604] <=  8'h66;        memory[8605] <=  8'h79;        memory[8606] <=  8'h67;        memory[8607] <=  8'h69;        memory[8608] <=  8'h75;        memory[8609] <=  8'h68;        memory[8610] <=  8'h6c;        memory[8611] <=  8'h6a;        memory[8612] <=  8'h62;        memory[8613] <=  8'h6b;        memory[8614] <=  8'h68;        memory[8615] <=  8'h76;        memory[8616] <=  8'h67;        memory[8617] <=  8'h63;        memory[8618] <=  8'h66;        memory[8619] <=  8'h78;        memory[8620] <=  8'h64;        memory[8621] <=  8'h74;        memory[8622] <=  8'h75;        memory[8623] <=  8'h79;        memory[8624] <=  8'h69;        memory[8625] <=  8'h75;        memory[8626] <=  8'h68;        memory[8627] <=  8'h6c;        memory[8628] <=  8'h6a;        memory[8629] <=  8'h6b;        memory[8630] <=  8'h67;        memory[8631] <=  8'h6a;        memory[8632] <=  8'h63;        memory[8633] <=  8'h66;        memory[8634] <=  8'h68;        memory[8635] <=  8'h64;        memory[8636] <=  8'h67;        memory[8637] <=  8'h72;        memory[8638] <=  8'h79;        memory[8639] <=  8'h74;        memory[8640] <=  8'h66;        memory[8641] <=  8'h75;        memory[8642] <=  8'h79;        memory[8643] <=  8'h69;        memory[8644] <=  8'h68;        memory[8645] <=  8'h6c;        memory[8646] <=  8'h62;        memory[8647] <=  8'h6d;        memory[8648] <=  8'h76;        memory[8649] <=  8'h6e;        memory[8650] <=  8'h63;        memory[8651] <=  8'h66;        memory[8652] <=  8'h68;        memory[8653] <=  8'h64;        memory[8654] <=  8'h74;        memory[8655] <=  8'h75;        memory[8656] <=  8'h67;        memory[8657] <=  8'h79;        memory[8658] <=  8'h69;        memory[8659] <=  8'h68;        memory[8660] <=  8'h75;        memory[8661] <=  8'h6a;        memory[8662] <=  8'h6c;        memory[8663] <=  8'h62;        memory[8664] <=  8'h6d;        memory[8665] <=  8'h76;        memory[8666] <=  8'h6e;        memory[8667] <=  8'h63;        memory[8668] <=  8'h66;        memory[8669] <=  8'h68;        memory[8670] <=  8'h67;        memory[8671] <=  8'h79;        memory[8672] <=  8'h68;        memory[8673] <=  8'h75;        memory[8674] <=  8'h6a;        memory[8675] <=  8'h6e;        memory[8676] <=  8'h2c;        memory[8677] <=  8'h62;        memory[8678] <=  8'h6e;        memory[8679] <=  8'h6d;        memory[8680] <=  8'h76;        memory[8681] <=  8'h6e;        memory[8682] <=  8'h63;        memory[8683] <=  8'h66;        memory[8684] <=  8'h68;        memory[8685] <=  8'h74;        memory[8686] <=  8'h79;        memory[8687] <=  8'h69;        memory[8688] <=  8'h75;        memory[8689] <=  8'h6c;        memory[8690] <=  8'h6a;        memory[8691] <=  8'h62;        memory[8692] <=  8'h6d;        memory[8693] <=  8'h76;        memory[8694] <=  8'h6e;        memory[8695] <=  8'h63;        memory[8696] <=  8'h66;        memory[8697] <=  8'h74;        memory[8698] <=  8'h75;        memory[8699] <=  8'h79;        memory[8700] <=  8'h69;        memory[8701] <=  8'h68;        memory[8702] <=  8'h6b;        memory[8703] <=  8'h62;        memory[8704] <=  8'h76;        memory[8705] <=  8'h63;        memory[8706] <=  8'h66;        memory[8707] <=  8'h67;        memory[8708] <=  8'h74;        memory[8709] <=  8'h75;        memory[8710] <=  8'h79;        memory[8711] <=  8'h69;        memory[8712] <=  8'h75;        memory[8713] <=  8'h68;        memory[8714] <=  8'h6a;        memory[8715] <=  8'h6b;        memory[8716] <=  8'h62;        memory[8717] <=  8'h76;        memory[8718] <=  8'h63;        memory[8719] <=  8'h66;        memory[8720] <=  8'h74;        memory[8721] <=  8'h75;        memory[8722] <=  8'h79;        memory[8723] <=  8'h69;        memory[8724] <=  8'h75;        memory[8725] <=  8'h6a;        memory[8726] <=  8'h6b;        memory[8727] <=  8'h6e;        memory[8728] <=  8'h62;        memory[8729] <=  8'h76;        memory[8730] <=  8'h67;        memory[8731] <=  8'h66;        memory[8732] <=  8'h74;        memory[8733] <=  8'h79;        memory[8734] <=  8'h75;        memory[8735] <=  8'h75;        memory[8736] <=  8'h69;        memory[8737] <=  8'h6a;        memory[8738] <=  8'h6b;        memory[8739] <=  8'h68;        memory[8740] <=  8'h62;        memory[8741] <=  8'h6a;        memory[8742] <=  8'h67;        memory[8743] <=  8'h68;        memory[8744] <=  8'h66;        memory[8745] <=  8'h79;        memory[8746] <=  8'h74;        memory[8747] <=  8'h79;        memory[8748] <=  8'h69;        memory[8749] <=  8'h75;        memory[8750] <=  8'h64;        memory[8751] <=  8'h6a;        memory[8752] <=  8'h6b;        memory[8753] <=  8'h68;        memory[8754] <=  8'h63;        memory[8755] <=  8'h7a;        memory[8756] <=  8'h67;        memory[8757] <=  8'h68;        memory[8758] <=  8'h74;        memory[8759] <=  8'h75;        memory[8760] <=  8'h79;        memory[8761] <=  8'h69;        memory[8762] <=  8'h61;        memory[8763] <=  8'h73;        memory[8764] <=  8'h75;        memory[8765] <=  8'h6a;        memory[8766] <=  8'h6b;        memory[8767] <=  8'h62;        memory[8768] <=  8'h6e;        memory[8769] <=  8'h61;        memory[8770] <=  8'h76;        memory[8771] <=  8'h63;        memory[8772] <=  8'h66;        memory[8773] <=  8'h68;        memory[8774] <=  8'h75;        memory[8775] <=  8'h61;        memory[8776] <=  8'h73;        memory[8777] <=  8'h79;        memory[8778] <=  8'h64;        memory[8779] <=  8'h75;        memory[8780] <=  8'h69;        memory[8781] <=  8'h6a;        memory[8782] <=  8'h61;        memory[8783] <=  8'h6b;        memory[8784] <=  8'h62;        memory[8785] <=  8'h63;        memory[8786] <=  8'h78;        memory[8787] <=  8'h68;        memory[8788] <=  8'h67;        memory[8789] <=  8'h79;        memory[8790] <=  8'h75;        memory[8791] <=  8'h7a;        memory[8792] <=  8'h63;        memory[8793] <=  8'h61;        memory[8794] <=  8'h73;        memory[8795] <=  8'h69;        memory[8796] <=  8'h75;        memory[8797] <=  8'h6f;        memory[8798] <=  8'h69;        memory[8799] <=  8'h6a;        memory[8800] <=  8'h61;        memory[8801] <=  8'h6c;        memory[8802] <=  8'h63;        memory[8803] <=  8'h78;        memory[8804] <=  8'h62;        memory[8805] <=  8'h63;        memory[8806] <=  8'h20;        memory[8807] <=  8'h6e;        memory[8808] <=  8'h76;        memory[8809] <=  8'h63;        memory[8810] <=  8'h61;        memory[8811] <=  8'h64;        memory[8812] <=  8'h73;        memory[8813] <=  8'h67;        memory[8814] <=  8'h79;        memory[8815] <=  8'h68;        memory[8816] <=  8'h75;        memory[8817] <=  8'h61;        memory[8818] <=  8'h6a;        memory[8819] <=  8'h6b;        memory[8820] <=  8'h78;        memory[8821] <=  8'h62;        memory[8822] <=  8'h20;        memory[8823] <=  8'h6e;        memory[8824] <=  8'h76;        memory[8825] <=  8'h63;        memory[8826] <=  8'h61;        memory[8827] <=  8'h73;        memory[8828] <=  8'h67;        memory[8829] <=  8'h68;        memory[8830] <=  8'h75;        memory[8831] <=  8'h6a;        memory[8832] <=  8'h6c;        memory[8833] <=  8'h6b;        memory[8834] <=  8'h63;        memory[8835] <=  8'h78;        memory[8836] <=  8'h20;        memory[8837] <=  8'h6a;        memory[8838] <=  8'h6b;        memory[8839] <=  8'h68;        memory[8840] <=  8'h61;        memory[8841] <=  8'h73;        memory[8842] <=  8'h76;        memory[8843] <=  8'h64;        memory[8844] <=  8'h6e;        memory[8845] <=  8'h20;        memory[8846] <=  8'h62;        memory[8847] <=  8'h6e;        memory[8848] <=  8'h6d;        memory[8849] <=  8'h6b;        memory[8850] <=  8'h77;        memory[8851] <=  8'h64;        memory[8852] <=  8'h6f;        memory[8853] <=  8'h77;        memory[8854] <=  8'h69;        memory[8855] <=  8'h6f;        memory[8856] <=  8'h75;        memory[8857] <=  8'h69;        memory[8858] <=  8'h68;        memory[8859] <=  8'h62;        memory[8860] <=  8'h6e;        memory[8861] <=  8'h6b;        memory[8862] <=  8'h77;        memory[8863] <=  8'h69;        memory[8864] <=  8'h6f;        memory[8865] <=  8'h75;        memory[8866] <=  8'h71;        memory[8867] <=  8'h69;        memory[8868] <=  8'h79;        memory[8869] <=  8'h67;        memory[8870] <=  8'h6a;        memory[8871] <=  8'h64;        memory[8872] <=  8'h61;        memory[8873] <=  8'h76;        memory[8874] <=  8'h62;        memory[8875] <=  8'h6e;        memory[8876] <=  8'h6b;        memory[8877] <=  8'h6f;        memory[8878] <=  8'h70;        memory[8879] <=  8'h64;        memory[8880] <=  8'h76;        memory[8881] <=  8'h69;        memory[8882] <=  8'h6f;        memory[8883] <=  8'h75;        memory[8884] <=  8'h69;        memory[8885] <=  8'h48;        memory[8886] <=  8'h42;        memory[8887] <=  8'h6b;        memory[8888] <=  8'h64;        memory[8889] <=  8'h6e;        memory[8890] <=  8'h6c;        memory[8891] <=  8'h71;        memory[8892] <=  8'h6b;        memory[8893] <=  8'h6d;        memory[8894] <=  8'h6a;        memory[8895] <=  8'h70;        memory[8896] <=  8'h69;        memory[8897] <=  8'h6f;        memory[8898] <=  8'h68;        memory[8899] <=  8'h65;        memory[8900] <=  8'h66;        memory[8901] <=  8'h75;        memory[8902] <=  8'h67;        memory[8903] <=  8'h69;        memory[8904] <=  8'h73;        memory[8905] <=  8'h61;        memory[8906] <=  8'h62;        memory[8907] <=  8'h64;        memory[8908] <=  8'h6b;        memory[8909] <=  8'h6a;        memory[8910] <=  8'h6b;        memory[8911] <=  8'h6c;        memory[8912] <=  8'h6a;        memory[8913] <=  8'h69;        memory[8914] <=  8'h73;        memory[8915] <=  8'h6f;        memory[8916] <=  8'h71;        memory[8917] <=  8'h68;        memory[8918] <=  8'h77;        memory[8919] <=  8'h67;        memory[8920] <=  8'h69;        memory[8921] <=  8'h79;        memory[8922] <=  8'h6a;        memory[8923] <=  8'h64;        memory[8924] <=  8'h76;        memory[8925] <=  8'h62;        memory[8926] <=  8'h6e;        memory[8927] <=  8'h61;        memory[8928] <=  8'h73;        memory[8929] <=  8'h66;        memory[8930] <=  8'h6c;        memory[8931] <=  8'h6b;        memory[8932] <=  8'h64;        memory[8933] <=  8'h6a;        memory[8934] <=  8'h68;        memory[8935] <=  8'h63;        memory[8936] <=  8'h67;        memory[8937] <=  8'h6a;        memory[8938] <=  8'h76;        memory[8939] <=  8'h73;        memory[8940] <=  8'h64;        memory[8941] <=  8'h62;        memory[8942] <=  8'h62;        memory[8943] <=  8'h61;        memory[8944] <=  8'h72;        memory[8945] <=  8'h62;        memory[8946] <=  8'h62;        memory[8947] <=  8'h73;        memory[8948] <=  8'h62;        memory[8949] <=  8'h67;        memory[8950] <=  8'h73;        memory[8951] <=  8'h66;        memory[8952] <=  8'h67;        memory[8953] <=  8'h61;        memory[8954] <=  8'h68;        memory[8955] <=  8'h66;        memory[8956] <=  8'h73;        memory[8957] <=  8'h68;        memory[8958] <=  8'h61;        memory[8959] <=  8'h66;        memory[8960] <=  8'h73;        memory[8961] <=  8'h66;        memory[8962] <=  8'h68;        memory[8963] <=  8'h61;        memory[8964] <=  8'h69;        memory[8965] <=  8'h64;        memory[8966] <=  8'h75;        memory[8967] <=  8'h67;        memory[8968] <=  8'h64;        memory[8969] <=  8'h77;        memory[8970] <=  8'h62;        memory[8971] <=  8'h61;        memory[8972] <=  8'h62;        memory[8973] <=  8'h72;        memory[8974] <=  8'h62;        memory[8975] <=  8'h61;        memory[8976] <=  8'h62;        memory[8977] <=  8'h62;        memory[8978] <=  8'h74;        memory[8979] <=  8'h62;        memory[8980] <=  8'h62;        memory[8981] <=  8'h62;        memory[8982] <=  8'h62;        memory[8983] <=  8'h62;        memory[8984] <=  8'h62;        memory[8985] <=  8'h62;        memory[8986] <=  8'h62;        memory[8987] <=  8'h61;        memory[8988] <=  8'h62;        memory[8989] <=  8'h62;        memory[8990] <=  8'h72;        memory[8991] <=  8'h74;        memory[8992] <=  8'h62;        memory[8993] <=  8'h62;        memory[8994] <=  8'h61;        memory[8995] <=  8'h62;        memory[8996] <=  8'h72;        memory[8997] <=  8'h62;        memory[8998] <=  8'h74;        memory[8999] <=  8'h62;        memory[9000] <=  8'h62;        memory[9001] <=  8'h62;        memory[9002] <=  8'h63;        memory[9003] <=  8'h61;        memory[9004] <=  8'h72;        memory[9005] <=  8'h74;        memory[9006] <=  8'h73;        memory[9007] <=  8'h62;        memory[9008] <=  8'h61;        memory[9009] <=  8'h72;        memory[9010] <=  8'h74;        memory[9011] <=  8'h74;        memory[9012] <=  8'h62;        memory[9013] <=  8'h61;        memory[9014] <=  8'h72;        memory[9015] <=  8'h74;        memory[9016] <=  8'h78;        memory[9017] <=  8'h61;        memory[9018] <=  8'h74;        memory[9019] <=  8'h6b;        memory[9020] <=  8'h73;        memory[9021] <=  8'h68;        memory[9022] <=  8'h63;        memory[9023] <=  8'h66;        memory[9024] <=  8'h69;        memory[9025] <=  8'h77;        memory[9026] <=  8'h68;        memory[9027] <=  8'h61;        memory[9028] <=  8'h74;        memory[9029] <=  8'h61;        memory[9030] <=  8'h6e;        memory[9031] <=  8'h61;        memory[9032] <=  8'h62;        memory[9033] <=  8'h61;        memory[9034] <=  8'h63;        memory[9035] <=  8'h61;        memory[9036] <=  8'h74;        memory[9037] <=  8'h61;        memory[9038] <=  8'h62;        memory[9039] <=  8'h61;        memory[9040] <=  8'h72;        memory[9041] <=  8'h63;        memory[9042] <=  8'h61;        memory[9043] <=  8'h68;        memory[9044] <=  8'h64;        memory[9045] <=  8'h75;        memory[9046] <=  8'h63;        memory[9047] <=  8'h74;        memory[9048] <=  8'h61;        memory[9049] <=  8'h64;        memory[9050] <=  8'h61;        memory[9051] <=  8'h61;        memory[9052] <=  8'h63;        memory[9053] <=  8'h61;        memory[9054] <=  8'h72;        memory[9055] <=  8'h63;        memory[9056] <=  8'h74;        memory[9057] <=  8'h72;        memory[9058] <=  8'h63;        memory[9059] <=  8'h61;        memory[9060] <=  8'h74;        memory[9061] <=  8'h72;        memory[9062] <=  8'h63;        memory[9063] <=  8'h61;        memory[9064] <=  8'h74;        memory[9065] <=  8'h63;        memory[9066] <=  8'h62;        memory[9067] <=  8'h61;        memory[9068] <=  8'h74;        memory[9069] <=  8'h62;        memory[9070] <=  8'h72;        memory[9071] <=  8'h63;        memory[9072] <=  8'h61;        memory[9073] <=  8'h74;        memory[9074] <=  8'h72;        memory[9075] <=  8'h6e;        memory[9076] <=  8'h62;        memory[9077] <=  8'h61;        memory[9078] <=  8'h63;        memory[9079] <=  8'h61;        memory[9080] <=  8'h74;        memory[9081] <=  8'h79;        memory[9082] <=  8'h73;        memory[9083] <=  8'h6e;        memory[9084] <=  8'h63;        memory[9085] <=  8'h74;        memory[9086] <=  8'h61;        memory[9087] <=  8'h6e;        memory[9088] <=  8'h62;        memory[9089] <=  8'h61;        memory[9090] <=  8'h63;        memory[9091] <=  8'h72;        memory[9092] <=  8'h6e;        memory[9093] <=  8'h74;        memory[9094] <=  8'h61;        memory[9095] <=  8'h62;        memory[9096] <=  8'h74;        memory[9097] <=  8'h6e;        memory[9098] <=  8'h61;        memory[9099] <=  8'h72;        memory[9100] <=  8'h62;        memory[9101] <=  8'h78;        memory[9102] <=  8'h74;        memory[9103] <=  8'h61;        memory[9104] <=  8'h72;        memory[9105] <=  8'h62;        memory[9106] <=  8'h61;        memory[9107] <=  8'h72;        memory[9108] <=  8'h74;        memory[9109] <=  8'h74;        memory[9110] <=  8'h62;        memory[9111] <=  8'h61;        memory[9112] <=  8'h72;        memory[9113] <=  8'h74;        memory[9114] <=  8'h78;        memory[9115] <=  8'h61;        memory[9116] <=  8'h74;        memory[9117] <=  8'h6b;        memory[9118] <=  8'h73;        memory[9119] <=  8'h68;        memory[9120] <=  8'h63;        memory[9121] <=  8'h66;        memory[9122] <=  8'h69;        memory[9123] <=  8'h77;        memory[9124] <=  8'h68;        memory[9125] <=  8'h61;        memory[9126] <=  8'h74;        memory[9127] <=  8'h61;        memory[9128] <=  8'h6e;        memory[9129] <=  8'h61;        memory[9130] <=  8'h62;        memory[9131] <=  8'h61;        memory[9132] <=  8'h63;        memory[9133] <=  8'h61;        memory[9134] <=  8'h74;        memory[9135] <=  8'h61;        memory[9136] <=  8'h62;        memory[9137] <=  8'h61;        memory[9138] <=  8'h72;        memory[9139] <=  8'h63;        memory[9140] <=  8'h61;        memory[9141] <=  8'h68;        memory[9142] <=  8'h64;        memory[9143] <=  8'h75;        memory[9144] <=  8'h63;        memory[9145] <=  8'h74;        memory[9146] <=  8'h61;        memory[9147] <=  8'h64;        memory[9148] <=  8'h61;        memory[9149] <=  8'h61;        memory[9150] <=  8'h63;        memory[9151] <=  8'h61;        memory[9152] <=  8'h72;        memory[9153] <=  8'h63;        memory[9154] <=  8'h74;        memory[9155] <=  8'h72;        memory[9156] <=  8'h63;        memory[9157] <=  8'h61;        memory[9158] <=  8'h74;        memory[9159] <=  8'h72;        memory[9160] <=  8'h63;        memory[9161] <=  8'h61;        memory[9162] <=  8'h74;        memory[9163] <=  8'h63;        memory[9164] <=  8'h62;        memory[9165] <=  8'h61;        memory[9166] <=  8'h74;        memory[9167] <=  8'h62;        memory[9168] <=  8'h72;        memory[9169] <=  8'h63;        memory[9170] <=  8'h61;        memory[9171] <=  8'h74;        memory[9172] <=  8'h72;        memory[9173] <=  8'h6e;        memory[9174] <=  8'h62;        memory[9175] <=  8'h61;        memory[9176] <=  8'h63;        memory[9177] <=  8'h61;        memory[9178] <=  8'h74;        memory[9179] <=  8'h79;        memory[9180] <=  8'h73;        memory[9181] <=  8'h6e;        memory[9182] <=  8'h63;        memory[9183] <=  8'h74;        memory[9184] <=  8'h61;        memory[9185] <=  8'h6e;        memory[9186] <=  8'h62;        memory[9187] <=  8'h61;        memory[9188] <=  8'h63;        memory[9189] <=  8'h72;        memory[9190] <=  8'h6e;        memory[9191] <=  8'h74;        memory[9192] <=  8'h61;        memory[9193] <=  8'h62;        memory[9194] <=  8'h74;        memory[9195] <=  8'h6e;        memory[9196] <=  8'h61;        memory[9197] <=  8'h72;        memory[9198] <=  8'h62;        memory[9199] <=  8'h78;        memory[9200] <=  8'h74;        memory[9201] <=  8'h61;        memory[9202] <=  8'h72;        memory[9203] <=  8'h62;        memory[9204] <=  8'h61;        memory[9205] <=  8'h72;        memory[9206] <=  8'h74;        memory[9207] <=  8'h74;        memory[9208] <=  8'h62;        memory[9209] <=  8'h61;        memory[9210] <=  8'h72;        memory[9211] <=  8'h74;        memory[9212] <=  8'h78;        memory[9213] <=  8'h61;        memory[9214] <=  8'h74;        memory[9215] <=  8'h6b;        memory[9216] <=  8'h73;        memory[9217] <=  8'h68;        memory[9218] <=  8'h63;        memory[9219] <=  8'h66;        memory[9220] <=  8'h69;        memory[9221] <=  8'h77;        memory[9222] <=  8'h68;        memory[9223] <=  8'h61;        memory[9224] <=  8'h74;        memory[9225] <=  8'h61;        memory[9226] <=  8'h6e;        memory[9227] <=  8'h61;        memory[9228] <=  8'h62;        memory[9229] <=  8'h61;        memory[9230] <=  8'h63;        memory[9231] <=  8'h61;        memory[9232] <=  8'h74;        memory[9233] <=  8'h61;        memory[9234] <=  8'h62;        memory[9235] <=  8'h61;        memory[9236] <=  8'h72;        memory[9237] <=  8'h63;        memory[9238] <=  8'h61;        memory[9239] <=  8'h68;        memory[9240] <=  8'h64;        memory[9241] <=  8'h75;        memory[9242] <=  8'h63;        memory[9243] <=  8'h74;        memory[9244] <=  8'h61;        memory[9245] <=  8'h64;        memory[9246] <=  8'h61;        memory[9247] <=  8'h61;        memory[9248] <=  8'h63;        memory[9249] <=  8'h61;        memory[9250] <=  8'h72;        memory[9251] <=  8'h63;        memory[9252] <=  8'h74;        memory[9253] <=  8'h72;        memory[9254] <=  8'h63;        memory[9255] <=  8'h61;        memory[9256] <=  8'h74;        memory[9257] <=  8'h72;        memory[9258] <=  8'h63;        memory[9259] <=  8'h61;        memory[9260] <=  8'h74;        memory[9261] <=  8'h63;        memory[9262] <=  8'h62;        memory[9263] <=  8'h61;        memory[9264] <=  8'h74;        memory[9265] <=  8'h62;        memory[9266] <=  8'h72;        memory[9267] <=  8'h63;        memory[9268] <=  8'h61;        memory[9269] <=  8'h74;        memory[9270] <=  8'h72;        memory[9271] <=  8'h6e;        memory[9272] <=  8'h62;        memory[9273] <=  8'h61;        memory[9274] <=  8'h63;        memory[9275] <=  8'h61;        memory[9276] <=  8'h74;        memory[9277] <=  8'h79;        memory[9278] <=  8'h73;        memory[9279] <=  8'h6e;        memory[9280] <=  8'h63;        memory[9281] <=  8'h74;        memory[9282] <=  8'h61;        memory[9283] <=  8'h6e;        memory[9284] <=  8'h62;        memory[9285] <=  8'h61;        memory[9286] <=  8'h63;        memory[9287] <=  8'h72;        memory[9288] <=  8'h6e;        memory[9289] <=  8'h74;        memory[9290] <=  8'h61;        memory[9291] <=  8'h62;        memory[9292] <=  8'h74;        memory[9293] <=  8'h6e;        memory[9294] <=  8'h61;        memory[9295] <=  8'h72;        memory[9296] <=  8'h62;        memory[9297] <=  8'h78;        memory[9298] <=  8'h74;        memory[9299] <=  8'h61;        memory[9300] <=  8'h72;        memory[9301] <=  8'h5d;        memory[9302] <=  8'h5d;        memory[9303] <=  8'h65;        memory[9304] <=  8'h66;        memory[9305] <=  8'h77;        memory[9306] <=  8'h65;        memory[9307] <=  8'h5d;        memory[9308] <=  8'h65;        memory[9309] <=  8'h67;        memory[9310] <=  8'h73;        memory[9311] <=  8'h67;        memory[9312] <=  8'h66;        memory[9313] <=  8'h62;        memory[9314] <=  8'h61;        memory[9315] <=  8'h72;        memory[9316] <=  8'h74;        memory[9317] <=  8'h74;        memory[9318] <=  8'h62;        memory[9319] <=  8'h61;        memory[9320] <=  8'h72;        memory[9321] <=  8'h74;        memory[9322] <=  8'h78;        memory[9323] <=  8'h61;        memory[9324] <=  8'h74;        memory[9325] <=  8'h6b;        memory[9326] <=  8'h73;        memory[9327] <=  8'h68;        memory[9328] <=  8'h63;        memory[9329] <=  8'h66;        memory[9330] <=  8'h69;        memory[9331] <=  8'h77;        memory[9332] <=  8'h68;        memory[9333] <=  8'h61;        memory[9334] <=  8'h74;        memory[9335] <=  8'h61;        memory[9336] <=  8'h6e;        memory[9337] <=  8'h61;        memory[9338] <=  8'h62;        memory[9339] <=  8'h61;        memory[9340] <=  8'h63;        memory[9341] <=  8'h61;        memory[9342] <=  8'h74;        memory[9343] <=  8'h61;        memory[9344] <=  8'h62;        memory[9345] <=  8'h61;        memory[9346] <=  8'h72;        memory[9347] <=  8'h63;        memory[9348] <=  8'h61;        memory[9349] <=  8'h68;        memory[9350] <=  8'h64;        memory[9351] <=  8'h75;        memory[9352] <=  8'h63;        memory[9353] <=  8'h74;        memory[9354] <=  8'h61;        memory[9355] <=  8'h64;        memory[9356] <=  8'h61;        memory[9357] <=  8'h61;        memory[9358] <=  8'h63;        memory[9359] <=  8'h61;        memory[9360] <=  8'h72;        memory[9361] <=  8'h63;        memory[9362] <=  8'h74;        memory[9363] <=  8'h72;        memory[9364] <=  8'h63;        memory[9365] <=  8'h61;        memory[9366] <=  8'h74;        memory[9367] <=  8'h72;        memory[9368] <=  8'h63;        memory[9369] <=  8'h61;        memory[9370] <=  8'h74;        memory[9371] <=  8'h63;        memory[9372] <=  8'h62;        memory[9373] <=  8'h61;        memory[9374] <=  8'h74;        memory[9375] <=  8'h62;        memory[9376] <=  8'h72;        memory[9377] <=  8'h63;        memory[9378] <=  8'h61;        memory[9379] <=  8'h74;        memory[9380] <=  8'h72;        memory[9381] <=  8'h6e;        memory[9382] <=  8'h62;        memory[9383] <=  8'h61;        memory[9384] <=  8'h63;        memory[9385] <=  8'h61;        memory[9386] <=  8'h74;        memory[9387] <=  8'h79;        memory[9388] <=  8'h73;        memory[9389] <=  8'h6e;        memory[9390] <=  8'h63;        memory[9391] <=  8'h74;        memory[9392] <=  8'h61;        memory[9393] <=  8'h6e;        memory[9394] <=  8'h62;        memory[9395] <=  8'h61;        memory[9396] <=  8'h63;        memory[9397] <=  8'h72;        memory[9398] <=  8'h6e;        memory[9399] <=  8'h74;        memory[9400] <=  8'h61;        memory[9401] <=  8'h62;        memory[9402] <=  8'h74;        memory[9403] <=  8'h6e;        memory[9404] <=  8'h61;        memory[9405] <=  8'h72;        memory[9406] <=  8'h62;        memory[9407] <=  8'h78;        memory[9408] <=  8'h74;        memory[9409] <=  8'h61;        memory[9410] <=  8'h72;        memory[9411] <=  8'h62;        memory[9412] <=  8'h61;        memory[9413] <=  8'h72;        memory[9414] <=  8'h74;        memory[9415] <=  8'h74;        memory[9416] <=  8'h62;        memory[9417] <=  8'h61;        memory[9418] <=  8'h72;        memory[9419] <=  8'h74;        memory[9420] <=  8'h78;        memory[9421] <=  8'h61;        memory[9422] <=  8'h74;        memory[9423] <=  8'h6b;        memory[9424] <=  8'h73;        memory[9425] <=  8'h68;        memory[9426] <=  8'h63;        memory[9427] <=  8'h66;        memory[9428] <=  8'h69;        memory[9429] <=  8'h77;        memory[9430] <=  8'h68;        memory[9431] <=  8'h61;        memory[9432] <=  8'h74;        memory[9433] <=  8'h61;        memory[9434] <=  8'h6e;        memory[9435] <=  8'h61;        memory[9436] <=  8'h62;        memory[9437] <=  8'h61;        memory[9438] <=  8'h63;        memory[9439] <=  8'h61;        memory[9440] <=  8'h74;        memory[9441] <=  8'h61;        memory[9442] <=  8'h62;        memory[9443] <=  8'h61;        memory[9444] <=  8'h72;        memory[9445] <=  8'h63;        memory[9446] <=  8'h61;        memory[9447] <=  8'h68;        memory[9448] <=  8'h64;        memory[9449] <=  8'h75;        memory[9450] <=  8'h63;        memory[9451] <=  8'h74;        memory[9452] <=  8'h61;        memory[9453] <=  8'h64;        memory[9454] <=  8'h61;        memory[9455] <=  8'h61;        memory[9456] <=  8'h63;        memory[9457] <=  8'h61;        memory[9458] <=  8'h72;        memory[9459] <=  8'h63;        memory[9460] <=  8'h74;        memory[9461] <=  8'h72;        memory[9462] <=  8'h63;        memory[9463] <=  8'h61;        memory[9464] <=  8'h74;        memory[9465] <=  8'h72;        memory[9466] <=  8'h63;        memory[9467] <=  8'h61;        memory[9468] <=  8'h74;        memory[9469] <=  8'h63;        memory[9470] <=  8'h62;        memory[9471] <=  8'h61;        memory[9472] <=  8'h74;        memory[9473] <=  8'h62;        memory[9474] <=  8'h72;        memory[9475] <=  8'h63;        memory[9476] <=  8'h61;        memory[9477] <=  8'h74;        memory[9478] <=  8'h72;        memory[9479] <=  8'h6e;        memory[9480] <=  8'h62;        memory[9481] <=  8'h61;        memory[9482] <=  8'h63;        memory[9483] <=  8'h61;        memory[9484] <=  8'h74;        memory[9485] <=  8'h79;        memory[9486] <=  8'h73;        memory[9487] <=  8'h6e;        memory[9488] <=  8'h63;        memory[9489] <=  8'h74;        memory[9490] <=  8'h61;        memory[9491] <=  8'h6e;        memory[9492] <=  8'h62;        memory[9493] <=  8'h61;        memory[9494] <=  8'h63;        memory[9495] <=  8'h72;        memory[9496] <=  8'h6e;        memory[9497] <=  8'h74;        memory[9498] <=  8'h61;        memory[9499] <=  8'h62;        memory[9500] <=  8'h74;        memory[9501] <=  8'h6e;        memory[9502] <=  8'h61;        memory[9503] <=  8'h72;        memory[9504] <=  8'h62;        memory[9505] <=  8'h78;        memory[9506] <=  8'h74;        memory[9507] <=  8'h61;        memory[9508] <=  8'h72;        memory[9509] <=  8'h64;        memory[9510] <=  8'h66;        memory[9511] <=  8'h73;        memory[9512] <=  8'h67;        memory[9513] <=  8'h76;        memory[9514] <=  8'h68;        memory[9515] <=  8'h62;        memory[9516] <=  8'h6b;        memory[9517] <=  8'h6a;        memory[9518] <=  8'h6e;        memory[9519] <=  8'h6d;        memory[9520] <=  8'h62;        memory[9521] <=  8'h76;        memory[9522] <=  8'h78;        memory[9523] <=  8'h63;        memory[9524] <=  8'h73;        memory[9525] <=  8'h66;        memory[9526] <=  8'h72;        memory[9527] <=  8'h74;        memory[9528] <=  8'h79;        memory[9529] <=  8'h75;        memory[9530] <=  8'h6a;        memory[9531] <=  8'h6e;        memory[9532] <=  8'h62;        memory[9533] <=  8'h76;        memory[9534] <=  8'h63;        memory[9535] <=  8'h64;        memory[9536] <=  8'h74;        memory[9537] <=  8'h79;        memory[9538] <=  8'h75;        memory[9539] <=  8'h69;        memory[9540] <=  8'h6b;        memory[9541] <=  8'h6d;        memory[9542] <=  8'h6e;        memory[9543] <=  8'h62;        memory[9544] <=  8'h76;        memory[9545] <=  8'h63;        memory[9546] <=  8'h78;        memory[9547] <=  8'h73;        memory[9548] <=  8'h64;        memory[9549] <=  8'h72;        memory[9550] <=  8'h74;        memory[9551] <=  8'h79;        memory[9552] <=  8'h75;        memory[9553] <=  8'h69;        memory[9554] <=  8'h6b;        memory[9555] <=  8'h6d;        memory[9556] <=  8'h6e;        memory[9557] <=  8'h62;        memory[9558] <=  8'h76;        memory[9559] <=  8'h63;        memory[9560] <=  8'h73;        memory[9561] <=  8'h77;        memory[9562] <=  8'h33;        memory[9563] <=  8'h34;        memory[9564] <=  8'h35;        memory[9565] <=  8'h36;        memory[9566] <=  8'h37;        memory[9567] <=  8'h38;        memory[9568] <=  8'h69;        memory[9569] <=  8'h6b;        memory[9570] <=  8'h6d;        memory[9571] <=  8'h6e;        memory[9572] <=  8'h62;        memory[9573] <=  8'h76;        memory[9574] <=  8'h63;        memory[9575] <=  8'h64;        memory[9576] <=  8'h65;        memory[9577] <=  8'h72;        memory[9578] <=  8'h36;        memory[9579] <=  8'h37;        memory[9580] <=  8'h38;        memory[9581] <=  8'h69;        memory[9582] <=  8'h6f;        memory[9583] <=  8'h6b;        memory[9584] <=  8'h6a;        memory[9585] <=  8'h6e;        memory[9586] <=  8'h62;        memory[9587] <=  8'h76;        memory[9588] <=  8'h63;        memory[9589] <=  8'h64;        memory[9590] <=  8'h72;        memory[9591] <=  8'h74;        memory[9592] <=  8'h79;        memory[9593] <=  8'h75;        memory[9594] <=  8'h73;        memory[9595] <=  8'h6a;        memory[9596] <=  8'h63;        memory[9597] <=  8'h6e;        memory[9598] <=  8'h62;        memory[9599] <=  8'h64;        memory[9600] <=  8'h66;        memory[9601] <=  8'h73;        memory[9602] <=  8'h74;        memory[9603] <=  8'h79;        memory[9604] <=  8'h75;        memory[9605] <=  8'h61;        memory[9606] <=  8'h69;        memory[9607] <=  8'h6b;        memory[9608] <=  8'h78;        memory[9609] <=  8'h6d;        memory[9610] <=  8'h6e;        memory[9611] <=  8'h73;        memory[9612] <=  8'h6a;        memory[9613] <=  8'h6f;        memory[9614] <=  8'h64;        memory[9615] <=  8'h6c;        memory[9616] <=  8'h63;        memory[9617] <=  8'h78;        memory[9618] <=  8'h62;        memory[9619] <=  8'h61;        memory[9620] <=  8'h72;        memory[9621] <=  8'h74;        memory[9622] <=  8'h78;        memory[9623] <=  8'h61;        memory[9624] <=  8'h74;        memory[9625] <=  8'h6b;        memory[9626] <=  8'h73;        memory[9627] <=  8'h68;        memory[9628] <=  8'h63;        memory[9629] <=  8'h66;        memory[9630] <=  8'h69;        memory[9631] <=  8'h77;        memory[9632] <=  8'h68;        memory[9633] <=  8'h61;        memory[9634] <=  8'h74;        memory[9635] <=  8'h61;        memory[9636] <=  8'h6e;        memory[9637] <=  8'h61;        memory[9638] <=  8'h62;        memory[9639] <=  8'h61;        memory[9640] <=  8'h63;        memory[9641] <=  8'h61;        memory[9642] <=  8'h74;        memory[9643] <=  8'h61;        memory[9644] <=  8'h62;        memory[9645] <=  8'h61;        memory[9646] <=  8'h72;        memory[9647] <=  8'h63;        memory[9648] <=  8'h61;        memory[9649] <=  8'h68;        memory[9650] <=  8'h64;        memory[9651] <=  8'h75;        memory[9652] <=  8'h63;        memory[9653] <=  8'h74;        memory[9654] <=  8'h61;        memory[9655] <=  8'h64;        memory[9656] <=  8'h61;        memory[9657] <=  8'h61;        memory[9658] <=  8'h63;        memory[9659] <=  8'h61;        memory[9660] <=  8'h72;        memory[9661] <=  8'h62;        memory[9662] <=  8'h61;        memory[9663] <=  8'h72;        memory[9664] <=  8'h74;        memory[9665] <=  8'h78;        memory[9666] <=  8'h61;        memory[9667] <=  8'h74;        memory[9668] <=  8'h6b;        memory[9669] <=  8'h73;        memory[9670] <=  8'h68;        memory[9671] <=  8'h63;        memory[9672] <=  8'h66;        memory[9673] <=  8'h69;        memory[9674] <=  8'h77;        memory[9675] <=  8'h68;        memory[9676] <=  8'h61;        memory[9677] <=  8'h74;        memory[9678] <=  8'h61;        memory[9679] <=  8'h6e;        memory[9680] <=  8'h61;        memory[9681] <=  8'h62;        memory[9682] <=  8'h61;        memory[9683] <=  8'h63;        memory[9684] <=  8'h61;        memory[9685] <=  8'h74;        memory[9686] <=  8'h61;        memory[9687] <=  8'h62;        memory[9688] <=  8'h61;        memory[9689] <=  8'h72;        memory[9690] <=  8'h63;        memory[9691] <=  8'h61;        memory[9692] <=  8'h68;        memory[9693] <=  8'h64;        memory[9694] <=  8'h75;        memory[9695] <=  8'h63;        memory[9696] <=  8'h74;        memory[9697] <=  8'h61;        memory[9698] <=  8'h64;        memory[9699] <=  8'h61;        memory[9700] <=  8'h61;        memory[9701] <=  8'h63;        memory[9702] <=  8'h61;        memory[9703] <=  8'h72;        memory[9704] <=  8'h62;        memory[9705] <=  8'h61;        memory[9706] <=  8'h72;        memory[9707] <=  8'h74;        memory[9708] <=  8'h78;        memory[9709] <=  8'h61;        memory[9710] <=  8'h74;        memory[9711] <=  8'h6b;        memory[9712] <=  8'h73;        memory[9713] <=  8'h68;        memory[9714] <=  8'h63;        memory[9715] <=  8'h66;        memory[9716] <=  8'h69;        memory[9717] <=  8'h77;        memory[9718] <=  8'h68;        memory[9719] <=  8'h61;        memory[9720] <=  8'h74;        memory[9721] <=  8'h61;        memory[9722] <=  8'h6e;        memory[9723] <=  8'h61;        memory[9724] <=  8'h62;        memory[9725] <=  8'h61;        memory[9726] <=  8'h63;        memory[9727] <=  8'h61;        memory[9728] <=  8'h74;        memory[9729] <=  8'h61;        memory[9730] <=  8'h62;        memory[9731] <=  8'h61;        memory[9732] <=  8'h72;        memory[9733] <=  8'h63;        memory[9734] <=  8'h61;        memory[9735] <=  8'h68;        memory[9736] <=  8'h64;        memory[9737] <=  8'h75;        memory[9738] <=  8'h63;        memory[9739] <=  8'h74;        memory[9740] <=  8'h61;        memory[9741] <=  8'h64;        memory[9742] <=  8'h61;        memory[9743] <=  8'h61;        memory[9744] <=  8'h63;        memory[9745] <=  8'h61;        memory[9746] <=  8'h72;        memory[9747] <=  8'h62;        memory[9748] <=  8'h61;        memory[9749] <=  8'h72;        memory[9750] <=  8'h74;        memory[9751] <=  8'h78;        memory[9752] <=  8'h61;        memory[9753] <=  8'h74;        memory[9754] <=  8'h6b;        memory[9755] <=  8'h73;        memory[9756] <=  8'h68;        memory[9757] <=  8'h63;        memory[9758] <=  8'h66;        memory[9759] <=  8'h69;        memory[9760] <=  8'h77;        memory[9761] <=  8'h68;        memory[9762] <=  8'h61;        memory[9763] <=  8'h74;        memory[9764] <=  8'h61;        memory[9765] <=  8'h6e;        memory[9766] <=  8'h61;        memory[9767] <=  8'h62;        memory[9768] <=  8'h61;        memory[9769] <=  8'h63;        memory[9770] <=  8'h61;        memory[9771] <=  8'h74;        memory[9772] <=  8'h61;        memory[9773] <=  8'h62;        memory[9774] <=  8'h61;        memory[9775] <=  8'h72;        memory[9776] <=  8'h63;        memory[9777] <=  8'h61;        memory[9778] <=  8'h68;        memory[9779] <=  8'h64;        memory[9780] <=  8'h75;        memory[9781] <=  8'h63;        memory[9782] <=  8'h74;        memory[9783] <=  8'h61;        memory[9784] <=  8'h64;        memory[9785] <=  8'h61;        memory[9786] <=  8'h61;        memory[9787] <=  8'h63;        memory[9788] <=  8'h61;        memory[9789] <=  8'h72;        memory[9790] <=  8'h62;        memory[9791] <=  8'h61;        memory[9792] <=  8'h72;        memory[9793] <=  8'h74;        memory[9794] <=  8'h78;        memory[9795] <=  8'h61;        memory[9796] <=  8'h74;        memory[9797] <=  8'h6b;        memory[9798] <=  8'h73;        memory[9799] <=  8'h68;        memory[9800] <=  8'h63;        memory[9801] <=  8'h66;        memory[9802] <=  8'h69;        memory[9803] <=  8'h77;        memory[9804] <=  8'h68;        memory[9805] <=  8'h61;        memory[9806] <=  8'h74;        memory[9807] <=  8'h61;        memory[9808] <=  8'h6e;        memory[9809] <=  8'h61;        memory[9810] <=  8'h62;        memory[9811] <=  8'h61;        memory[9812] <=  8'h63;        memory[9813] <=  8'h61;        memory[9814] <=  8'h74;        memory[9815] <=  8'h61;        memory[9816] <=  8'h62;        memory[9817] <=  8'h61;        memory[9818] <=  8'h72;        memory[9819] <=  8'h63;        memory[9820] <=  8'h61;        memory[9821] <=  8'h68;        memory[9822] <=  8'h64;        memory[9823] <=  8'h75;        memory[9824] <=  8'h63;        memory[9825] <=  8'h74;        memory[9826] <=  8'h61;        memory[9827] <=  8'h64;        memory[9828] <=  8'h61;        memory[9829] <=  8'h61;        memory[9830] <=  8'h63;        memory[9831] <=  8'h61;        memory[9832] <=  8'h72;        memory[9833] <=  8'h62;        memory[9834] <=  8'h61;        memory[9835] <=  8'h72;        memory[9836] <=  8'h74;        memory[9837] <=  8'h78;        memory[9838] <=  8'h61;        memory[9839] <=  8'h74;        memory[9840] <=  8'h6b;        memory[9841] <=  8'h73;        memory[9842] <=  8'h68;        memory[9843] <=  8'h63;        memory[9844] <=  8'h66;        memory[9845] <=  8'h69;        memory[9846] <=  8'h77;        memory[9847] <=  8'h68;        memory[9848] <=  8'h61;        memory[9849] <=  8'h74;        memory[9850] <=  8'h61;        memory[9851] <=  8'h6e;        memory[9852] <=  8'h61;        memory[9853] <=  8'h62;        memory[9854] <=  8'h61;        memory[9855] <=  8'h63;        memory[9856] <=  8'h61;        memory[9857] <=  8'h74;        memory[9858] <=  8'h61;        memory[9859] <=  8'h62;        memory[9860] <=  8'h61;        memory[9861] <=  8'h72;        memory[9862] <=  8'h63;        memory[9863] <=  8'h61;        memory[9864] <=  8'h68;        memory[9865] <=  8'h64;        memory[9866] <=  8'h75;        memory[9867] <=  8'h63;        memory[9868] <=  8'h74;        memory[9869] <=  8'h61;        memory[9870] <=  8'h64;        memory[9871] <=  8'h61;        memory[9872] <=  8'h61;        memory[9873] <=  8'h63;        memory[9874] <=  8'h61;        memory[9875] <=  8'h72;        memory[9876] <=  8'h62;        memory[9877] <=  8'h61;        memory[9878] <=  8'h72;        memory[9879] <=  8'h74;        memory[9880] <=  8'h78;        memory[9881] <=  8'h61;        memory[9882] <=  8'h74;        memory[9883] <=  8'h6b;        memory[9884] <=  8'h73;        memory[9885] <=  8'h68;        memory[9886] <=  8'h63;        memory[9887] <=  8'h66;        memory[9888] <=  8'h69;        memory[9889] <=  8'h77;        memory[9890] <=  8'h68;        memory[9891] <=  8'h61;        memory[9892] <=  8'h74;        memory[9893] <=  8'h61;        memory[9894] <=  8'h6e;        memory[9895] <=  8'h61;        memory[9896] <=  8'h62;        memory[9897] <=  8'h61;        memory[9898] <=  8'h63;        memory[9899] <=  8'h61;        memory[9900] <=  8'h74;        memory[9901] <=  8'h61;        memory[9902] <=  8'h62;        memory[9903] <=  8'h61;        memory[9904] <=  8'h72;        memory[9905] <=  8'h63;        memory[9906] <=  8'h61;        memory[9907] <=  8'h68;        memory[9908] <=  8'h64;        memory[9909] <=  8'h75;        memory[9910] <=  8'h63;        memory[9911] <=  8'h74;        memory[9912] <=  8'h61;        memory[9913] <=  8'h64;        memory[9914] <=  8'h61;        memory[9915] <=  8'h61;        memory[9916] <=  8'h63;        memory[9917] <=  8'h61;        memory[9918] <=  8'h72;        memory[9919] <=  8'h62;        memory[9920] <=  8'h61;        memory[9921] <=  8'h72;        memory[9922] <=  8'h74;        memory[9923] <=  8'h78;        memory[9924] <=  8'h61;        memory[9925] <=  8'h74;        memory[9926] <=  8'h6b;        memory[9927] <=  8'h73;        memory[9928] <=  8'h68;        memory[9929] <=  8'h63;        memory[9930] <=  8'h66;        memory[9931] <=  8'h69;        memory[9932] <=  8'h77;        memory[9933] <=  8'h68;        memory[9934] <=  8'h61;        memory[9935] <=  8'h74;        memory[9936] <=  8'h61;        memory[9937] <=  8'h6e;        memory[9938] <=  8'h61;        memory[9939] <=  8'h62;        memory[9940] <=  8'h61;        memory[9941] <=  8'h63;        memory[9942] <=  8'h61;        memory[9943] <=  8'h74;        memory[9944] <=  8'h61;        memory[9945] <=  8'h62;        memory[9946] <=  8'h61;        memory[9947] <=  8'h72;        memory[9948] <=  8'h63;        memory[9949] <=  8'h61;        memory[9950] <=  8'h68;        memory[9951] <=  8'h64;        memory[9952] <=  8'h75;        memory[9953] <=  8'h63;        memory[9954] <=  8'h74;        memory[9955] <=  8'h61;        memory[9956] <=  8'h64;        memory[9957] <=  8'h61;        memory[9958] <=  8'h61;        memory[9959] <=  8'h63;        memory[9960] <=  8'h61;        memory[9961] <=  8'h72;        memory[9962] <=  8'h62;        memory[9963] <=  8'h61;        memory[9964] <=  8'h72;        memory[9965] <=  8'h74;        memory[9966] <=  8'h78;        memory[9967] <=  8'h61;        memory[9968] <=  8'h74;        memory[9969] <=  8'h6b;        memory[9970] <=  8'h73;        memory[9971] <=  8'h68;        memory[9972] <=  8'h63;        memory[9973] <=  8'h66;        memory[9974] <=  8'h69;        memory[9975] <=  8'h77;        memory[9976] <=  8'h68;        memory[9977] <=  8'h61;        memory[9978] <=  8'h74;        memory[9979] <=  8'h61;        memory[9980] <=  8'h6e;        memory[9981] <=  8'h61;        memory[9982] <=  8'h62;        memory[9983] <=  8'h61;        memory[9984] <=  8'h63;        memory[9985] <=  8'h61;        memory[9986] <=  8'h74;        memory[9987] <=  8'h61;        memory[9988] <=  8'h62;        memory[9989] <=  8'h61;        memory[9990] <=  8'h72;        memory[9991] <=  8'h63;        memory[9992] <=  8'h61;        memory[9993] <=  8'h68;        memory[9994] <=  8'h64;        memory[9995] <=  8'h75;        memory[9996] <=  8'h63;        memory[9997] <=  8'h74;        memory[9998] <=  8'h61;        memory[9999] <=  8'h64;        memory[10000] <=  8'h61;        memory[10001] <=  8'h61;        memory[10002] <=  8'h63;        memory[10003] <=  8'h61;        memory[10004] <=  8'h72;        memory[10005] <=  8'h62;        memory[10006] <=  8'h61;        memory[10007] <=  8'h72;        memory[10008] <=  8'h74;        memory[10009] <=  8'h74;        memory[10010] <=  8'h62;        memory[10011] <=  8'h61;        memory[10012] <=  8'h72;        memory[10013] <=  8'h74;        memory[10014] <=  8'h78;        memory[10015] <=  8'h61;        memory[10016] <=  8'h74;        memory[10017] <=  8'h6b;        memory[10018] <=  8'h73;        memory[10019] <=  8'h68;        memory[10020] <=  8'h63;        memory[10021] <=  8'h66;        memory[10022] <=  8'h69;        memory[10023] <=  8'h77;        memory[10024] <=  8'h68;        memory[10025] <=  8'h61;        memory[10026] <=  8'h74;        memory[10027] <=  8'h61;        memory[10028] <=  8'h6e;        memory[10029] <=  8'h61;        memory[10030] <=  8'h62;        memory[10031] <=  8'h61;        memory[10032] <=  8'h63;        memory[10033] <=  8'h61;        memory[10034] <=  8'h74;        memory[10035] <=  8'h61;        memory[10036] <=  8'h62;        memory[10037] <=  8'h61;        memory[10038] <=  8'h72;        memory[10039] <=  8'h63;        memory[10040] <=  8'h61;        memory[10041] <=  8'h68;        memory[10042] <=  8'h64;        memory[10043] <=  8'h75;        memory[10044] <=  8'h63;        memory[10045] <=  8'h74;        memory[10046] <=  8'h61;        memory[10047] <=  8'h64;        memory[10048] <=  8'h61;        memory[10049] <=  8'h61;        memory[10050] <=  8'h63;        memory[10051] <=  8'h61;        memory[10052] <=  8'h72;        memory[10053] <=  8'h63;        memory[10054] <=  8'h74;        memory[10055] <=  8'h72;        memory[10056] <=  8'h63;        memory[10057] <=  8'h61;        memory[10058] <=  8'h74;        memory[10059] <=  8'h72;        memory[10060] <=  8'h63;        memory[10061] <=  8'h61;        memory[10062] <=  8'h74;        memory[10063] <=  8'h63;        memory[10064] <=  8'h62;        memory[10065] <=  8'h61;        memory[10066] <=  8'h74;        memory[10067] <=  8'h62;        memory[10068] <=  8'h72;        memory[10069] <=  8'h63;        memory[10070] <=  8'h61;        memory[10071] <=  8'h72;        memory[10072] <=  8'h62;        memory[10073] <=  8'h78;        memory[10074] <=  8'h74;        memory[10075] <=  8'h61;        memory[10076] <=  8'h72;        memory[10077] <=  8'h64;        memory[10078] <=  8'h66;        memory[10079] <=  8'h73;        memory[10080] <=  8'h67;        memory[10081] <=  8'h76;        memory[10082] <=  8'h68;        memory[10083] <=  8'h62;        memory[10084] <=  8'h6b;        memory[10085] <=  8'h6a;        memory[10086] <=  8'h6e;        memory[10087] <=  8'h6d;        memory[10088] <=  8'h62;        memory[10089] <=  8'h76;        memory[10090] <=  8'h78;        memory[10091] <=  8'h63;        memory[10092] <=  8'h73;        memory[10093] <=  8'h66;        memory[10094] <=  8'h72;        memory[10095] <=  8'h74;        memory[10096] <=  8'h79;        memory[10097] <=  8'h75;        memory[10098] <=  8'h6a;        memory[10099] <=  8'h6e;        memory[10100] <=  8'h62;        memory[10101] <=  8'h76;        memory[10102] <=  8'h63;        memory[10103] <=  8'h64;        memory[10104] <=  8'h74;        memory[10105] <=  8'h79;        memory[10106] <=  8'h75;        memory[10107] <=  8'h69;        memory[10108] <=  8'h6b;        memory[10109] <=  8'h6d;        memory[10110] <=  8'h6e;        memory[10111] <=  8'h62;        memory[10112] <=  8'h76;        memory[10113] <=  8'h63;        memory[10114] <=  8'h78;        memory[10115] <=  8'h73;        memory[10116] <=  8'h64;        memory[10117] <=  8'h72;        memory[10118] <=  8'h74;        memory[10119] <=  8'h79;        memory[10120] <=  8'h75;        memory[10121] <=  8'h69;        memory[10122] <=  8'h6b;        memory[10123] <=  8'h6d;        memory[10124] <=  8'h6e;        memory[10125] <=  8'h62;        memory[10126] <=  8'h76;        memory[10127] <=  8'h63;        memory[10128] <=  8'h73;        memory[10129] <=  8'h77;        memory[10130] <=  8'h33;        memory[10131] <=  8'h34;        memory[10132] <=  8'h35;        memory[10133] <=  8'h36;        memory[10134] <=  8'h37;        memory[10135] <=  8'h38;        memory[10136] <=  8'h69;        memory[10137] <=  8'h6b;        memory[10138] <=  8'h6d;        memory[10139] <=  8'h6e;        memory[10140] <=  8'h62;        memory[10141] <=  8'h76;        memory[10142] <=  8'h63;        memory[10143] <=  8'h64;        memory[10144] <=  8'h65;        memory[10145] <=  8'h72;        memory[10146] <=  8'h36;        memory[10147] <=  8'h37;        memory[10148] <=  8'h38;        memory[10149] <=  8'h69;        memory[10150] <=  8'h6f;        memory[10151] <=  8'h6b;        memory[10152] <=  8'h6a;        memory[10153] <=  8'h6e;        memory[10154] <=  8'h62;        memory[10155] <=  8'h76;        memory[10156] <=  8'h63;        memory[10157] <=  8'h64;        memory[10158] <=  8'h72;        memory[10159] <=  8'h74;        memory[10160] <=  8'h79;        memory[10161] <=  8'h75;        memory[10162] <=  8'h73;        memory[10163] <=  8'h6a;        memory[10164] <=  8'h63;        memory[10165] <=  8'h6e;        memory[10166] <=  8'h62;        memory[10167] <=  8'h64;        memory[10168] <=  8'h66;        memory[10169] <=  8'h73;        memory[10170] <=  8'h74;        memory[10171] <=  8'h79;        memory[10172] <=  8'h75;        memory[10173] <=  8'h61;        memory[10174] <=  8'h69;        memory[10175] <=  8'h6b;        memory[10176] <=  8'h78;        memory[10177] <=  8'h6d;        memory[10178] <=  8'h6e;        memory[10179] <=  8'h73;        memory[10180] <=  8'h6a;        memory[10181] <=  8'h6f;        memory[10182] <=  8'h64;        memory[10183] <=  8'h6c;        memory[10184] <=  8'h63;        memory[10185] <=  8'h78;        memory[10186] <=  8'h2c;        memory[10187] <=  8'h6d;        memory[10188] <=  8'h73;        memory[10189] <=  8'h6b;        memory[10190] <=  8'h64;        memory[10191] <=  8'h6c;        memory[10192] <=  8'h70;        memory[10193] <=  8'h5b;        memory[10194] <=  8'h3b;        memory[10195] <=  8'h73;        memory[10196] <=  8'h6c;        memory[10197] <=  8'h64;        memory[10198] <=  8'h70;        memory[10199] <=  8'h76;        memory[10200] <=  8'h63;        memory[10201] <=  8'h5b;        memory[10202] <=  8'h78;        memory[10203] <=  8'h76;        memory[10204] <=  8'h63;        memory[10205] <=  8'h5b;        memory[10206] <=  8'h78;        memory[10207] <=  8'h70;        memory[10208] <=  8'h6f;        memory[10209] <=  8'h20;        memory[10210] <=  8'h62;        memory[10211] <=  8'h61;        memory[10212] <=  8'h72;        memory[10213] <=  8'h74;        memory[10214] <=  8'h74;        memory[10215] <=  8'h62;        memory[10216] <=  8'h61;        memory[10217] <=  8'h72;        memory[10218] <=  8'h74;        memory[10219] <=  8'h78;        memory[10220] <=  8'h61;        memory[10221] <=  8'h74;        memory[10222] <=  8'h6b;        memory[10223] <=  8'h73;        memory[10224] <=  8'h68;        memory[10225] <=  8'h63;        memory[10226] <=  8'h66;        memory[10227] <=  8'h69;        memory[10228] <=  8'h77;        memory[10229] <=  8'h68;        memory[10230] <=  8'h61;        memory[10231] <=  8'h69;        memory[10232] <=  8'h6a;        memory[10233] <=  8'h78;        memory[10234] <=  8'h5d;        memory[10235] <=  8'h65;        memory[10236] <=  8'h6b;        memory[10237] <=  8'h6f;        memory[10238] <=  8'h39;        memory[10239] <=  8'h64;        memory[10240] <=  8'h75;        memory[10241] <=  8'h38;        memory[10242] <=  8'h79;        memory[10243] <=  8'h20;        memory[10244] <=  8'h37;        memory[10245] <=  8'h63;        memory[10246] <=  8'h67;        memory[10247] <=  8'h78;        memory[10248] <=  8'h63;        memory[10249] <=  8'h75;        memory[10250] <=  8'h68;        memory[10251] <=  8'h69;        memory[10252] <=  8'h6a;        memory[10253] <=  8'h77;        memory[10254] <=  8'h69;        memory[10255] <=  8'h64;        memory[10256] <=  8'h66;        memory[10257] <=  8'h68;        memory[10258] <=  8'h75;        memory[10259] <=  8'h76;        memory[10260] <=  8'h64;        memory[10261] <=  8'h62;        memory[10262] <=  8'h66;        memory[10263] <=  8'h6a;        memory[10264] <=  8'h6e;        memory[10265] <=  8'h6b;        memory[10266] <=  8'h6a;        memory[10267] <=  8'h65;        memory[10268] <=  8'h38;        memory[10269] <=  8'h66;        memory[10270] <=  8'h37;        memory[10271] <=  8'h67;        memory[10272] <=  8'h79;        memory[10273] <=  8'h76;        memory[10274] <=  8'h63;        memory[10275] <=  8'h68;        memory[10276] <=  8'h69;        memory[10277] <=  8'h6a;        memory[10278] <=  8'h33;        memory[10279] <=  8'h65;        memory[10280] <=  8'h67;        memory[10281] <=  8'h79;        memory[10282] <=  8'h72;        memory[10283] <=  8'h64;        memory[10284] <=  8'h62;        memory[10285] <=  8'h6e;        memory[10286] <=  8'h63;        memory[10287] <=  8'h7a;        memory[10288] <=  8'h6a;        memory[10289] <=  8'h6f;        memory[10290] <=  8'h66;        memory[10291] <=  8'h78;        memory[10292] <=  8'h6a;        memory[10293] <=  8'h69;        memory[10294] <=  8'h63;        memory[10295] <=  8'h68;        memory[10296] <=  8'h62;        memory[10297] <=  8'h6e;        memory[10298] <=  8'h6d;        memory[10299] <=  8'h63;        memory[10300] <=  8'h73;        memory[10301] <=  8'h6c;        memory[10302] <=  8'h6b;        memory[10303] <=  8'h6a;        memory[10304] <=  8'h69;        memory[10305] <=  8'h68;        memory[10306] <=  8'h76;        memory[10307] <=  8'h75;        memory[10308] <=  8'h69;        memory[10309] <=  8'h64;        memory[10310] <=  8'h68;        memory[10311] <=  8'h75;        memory[10312] <=  8'h67;        memory[10313] <=  8'h79;        memory[10314] <=  8'h62;        memory[10315] <=  8'h68;        memory[10316] <=  8'h65;        memory[10317] <=  8'h6a;        memory[10318] <=  8'h72;        memory[10319] <=  8'h6b;        memory[10320] <=  8'h6a;        memory[10321] <=  8'h6f;        memory[10322] <=  8'h64;        memory[10323] <=  8'h67;        memory[10324] <=  8'h69;        memory[10325] <=  8'h75;        memory[10326] <=  8'h69;        memory[10327] <=  8'h67;        memory[10328] <=  8'h76;        memory[10329] <=  8'h79;        memory[10330] <=  8'h75;        memory[10331] <=  8'h67;        memory[10332] <=  8'h78;        memory[10333] <=  8'h68;        memory[10334] <=  8'h63;        memory[10335] <=  8'h20;        memory[10336] <=  8'h20;        memory[10337] <=  8'h20;        memory[10338] <=  8'h78;        memory[10339] <=  8'h76;        memory[10340] <=  8'h20;        memory[10341] <=  8'h63;        memory[10342] <=  8'h78;        memory[10343] <=  8'h67;        memory[10344] <=  8'h79;        memory[10345] <=  8'h63;        memory[10346] <=  8'h75;        memory[10347] <=  8'h68;        memory[10348] <=  8'h6a;        memory[10349] <=  8'h6b;        memory[10350] <=  8'h61;        memory[10351] <=  8'h6c;        memory[10352] <=  8'h78;        memory[10353] <=  8'h76;        memory[10354] <=  8'h70;        memory[10355] <=  8'h6f;        memory[10356] <=  8'h69;        memory[10357] <=  8'h6a;        memory[10358] <=  8'h69;        memory[10359] <=  8'h68;        memory[10360] <=  8'h6a;        memory[10361] <=  8'h62;        memory[10362] <=  8'h77;        memory[10363] <=  8'h65;        memory[10364] <=  8'h6e;        memory[10365] <=  8'h61;        memory[10366] <=  8'h66;        memory[10367] <=  8'h6d;        memory[10368] <=  8'h64;        memory[10369] <=  8'h6b;        memory[10370] <=  8'h6d;        memory[10371] <=  8'h76;        memory[10372] <=  8'h6c;        memory[10373] <=  8'h63;        memory[10374] <=  8'h6f;        memory[10375] <=  8'h64;        memory[10376] <=  8'h69;        memory[10377] <=  8'h75;        memory[10378] <=  8'h68;        memory[10379] <=  8'h73;        memory[10380] <=  8'h66;        memory[10381] <=  8'h65;        memory[10382] <=  8'h62;        memory[10383] <=  8'h6e;        memory[10384] <=  8'h64;        memory[10385] <=  8'h73;        memory[10386] <=  8'h63;        memory[10387] <=  8'h6b;        memory[10388] <=  8'h20;        memory[10389] <=  8'h78;        memory[10390] <=  8'h6a;        memory[10391] <=  8'h78;        memory[10392] <=  8'h63;        memory[10393] <=  8'h73;        memory[10394] <=  8'h64;        memory[10395] <=  8'h66;        memory[10396] <=  8'h6b;        memory[10397] <=  8'h64;        memory[10398] <=  8'h6e;        memory[10399] <=  8'h6d;        memory[10400] <=  8'h64;        memory[10401] <=  8'h73;        memory[10402] <=  8'h63;        memory[10403] <=  8'h6b;        memory[10404] <=  8'h78;        memory[10405] <=  8'h6c;        memory[10406] <=  8'h6f;        memory[10407] <=  8'h66;        memory[10408] <=  8'h6a;        memory[10409] <=  8'h69;        memory[10410] <=  8'h61;        memory[10411] <=  8'h62;        memory[10412] <=  8'h6e;        memory[10413] <=  8'h20;        memory[10414] <=  8'h78;        memory[10415] <=  8'h6b;        memory[10416] <=  8'h6d;        memory[10417] <=  8'h20;        memory[10418] <=  8'h6f;        memory[10419] <=  8'h63;        memory[10420] <=  8'h76;        memory[10421] <=  8'h73;        memory[10422] <=  8'h64;        memory[10423] <=  8'h69;        memory[10424] <=  8'h66;        memory[10425] <=  8'h68;        memory[10426] <=  8'h65;        memory[10427] <=  8'h71;        memory[10428] <=  8'h6a;        memory[10429] <=  8'h77;        memory[10430] <=  8'h62;        memory[10431] <=  8'h65;        memory[10432] <=  8'h6e;        memory[10433] <=  8'h20;        memory[10434] <=  8'h6d;        memory[10435] <=  8'h64;        memory[10436] <=  8'h73;        memory[10437] <=  8'h6c;        memory[10438] <=  8'h76;        memory[10439] <=  8'h6b;        memory[10440] <=  8'h63;        memory[10441] <=  8'h78;        memory[10442] <=  8'h20;        memory[10443] <=  8'h6f;        memory[10444] <=  8'h78;        memory[10445] <=  8'h69;        memory[10446] <=  8'h63;        memory[10447] <=  8'h6a;        memory[10448] <=  8'h76;        memory[10449] <=  8'h64;        memory[10450] <=  8'h66;        memory[10451] <=  8'h65;        memory[10452] <=  8'h71;        memory[10453] <=  8'h6e;        memory[10454] <=  8'h20;        memory[10455] <=  8'h64;        memory[10456] <=  8'h6d;        memory[10457] <=  8'h73;        memory[10458] <=  8'h6c;        memory[10459] <=  8'h63;        memory[10460] <=  8'h78;        memory[10461] <=  8'h6b;        memory[10462] <=  8'h20;        memory[10463] <=  8'h6f;        memory[10464] <=  8'h78;        memory[10465] <=  8'h63;        memory[10466] <=  8'h76;        memory[10467] <=  8'h6a;        memory[10468] <=  8'h64;        memory[10469] <=  8'h62;        memory[10470] <=  8'h71;        memory[10471] <=  8'h77;        memory[10472] <=  8'h65;        memory[10473] <=  8'h6e;        memory[10474] <=  8'h6d;        memory[10475] <=  8'h64;        memory[10476] <=  8'h6c;        memory[10477] <=  8'h73;        memory[10478] <=  8'h2c;        memory[10479] <=  8'h76;        memory[10480] <=  8'h63;        memory[10481] <=  8'h78;        memory[10482] <=  8'h20;        memory[10483] <=  8'h63;        memory[10484] <=  8'h6f;        memory[10485] <=  8'h69;        memory[10486] <=  8'h76;        memory[10487] <=  8'h68;        memory[10488] <=  8'h73;        memory[10489] <=  8'h64;        memory[10490] <=  8'h62;        memory[10491] <=  8'h71;        memory[10492] <=  8'h77;        memory[10493] <=  8'h65;        memory[10494] <=  8'h6e;        memory[10495] <=  8'h64;        memory[10496] <=  8'h6b;        memory[10497] <=  8'h73;        memory[10498] <=  8'h76;        memory[10499] <=  8'h6f;        memory[10500] <=  8'h63;        memory[10501] <=  8'h20;        memory[10502] <=  8'h76;        memory[10503] <=  8'h69;        memory[10504] <=  8'h75;        memory[10505] <=  8'h69;        memory[10506] <=  8'h68;        memory[10507] <=  8'h63;        memory[10508] <=  8'h78;        memory[10509] <=  8'h69;        memory[10510] <=  8'h6f;        memory[10511] <=  8'h76;        memory[10512] <=  8'h73;        memory[10513] <=  8'h64;        memory[10514] <=  8'h61;        memory[10515] <=  8'h64;        memory[10516] <=  8'h6e;        memory[10517] <=  8'h77;        memory[10518] <=  8'h71;        memory[10519] <=  8'h6b;        memory[10520] <=  8'h6c;        memory[10521] <=  8'h73;        memory[10522] <=  8'h76;        memory[10523] <=  8'h6e;        memory[10524] <=  8'h62;        memory[10525] <=  8'h20;        memory[10526] <=  8'h64;        memory[10527] <=  8'h66;        memory[10528] <=  8'h6a;        memory[10529] <=  8'h6b;        memory[10530] <=  8'h71;        memory[10531] <=  8'h64;        memory[10532] <=  8'h77;        memory[10533] <=  8'h65;        memory[10534] <=  8'h6e;        memory[10535] <=  8'h62;        memory[10536] <=  8'h20;        memory[10537] <=  8'h64;        memory[10538] <=  8'h73;        memory[10539] <=  8'h76;        memory[10540] <=  8'h68;        memory[10541] <=  8'h64;        memory[10542] <=  8'h61;        memory[10543] <=  8'h71;        memory[10544] <=  8'h77;        memory[10545] <=  8'h6a;        memory[10546] <=  8'h65;        memory[10547] <=  8'h6e;        memory[10548] <=  8'h64;        memory[10549] <=  8'h20;        memory[10550] <=  8'h61;        memory[10551] <=  8'h63;        memory[10552] <=  8'h62;        memory[10553] <=  8'h68;        memory[10554] <=  8'h64;        memory[10555] <=  8'h61;        memory[10556] <=  8'h77;        memory[10557] <=  8'h71;        memory[10558] <=  8'h6e;        memory[10559] <=  8'h20;        memory[10560] <=  8'h62;        memory[10561] <=  8'h73;        memory[10562] <=  8'h76;        memory[10563] <=  8'h61;        memory[10564] <=  8'h67;        memory[10565] <=  8'h76;        memory[10566] <=  8'h68;        memory[10567] <=  8'h67;        memory[10568] <=  8'h61;        memory[10569] <=  8'h73;        memory[10570] <=  8'h6a;        memory[10571] <=  8'h6b;        memory[10572] <=  8'h63;        memory[10573] <=  8'h78;        memory[10574] <=  8'h76;        memory[10575] <=  8'h6e;        memory[10576] <=  8'h73;        memory[10577] <=  8'h64;        memory[10578] <=  8'h20;        memory[10579] <=  8'h66;        memory[10580] <=  8'h62;        memory[10581] <=  8'h64;        memory[10582] <=  8'h61;        memory[10583] <=  8'h73;        memory[10584] <=  8'h76;        memory[10585] <=  8'h67;        memory[10586] <=  8'h63;        memory[10587] <=  8'h79;        memory[10588] <=  8'h7a;        memory[10589] <=  8'h78;        memory[10590] <=  8'h79;        memory[10591] <=  8'h75;        memory[10592] <=  8'h20;        memory[10593] <=  8'h69;        memory[10594] <=  8'h6a;        memory[10595] <=  8'h64;        memory[10596] <=  8'h66;        memory[10597] <=  8'h6b;        memory[10598] <=  8'h61;        memory[10599] <=  8'h64;        memory[10600] <=  8'h63;        memory[10601] <=  8'h78;        memory[10602] <=  8'h68;        memory[10603] <=  8'h20;        memory[10604] <=  8'h67;        memory[10605] <=  8'h61;        memory[10606] <=  8'h68;        memory[10607] <=  8'h75;        memory[10608] <=  8'h64;        memory[10609] <=  8'h73;        memory[10610] <=  8'h69;        memory[10611] <=  8'h6a;        memory[10612] <=  8'h61;        memory[10613] <=  8'h6b;        memory[10614] <=  8'h63;        memory[10615] <=  8'h62;        memory[10616] <=  8'h61;        memory[10617] <=  8'h72;        memory[10618] <=  8'h73;        memory[10619] <=  8'h68;        memory[10620] <=  8'h64;        memory[10621] <=  8'h66;        memory[10622] <=  8'h67;        memory[10623] <=  8'h73;        memory[10624] <=  8'h68;        memory[10625] <=  8'h64;        memory[10626] <=  8'h66;        memory[10627] <=  8'h68;        memory[10628] <=  8'h64;        memory[10629] <=  8'h6a;        memory[10630] <=  8'h68;        memory[10631] <=  8'h62;        memory[10632] <=  8'h67;        memory[10633] <=  8'h63;        memory[10634] <=  8'h61;        memory[10635] <=  8'h66;        memory[10636] <=  8'h73;        memory[10637] <=  8'h79;        memory[10638] <=  8'h67;        memory[10639] <=  8'h6b;        memory[10640] <=  8'h75;        memory[10641] <=  8'h64;        memory[10642] <=  8'h68;        memory[10643] <=  8'h62;        memory[10644] <=  8'h77;        memory[10645] <=  8'h76;        memory[10646] <=  8'h67;        memory[10647] <=  8'h61;        memory[10648] <=  8'h66;        memory[10649] <=  8'h64;        memory[10650] <=  8'h74;        memory[10651] <=  8'h75;        memory[10652] <=  8'h66;        memory[10653] <=  8'h79;        memory[10654] <=  8'h67;        memory[10655] <=  8'h69;        memory[10656] <=  8'h75;        memory[10657] <=  8'h68;        memory[10658] <=  8'h6c;        memory[10659] <=  8'h6a;        memory[10660] <=  8'h62;        memory[10661] <=  8'h6b;        memory[10662] <=  8'h68;        memory[10663] <=  8'h76;        memory[10664] <=  8'h67;        memory[10665] <=  8'h63;        memory[10666] <=  8'h66;        memory[10667] <=  8'h78;        memory[10668] <=  8'h64;        memory[10669] <=  8'h74;        memory[10670] <=  8'h75;        memory[10671] <=  8'h79;        memory[10672] <=  8'h69;        memory[10673] <=  8'h75;        memory[10674] <=  8'h68;        memory[10675] <=  8'h6c;        memory[10676] <=  8'h6a;        memory[10677] <=  8'h6b;        memory[10678] <=  8'h67;        memory[10679] <=  8'h6a;        memory[10680] <=  8'h63;        memory[10681] <=  8'h66;        memory[10682] <=  8'h68;        memory[10683] <=  8'h64;        memory[10684] <=  8'h67;        memory[10685] <=  8'h72;        memory[10686] <=  8'h79;        memory[10687] <=  8'h74;        memory[10688] <=  8'h66;        memory[10689] <=  8'h75;        memory[10690] <=  8'h79;        memory[10691] <=  8'h69;        memory[10692] <=  8'h68;        memory[10693] <=  8'h6c;        memory[10694] <=  8'h62;        memory[10695] <=  8'h6d;        memory[10696] <=  8'h76;        memory[10697] <=  8'h6e;        memory[10698] <=  8'h63;        memory[10699] <=  8'h66;        memory[10700] <=  8'h68;        memory[10701] <=  8'h64;        memory[10702] <=  8'h74;        memory[10703] <=  8'h75;        memory[10704] <=  8'h67;        memory[10705] <=  8'h79;        memory[10706] <=  8'h69;        memory[10707] <=  8'h68;        memory[10708] <=  8'h75;        memory[10709] <=  8'h6a;        memory[10710] <=  8'h6c;        memory[10711] <=  8'h62;        memory[10712] <=  8'h6d;        memory[10713] <=  8'h76;        memory[10714] <=  8'h6e;        memory[10715] <=  8'h63;        memory[10716] <=  8'h66;        memory[10717] <=  8'h68;        memory[10718] <=  8'h67;        memory[10719] <=  8'h79;        memory[10720] <=  8'h68;        memory[10721] <=  8'h75;        memory[10722] <=  8'h6a;        memory[10723] <=  8'h6e;        memory[10724] <=  8'h2c;        memory[10725] <=  8'h62;        memory[10726] <=  8'h6e;        memory[10727] <=  8'h6d;        memory[10728] <=  8'h76;        memory[10729] <=  8'h6e;        memory[10730] <=  8'h63;        memory[10731] <=  8'h66;        memory[10732] <=  8'h68;        memory[10733] <=  8'h74;        memory[10734] <=  8'h79;        memory[10735] <=  8'h69;        memory[10736] <=  8'h75;        memory[10737] <=  8'h6c;        memory[10738] <=  8'h6a;        memory[10739] <=  8'h62;        memory[10740] <=  8'h6d;        memory[10741] <=  8'h76;        memory[10742] <=  8'h6e;        memory[10743] <=  8'h63;        memory[10744] <=  8'h66;        memory[10745] <=  8'h74;        memory[10746] <=  8'h75;        memory[10747] <=  8'h79;        memory[10748] <=  8'h69;        memory[10749] <=  8'h68;        memory[10750] <=  8'h6b;        memory[10751] <=  8'h62;        memory[10752] <=  8'h76;        memory[10753] <=  8'h63;        memory[10754] <=  8'h66;        memory[10755] <=  8'h67;        memory[10756] <=  8'h74;        memory[10757] <=  8'h75;        memory[10758] <=  8'h79;        memory[10759] <=  8'h69;        memory[10760] <=  8'h75;        memory[10761] <=  8'h68;        memory[10762] <=  8'h6a;        memory[10763] <=  8'h6b;        memory[10764] <=  8'h62;        memory[10765] <=  8'h76;        memory[10766] <=  8'h63;        memory[10767] <=  8'h66;        memory[10768] <=  8'h74;        memory[10769] <=  8'h75;        memory[10770] <=  8'h79;        memory[10771] <=  8'h69;        memory[10772] <=  8'h75;        memory[10773] <=  8'h6a;        memory[10774] <=  8'h6b;        memory[10775] <=  8'h6e;        memory[10776] <=  8'h62;        memory[10777] <=  8'h76;        memory[10778] <=  8'h67;        memory[10779] <=  8'h66;        memory[10780] <=  8'h74;        memory[10781] <=  8'h79;        memory[10782] <=  8'h75;        memory[10783] <=  8'h75;        memory[10784] <=  8'h69;        memory[10785] <=  8'h6a;        memory[10786] <=  8'h6b;        memory[10787] <=  8'h68;        memory[10788] <=  8'h62;        memory[10789] <=  8'h6a;        memory[10790] <=  8'h67;        memory[10791] <=  8'h68;        memory[10792] <=  8'h66;        memory[10793] <=  8'h79;        memory[10794] <=  8'h74;        memory[10795] <=  8'h79;        memory[10796] <=  8'h69;        memory[10797] <=  8'h75;        memory[10798] <=  8'h64;        memory[10799] <=  8'h6a;        memory[10800] <=  8'h6b;        memory[10801] <=  8'h68;        memory[10802] <=  8'h63;        memory[10803] <=  8'h7a;        memory[10804] <=  8'h67;        memory[10805] <=  8'h68;        memory[10806] <=  8'h74;        memory[10807] <=  8'h75;        memory[10808] <=  8'h79;        memory[10809] <=  8'h69;        memory[10810] <=  8'h61;        memory[10811] <=  8'h73;        memory[10812] <=  8'h75;        memory[10813] <=  8'h6a;        memory[10814] <=  8'h6b;        memory[10815] <=  8'h62;        memory[10816] <=  8'h6e;        memory[10817] <=  8'h61;        memory[10818] <=  8'h76;        memory[10819] <=  8'h63;        memory[10820] <=  8'h66;        memory[10821] <=  8'h68;        memory[10822] <=  8'h75;        memory[10823] <=  8'h61;        memory[10824] <=  8'h73;        memory[10825] <=  8'h79;        memory[10826] <=  8'h64;        memory[10827] <=  8'h75;        memory[10828] <=  8'h69;        memory[10829] <=  8'h6a;        memory[10830] <=  8'h61;        memory[10831] <=  8'h6b;        memory[10832] <=  8'h62;        memory[10833] <=  8'h63;        memory[10834] <=  8'h78;        memory[10835] <=  8'h68;        memory[10836] <=  8'h67;        memory[10837] <=  8'h79;        memory[10838] <=  8'h75;        memory[10839] <=  8'h7a;        memory[10840] <=  8'h63;        memory[10841] <=  8'h61;        memory[10842] <=  8'h73;        memory[10843] <=  8'h69;        memory[10844] <=  8'h75;        memory[10845] <=  8'h6f;        memory[10846] <=  8'h69;        memory[10847] <=  8'h6a;        memory[10848] <=  8'h61;        memory[10849] <=  8'h6c;        memory[10850] <=  8'h63;        memory[10851] <=  8'h78;        memory[10852] <=  8'h62;        memory[10853] <=  8'h63;        memory[10854] <=  8'h20;        memory[10855] <=  8'h6e;        memory[10856] <=  8'h76;        memory[10857] <=  8'h63;        memory[10858] <=  8'h61;        memory[10859] <=  8'h64;        memory[10860] <=  8'h73;        memory[10861] <=  8'h67;        memory[10862] <=  8'h79;        memory[10863] <=  8'h68;        memory[10864] <=  8'h75;        memory[10865] <=  8'h61;        memory[10866] <=  8'h6a;        memory[10867] <=  8'h6b;        memory[10868] <=  8'h78;        memory[10869] <=  8'h62;        memory[10870] <=  8'h20;        memory[10871] <=  8'h6e;        memory[10872] <=  8'h76;        memory[10873] <=  8'h63;        memory[10874] <=  8'h61;        memory[10875] <=  8'h73;        memory[10876] <=  8'h67;        memory[10877] <=  8'h68;        memory[10878] <=  8'h75;        memory[10879] <=  8'h6a;        memory[10880] <=  8'h6c;        memory[10881] <=  8'h6b;        memory[10882] <=  8'h63;        memory[10883] <=  8'h78;        memory[10884] <=  8'h20;        memory[10885] <=  8'h6a;        memory[10886] <=  8'h6b;        memory[10887] <=  8'h68;        memory[10888] <=  8'h61;        memory[10889] <=  8'h73;        memory[10890] <=  8'h76;        memory[10891] <=  8'h64;        memory[10892] <=  8'h6e;        memory[10893] <=  8'h20;        memory[10894] <=  8'h62;        memory[10895] <=  8'h6e;        memory[10896] <=  8'h6d;        memory[10897] <=  8'h6b;        memory[10898] <=  8'h77;        memory[10899] <=  8'h64;        memory[10900] <=  8'h6f;        memory[10901] <=  8'h77;        memory[10902] <=  8'h69;        memory[10903] <=  8'h6f;        memory[10904] <=  8'h75;        memory[10905] <=  8'h69;        memory[10906] <=  8'h68;        memory[10907] <=  8'h62;        memory[10908] <=  8'h6e;        memory[10909] <=  8'h6b;        memory[10910] <=  8'h77;        memory[10911] <=  8'h69;        memory[10912] <=  8'h6f;        memory[10913] <=  8'h75;        memory[10914] <=  8'h71;        memory[10915] <=  8'h69;        memory[10916] <=  8'h79;        memory[10917] <=  8'h67;        memory[10918] <=  8'h6a;        memory[10919] <=  8'h64;        memory[10920] <=  8'h61;        memory[10921] <=  8'h76;        memory[10922] <=  8'h62;        memory[10923] <=  8'h6e;        memory[10924] <=  8'h6b;        memory[10925] <=  8'h6f;        memory[10926] <=  8'h70;        memory[10927] <=  8'h64;        memory[10928] <=  8'h76;        memory[10929] <=  8'h69;        memory[10930] <=  8'h6f;        memory[10931] <=  8'h75;        memory[10932] <=  8'h69;        memory[10933] <=  8'h48;        memory[10934] <=  8'h42;        memory[10935] <=  8'h6b;        memory[10936] <=  8'h64;        memory[10937] <=  8'h6e;        memory[10938] <=  8'h6c;        memory[10939] <=  8'h71;        memory[10940] <=  8'h6b;        memory[10941] <=  8'h6d;        memory[10942] <=  8'h6a;        memory[10943] <=  8'h70;        memory[10944] <=  8'h69;        memory[10945] <=  8'h6f;        memory[10946] <=  8'h68;        memory[10947] <=  8'h65;        memory[10948] <=  8'h66;        memory[10949] <=  8'h75;        memory[10950] <=  8'h67;        memory[10951] <=  8'h69;        memory[10952] <=  8'h73;        memory[10953] <=  8'h61;        memory[10954] <=  8'h62;        memory[10955] <=  8'h64;        memory[10956] <=  8'h6b;        memory[10957] <=  8'h6a;        memory[10958] <=  8'h6b;        memory[10959] <=  8'h6c;        memory[10960] <=  8'h6a;        memory[10961] <=  8'h69;        memory[10962] <=  8'h73;        memory[10963] <=  8'h6f;        memory[10964] <=  8'h71;        memory[10965] <=  8'h68;        memory[10966] <=  8'h77;        memory[10967] <=  8'h67;        memory[10968] <=  8'h69;        memory[10969] <=  8'h79;        memory[10970] <=  8'h6a;        memory[10971] <=  8'h64;        memory[10972] <=  8'h76;        memory[10973] <=  8'h62;        memory[10974] <=  8'h6e;        memory[10975] <=  8'h61;        memory[10976] <=  8'h73;        memory[10977] <=  8'h66;        memory[10978] <=  8'h6c;        memory[10979] <=  8'h6b;        memory[10980] <=  8'h64;        memory[10981] <=  8'h6a;        memory[10982] <=  8'h68;        memory[10983] <=  8'h63;        memory[10984] <=  8'h67;        memory[10985] <=  8'h6a;        memory[10986] <=  8'h76;        memory[10987] <=  8'h73;        memory[10988] <=  8'h64;        memory[10989] <=  8'h62;        memory[10990] <=  8'h62;        memory[10991] <=  8'h61;        memory[10992] <=  8'h72;        memory[10993] <=  8'h62;        memory[10994] <=  8'h62;        memory[10995] <=  8'h73;        memory[10996] <=  8'h62;        memory[10997] <=  8'h67;        memory[10998] <=  8'h73;        memory[10999] <=  8'h66;        memory[11000] <=  8'h67;        memory[11001] <=  8'h61;        memory[11002] <=  8'h68;        memory[11003] <=  8'h66;        memory[11004] <=  8'h73;        memory[11005] <=  8'h68;        memory[11006] <=  8'h61;        memory[11007] <=  8'h66;        memory[11008] <=  8'h73;        memory[11009] <=  8'h66;        memory[11010] <=  8'h68;        memory[11011] <=  8'h61;        memory[11012] <=  8'h69;        memory[11013] <=  8'h64;        memory[11014] <=  8'h75;        memory[11015] <=  8'h67;        memory[11016] <=  8'h64;        memory[11017] <=  8'h77;        memory[11018] <=  8'h62;        memory[11019] <=  8'h61;        memory[11020] <=  8'h62;        memory[11021] <=  8'h72;        memory[11022] <=  8'h62;        memory[11023] <=  8'h61;        memory[11024] <=  8'h62;        memory[11025] <=  8'h62;        memory[11026] <=  8'h74;        memory[11027] <=  8'h62;        memory[11028] <=  8'h62;        memory[11029] <=  8'h62;        memory[11030] <=  8'h62;        memory[11031] <=  8'h62;        memory[11032] <=  8'h62;        memory[11033] <=  8'h62;        memory[11034] <=  8'h62;        memory[11035] <=  8'h61;        memory[11036] <=  8'h62;        memory[11037] <=  8'h62;        memory[11038] <=  8'h72;        memory[11039] <=  8'h74;        memory[11040] <=  8'h62;        memory[11041] <=  8'h62;        memory[11042] <=  8'h61;        memory[11043] <=  8'h62;        memory[11044] <=  8'h72;        memory[11045] <=  8'h62;        memory[11046] <=  8'h74;        memory[11047] <=  8'h62;        memory[11048] <=  8'h62;        memory[11049] <=  8'h62;        memory[11050] <=  8'h63;        memory[11051] <=  8'h61;        memory[11052] <=  8'h72;        memory[11053] <=  8'h74;        memory[11054] <=  8'h73;        memory[11055] <=  8'h62;        memory[11056] <=  8'h61;        memory[11057] <=  8'h72;        memory[11058] <=  8'h74;        memory[11059] <=  8'h74;        memory[11060] <=  8'h62;        memory[11061] <=  8'h61;        memory[11062] <=  8'h72;        memory[11063] <=  8'h74;        memory[11064] <=  8'h78;        memory[11065] <=  8'h61;        memory[11066] <=  8'h74;        memory[11067] <=  8'h6b;        memory[11068] <=  8'h73;        memory[11069] <=  8'h68;        memory[11070] <=  8'h63;        memory[11071] <=  8'h66;        memory[11072] <=  8'h69;        memory[11073] <=  8'h77;        memory[11074] <=  8'h68;        memory[11075] <=  8'h61;        memory[11076] <=  8'h74;        memory[11077] <=  8'h61;        memory[11078] <=  8'h6e;        memory[11079] <=  8'h61;        memory[11080] <=  8'h62;        memory[11081] <=  8'h61;        memory[11082] <=  8'h63;        memory[11083] <=  8'h61;        memory[11084] <=  8'h74;        memory[11085] <=  8'h61;        memory[11086] <=  8'h62;        memory[11087] <=  8'h61;        memory[11088] <=  8'h72;        memory[11089] <=  8'h63;        memory[11090] <=  8'h61;        memory[11091] <=  8'h68;        memory[11092] <=  8'h64;        memory[11093] <=  8'h75;        memory[11094] <=  8'h63;        memory[11095] <=  8'h74;        memory[11096] <=  8'h61;        memory[11097] <=  8'h64;        memory[11098] <=  8'h61;        memory[11099] <=  8'h61;        memory[11100] <=  8'h63;        memory[11101] <=  8'h61;        memory[11102] <=  8'h72;        memory[11103] <=  8'h63;        memory[11104] <=  8'h74;        memory[11105] <=  8'h72;        memory[11106] <=  8'h63;        memory[11107] <=  8'h61;        memory[11108] <=  8'h74;        memory[11109] <=  8'h72;        memory[11110] <=  8'h63;        memory[11111] <=  8'h61;        memory[11112] <=  8'h74;        memory[11113] <=  8'h63;        memory[11114] <=  8'h62;        memory[11115] <=  8'h61;        memory[11116] <=  8'h74;        memory[11117] <=  8'h62;        memory[11118] <=  8'h72;        memory[11119] <=  8'h63;        memory[11120] <=  8'h61;        memory[11121] <=  8'h74;        memory[11122] <=  8'h72;        memory[11123] <=  8'h6e;        memory[11124] <=  8'h62;        memory[11125] <=  8'h61;        memory[11126] <=  8'h63;        memory[11127] <=  8'h61;        memory[11128] <=  8'h74;        memory[11129] <=  8'h79;        memory[11130] <=  8'h73;        memory[11131] <=  8'h6e;        memory[11132] <=  8'h63;        memory[11133] <=  8'h74;        memory[11134] <=  8'h61;        memory[11135] <=  8'h6e;        memory[11136] <=  8'h62;        memory[11137] <=  8'h61;        memory[11138] <=  8'h63;        memory[11139] <=  8'h72;        memory[11140] <=  8'h6e;        memory[11141] <=  8'h74;        memory[11142] <=  8'h61;        memory[11143] <=  8'h62;        memory[11144] <=  8'h74;        memory[11145] <=  8'h6e;        memory[11146] <=  8'h61;        memory[11147] <=  8'h72;        memory[11148] <=  8'h62;        memory[11149] <=  8'h78;        memory[11150] <=  8'h74;        memory[11151] <=  8'h61;        memory[11152] <=  8'h72;        memory[11153] <=  8'h62;        memory[11154] <=  8'h61;        memory[11155] <=  8'h72;        memory[11156] <=  8'h74;        memory[11157] <=  8'h74;        memory[11158] <=  8'h62;        memory[11159] <=  8'h61;        memory[11160] <=  8'h72;        memory[11161] <=  8'h74;        memory[11162] <=  8'h78;        memory[11163] <=  8'h61;        memory[11164] <=  8'h74;        memory[11165] <=  8'h6b;        memory[11166] <=  8'h73;        memory[11167] <=  8'h68;        memory[11168] <=  8'h63;        memory[11169] <=  8'h66;        memory[11170] <=  8'h69;        memory[11171] <=  8'h77;        memory[11172] <=  8'h68;        memory[11173] <=  8'h61;        memory[11174] <=  8'h74;        memory[11175] <=  8'h61;        memory[11176] <=  8'h6e;        memory[11177] <=  8'h61;        memory[11178] <=  8'h62;        memory[11179] <=  8'h61;        memory[11180] <=  8'h63;        memory[11181] <=  8'h61;        memory[11182] <=  8'h74;        memory[11183] <=  8'h61;        memory[11184] <=  8'h62;        memory[11185] <=  8'h61;        memory[11186] <=  8'h72;        memory[11187] <=  8'h63;        memory[11188] <=  8'h61;        memory[11189] <=  8'h68;        memory[11190] <=  8'h64;        memory[11191] <=  8'h75;        memory[11192] <=  8'h63;        memory[11193] <=  8'h74;        memory[11194] <=  8'h61;        memory[11195] <=  8'h64;        memory[11196] <=  8'h61;        memory[11197] <=  8'h61;        memory[11198] <=  8'h63;        memory[11199] <=  8'h61;        memory[11200] <=  8'h72;        memory[11201] <=  8'h63;        memory[11202] <=  8'h74;        memory[11203] <=  8'h72;        memory[11204] <=  8'h63;        memory[11205] <=  8'h61;        memory[11206] <=  8'h74;        memory[11207] <=  8'h72;        memory[11208] <=  8'h63;        memory[11209] <=  8'h61;        memory[11210] <=  8'h74;        memory[11211] <=  8'h63;        memory[11212] <=  8'h62;        memory[11213] <=  8'h61;        memory[11214] <=  8'h74;        memory[11215] <=  8'h62;        memory[11216] <=  8'h72;        memory[11217] <=  8'h63;        memory[11218] <=  8'h61;        memory[11219] <=  8'h74;        memory[11220] <=  8'h72;        memory[11221] <=  8'h6e;        memory[11222] <=  8'h62;        memory[11223] <=  8'h61;        memory[11224] <=  8'h63;        memory[11225] <=  8'h61;        memory[11226] <=  8'h74;        memory[11227] <=  8'h79;        memory[11228] <=  8'h73;        memory[11229] <=  8'h6e;        memory[11230] <=  8'h63;        memory[11231] <=  8'h74;        memory[11232] <=  8'h61;        memory[11233] <=  8'h6e;        memory[11234] <=  8'h62;        memory[11235] <=  8'h61;        memory[11236] <=  8'h63;        memory[11237] <=  8'h72;        memory[11238] <=  8'h6e;        memory[11239] <=  8'h74;        memory[11240] <=  8'h61;        memory[11241] <=  8'h62;        memory[11242] <=  8'h74;        memory[11243] <=  8'h6e;        memory[11244] <=  8'h61;        memory[11245] <=  8'h72;        memory[11246] <=  8'h62;        memory[11247] <=  8'h78;        memory[11248] <=  8'h74;        memory[11249] <=  8'h61;        memory[11250] <=  8'h72;        memory[11251] <=  8'h62;        memory[11252] <=  8'h61;        memory[11253] <=  8'h72;        memory[11254] <=  8'h74;        memory[11255] <=  8'h74;        memory[11256] <=  8'h62;        memory[11257] <=  8'h61;        memory[11258] <=  8'h72;        memory[11259] <=  8'h74;        memory[11260] <=  8'h78;        memory[11261] <=  8'h61;        memory[11262] <=  8'h74;        memory[11263] <=  8'h6b;        memory[11264] <=  8'h73;        memory[11265] <=  8'h68;        memory[11266] <=  8'h63;        memory[11267] <=  8'h66;        memory[11268] <=  8'h69;        memory[11269] <=  8'h77;        memory[11270] <=  8'h68;        memory[11271] <=  8'h61;        memory[11272] <=  8'h74;        memory[11273] <=  8'h61;        memory[11274] <=  8'h6e;        memory[11275] <=  8'h61;        memory[11276] <=  8'h62;        memory[11277] <=  8'h61;        memory[11278] <=  8'h63;        memory[11279] <=  8'h61;        memory[11280] <=  8'h74;        memory[11281] <=  8'h61;        memory[11282] <=  8'h62;        memory[11283] <=  8'h61;        memory[11284] <=  8'h72;        memory[11285] <=  8'h63;        memory[11286] <=  8'h61;        memory[11287] <=  8'h68;        memory[11288] <=  8'h64;        memory[11289] <=  8'h75;        memory[11290] <=  8'h63;        memory[11291] <=  8'h74;        memory[11292] <=  8'h61;        memory[11293] <=  8'h64;        memory[11294] <=  8'h61;        memory[11295] <=  8'h61;        memory[11296] <=  8'h63;        memory[11297] <=  8'h61;        memory[11298] <=  8'h72;        memory[11299] <=  8'h63;        memory[11300] <=  8'h74;        memory[11301] <=  8'h72;        memory[11302] <=  8'h63;        memory[11303] <=  8'h61;        memory[11304] <=  8'h74;        memory[11305] <=  8'h72;        memory[11306] <=  8'h63;        memory[11307] <=  8'h61;        memory[11308] <=  8'h74;        memory[11309] <=  8'h63;        memory[11310] <=  8'h62;        memory[11311] <=  8'h61;        memory[11312] <=  8'h74;        memory[11313] <=  8'h62;        memory[11314] <=  8'h72;        memory[11315] <=  8'h63;        memory[11316] <=  8'h61;        memory[11317] <=  8'h74;        memory[11318] <=  8'h72;        memory[11319] <=  8'h6e;        memory[11320] <=  8'h62;        memory[11321] <=  8'h61;        memory[11322] <=  8'h63;        memory[11323] <=  8'h61;        memory[11324] <=  8'h74;        memory[11325] <=  8'h79;        memory[11326] <=  8'h73;        memory[11327] <=  8'h6e;        memory[11328] <=  8'h63;        memory[11329] <=  8'h74;        memory[11330] <=  8'h61;        memory[11331] <=  8'h6e;        memory[11332] <=  8'h62;        memory[11333] <=  8'h61;        memory[11334] <=  8'h63;        memory[11335] <=  8'h72;        memory[11336] <=  8'h6e;        memory[11337] <=  8'h74;        memory[11338] <=  8'h61;        memory[11339] <=  8'h62;        memory[11340] <=  8'h74;        memory[11341] <=  8'h6e;        memory[11342] <=  8'h61;        memory[11343] <=  8'h72;        memory[11344] <=  8'h62;        memory[11345] <=  8'h78;        memory[11346] <=  8'h74;        memory[11347] <=  8'h61;        memory[11348] <=  8'h72;        memory[11349] <=  8'h5d;        memory[11350] <=  8'h5d;        memory[11351] <=  8'h65;        memory[11352] <=  8'h66;        memory[11353] <=  8'h77;        memory[11354] <=  8'h65;        memory[11355] <=  8'h5d;        memory[11356] <=  8'h65;        memory[11357] <=  8'h67;        memory[11358] <=  8'h73;        memory[11359] <=  8'h67;        memory[11360] <=  8'h66;        memory[11361] <=  8'h62;        memory[11362] <=  8'h61;        memory[11363] <=  8'h72;        memory[11364] <=  8'h74;        memory[11365] <=  8'h74;        memory[11366] <=  8'h62;        memory[11367] <=  8'h61;        memory[11368] <=  8'h72;        memory[11369] <=  8'h74;        memory[11370] <=  8'h78;        memory[11371] <=  8'h61;        memory[11372] <=  8'h74;        memory[11373] <=  8'h6b;        memory[11374] <=  8'h73;        memory[11375] <=  8'h68;        memory[11376] <=  8'h63;        memory[11377] <=  8'h66;        memory[11378] <=  8'h69;        memory[11379] <=  8'h77;        memory[11380] <=  8'h68;        memory[11381] <=  8'h61;        memory[11382] <=  8'h74;        memory[11383] <=  8'h61;        memory[11384] <=  8'h6e;        memory[11385] <=  8'h61;        memory[11386] <=  8'h62;        memory[11387] <=  8'h61;        memory[11388] <=  8'h63;        memory[11389] <=  8'h61;        memory[11390] <=  8'h74;        memory[11391] <=  8'h61;        memory[11392] <=  8'h62;        memory[11393] <=  8'h61;        memory[11394] <=  8'h72;        memory[11395] <=  8'h63;        memory[11396] <=  8'h61;        memory[11397] <=  8'h68;        memory[11398] <=  8'h64;        memory[11399] <=  8'h75;        memory[11400] <=  8'h63;        memory[11401] <=  8'h74;        memory[11402] <=  8'h61;        memory[11403] <=  8'h64;        memory[11404] <=  8'h61;        memory[11405] <=  8'h61;        memory[11406] <=  8'h63;        memory[11407] <=  8'h61;        memory[11408] <=  8'h72;        memory[11409] <=  8'h63;        memory[11410] <=  8'h74;        memory[11411] <=  8'h72;        memory[11412] <=  8'h63;        memory[11413] <=  8'h61;        memory[11414] <=  8'h74;        memory[11415] <=  8'h72;        memory[11416] <=  8'h63;        memory[11417] <=  8'h61;        memory[11418] <=  8'h74;        memory[11419] <=  8'h63;        memory[11420] <=  8'h62;        memory[11421] <=  8'h61;        memory[11422] <=  8'h74;        memory[11423] <=  8'h62;        memory[11424] <=  8'h72;        memory[11425] <=  8'h63;        memory[11426] <=  8'h61;        memory[11427] <=  8'h74;        memory[11428] <=  8'h72;        memory[11429] <=  8'h6e;        memory[11430] <=  8'h62;        memory[11431] <=  8'h61;        memory[11432] <=  8'h63;        memory[11433] <=  8'h61;        memory[11434] <=  8'h74;        memory[11435] <=  8'h79;        memory[11436] <=  8'h73;        memory[11437] <=  8'h6e;        memory[11438] <=  8'h63;        memory[11439] <=  8'h74;        memory[11440] <=  8'h61;        memory[11441] <=  8'h6e;        memory[11442] <=  8'h62;        memory[11443] <=  8'h61;        memory[11444] <=  8'h63;        memory[11445] <=  8'h72;        memory[11446] <=  8'h6e;        memory[11447] <=  8'h74;        memory[11448] <=  8'h61;        memory[11449] <=  8'h62;        memory[11450] <=  8'h74;        memory[11451] <=  8'h6e;        memory[11452] <=  8'h61;        memory[11453] <=  8'h72;        memory[11454] <=  8'h62;        memory[11455] <=  8'h78;        memory[11456] <=  8'h74;        memory[11457] <=  8'h61;        memory[11458] <=  8'h72;        memory[11459] <=  8'h62;        memory[11460] <=  8'h61;        memory[11461] <=  8'h72;        memory[11462] <=  8'h74;        memory[11463] <=  8'h74;        memory[11464] <=  8'h62;        memory[11465] <=  8'h61;        memory[11466] <=  8'h72;        memory[11467] <=  8'h74;        memory[11468] <=  8'h78;        memory[11469] <=  8'h61;        memory[11470] <=  8'h74;        memory[11471] <=  8'h6b;        memory[11472] <=  8'h73;        memory[11473] <=  8'h68;        memory[11474] <=  8'h63;        memory[11475] <=  8'h66;        memory[11476] <=  8'h69;        memory[11477] <=  8'h77;        memory[11478] <=  8'h68;        memory[11479] <=  8'h61;        memory[11480] <=  8'h74;        memory[11481] <=  8'h61;        memory[11482] <=  8'h6e;        memory[11483] <=  8'h61;        memory[11484] <=  8'h62;        memory[11485] <=  8'h61;        memory[11486] <=  8'h63;        memory[11487] <=  8'h61;        memory[11488] <=  8'h74;        memory[11489] <=  8'h61;        memory[11490] <=  8'h62;        memory[11491] <=  8'h61;        memory[11492] <=  8'h72;        memory[11493] <=  8'h63;        memory[11494] <=  8'h61;        memory[11495] <=  8'h68;        memory[11496] <=  8'h64;        memory[11497] <=  8'h75;        memory[11498] <=  8'h63;        memory[11499] <=  8'h74;        memory[11500] <=  8'h61;        memory[11501] <=  8'h64;        memory[11502] <=  8'h61;        memory[11503] <=  8'h61;        memory[11504] <=  8'h63;        memory[11505] <=  8'h61;        memory[11506] <=  8'h72;        memory[11507] <=  8'h63;        memory[11508] <=  8'h74;        memory[11509] <=  8'h72;        memory[11510] <=  8'h63;        memory[11511] <=  8'h61;        memory[11512] <=  8'h74;        memory[11513] <=  8'h72;        memory[11514] <=  8'h63;        memory[11515] <=  8'h61;        memory[11516] <=  8'h74;        memory[11517] <=  8'h63;        memory[11518] <=  8'h62;        memory[11519] <=  8'h61;        memory[11520] <=  8'h74;        memory[11521] <=  8'h62;        memory[11522] <=  8'h72;        memory[11523] <=  8'h63;        memory[11524] <=  8'h61;        memory[11525] <=  8'h74;        memory[11526] <=  8'h72;        memory[11527] <=  8'h6e;        memory[11528] <=  8'h62;        memory[11529] <=  8'h61;        memory[11530] <=  8'h63;        memory[11531] <=  8'h61;        memory[11532] <=  8'h74;        memory[11533] <=  8'h79;        memory[11534] <=  8'h73;        memory[11535] <=  8'h6e;        memory[11536] <=  8'h63;        memory[11537] <=  8'h74;        memory[11538] <=  8'h61;        memory[11539] <=  8'h6e;        memory[11540] <=  8'h62;        memory[11541] <=  8'h61;        memory[11542] <=  8'h63;        memory[11543] <=  8'h72;        memory[11544] <=  8'h6e;        memory[11545] <=  8'h74;        memory[11546] <=  8'h61;        memory[11547] <=  8'h62;        memory[11548] <=  8'h74;        memory[11549] <=  8'h6e;        memory[11550] <=  8'h61;        memory[11551] <=  8'h72;        memory[11552] <=  8'h62;        memory[11553] <=  8'h78;        memory[11554] <=  8'h74;        memory[11555] <=  8'h61;        memory[11556] <=  8'h72;        memory[11557] <=  8'h64;        memory[11558] <=  8'h66;        memory[11559] <=  8'h73;        memory[11560] <=  8'h67;        memory[11561] <=  8'h76;        memory[11562] <=  8'h68;        memory[11563] <=  8'h62;        memory[11564] <=  8'h6b;        memory[11565] <=  8'h6a;        memory[11566] <=  8'h6e;        memory[11567] <=  8'h6d;        memory[11568] <=  8'h62;        memory[11569] <=  8'h76;        memory[11570] <=  8'h78;        memory[11571] <=  8'h63;        memory[11572] <=  8'h73;        memory[11573] <=  8'h66;        memory[11574] <=  8'h72;        memory[11575] <=  8'h74;        memory[11576] <=  8'h79;        memory[11577] <=  8'h75;        memory[11578] <=  8'h6a;        memory[11579] <=  8'h6e;        memory[11580] <=  8'h62;        memory[11581] <=  8'h76;        memory[11582] <=  8'h63;        memory[11583] <=  8'h64;        memory[11584] <=  8'h74;        memory[11585] <=  8'h79;        memory[11586] <=  8'h75;        memory[11587] <=  8'h69;        memory[11588] <=  8'h6b;        memory[11589] <=  8'h6d;        memory[11590] <=  8'h6e;        memory[11591] <=  8'h62;        memory[11592] <=  8'h76;        memory[11593] <=  8'h63;        memory[11594] <=  8'h78;        memory[11595] <=  8'h73;        memory[11596] <=  8'h64;        memory[11597] <=  8'h72;        memory[11598] <=  8'h74;        memory[11599] <=  8'h79;        memory[11600] <=  8'h75;        memory[11601] <=  8'h69;        memory[11602] <=  8'h6b;        memory[11603] <=  8'h6d;        memory[11604] <=  8'h6e;        memory[11605] <=  8'h62;        memory[11606] <=  8'h76;        memory[11607] <=  8'h63;        memory[11608] <=  8'h73;        memory[11609] <=  8'h77;        memory[11610] <=  8'h33;        memory[11611] <=  8'h34;        memory[11612] <=  8'h35;        memory[11613] <=  8'h36;        memory[11614] <=  8'h37;        memory[11615] <=  8'h38;        memory[11616] <=  8'h69;        memory[11617] <=  8'h6b;        memory[11618] <=  8'h6d;        memory[11619] <=  8'h6e;        memory[11620] <=  8'h62;        memory[11621] <=  8'h76;        memory[11622] <=  8'h63;        memory[11623] <=  8'h64;        memory[11624] <=  8'h65;        memory[11625] <=  8'h72;        memory[11626] <=  8'h36;        memory[11627] <=  8'h37;        memory[11628] <=  8'h38;        memory[11629] <=  8'h69;        memory[11630] <=  8'h6f;        memory[11631] <=  8'h6b;        memory[11632] <=  8'h6a;        memory[11633] <=  8'h6e;        memory[11634] <=  8'h62;        memory[11635] <=  8'h76;        memory[11636] <=  8'h63;        memory[11637] <=  8'h64;        memory[11638] <=  8'h72;        memory[11639] <=  8'h74;        memory[11640] <=  8'h79;        memory[11641] <=  8'h75;        memory[11642] <=  8'h73;        memory[11643] <=  8'h6a;        memory[11644] <=  8'h63;        memory[11645] <=  8'h6e;        memory[11646] <=  8'h62;        memory[11647] <=  8'h64;        memory[11648] <=  8'h66;        memory[11649] <=  8'h73;        memory[11650] <=  8'h74;        memory[11651] <=  8'h79;        memory[11652] <=  8'h75;        memory[11653] <=  8'h61;        memory[11654] <=  8'h69;        memory[11655] <=  8'h6b;        memory[11656] <=  8'h78;        memory[11657] <=  8'h6d;        memory[11658] <=  8'h6e;        memory[11659] <=  8'h73;        memory[11660] <=  8'h6a;        memory[11661] <=  8'h6f;        memory[11662] <=  8'h64;        memory[11663] <=  8'h6c;        memory[11664] <=  8'h63;        memory[11665] <=  8'h78;        memory[11666] <=  8'h62;        memory[11667] <=  8'h61;        memory[11668] <=  8'h72;        memory[11669] <=  8'h74;        memory[11670] <=  8'h78;        memory[11671] <=  8'h61;        memory[11672] <=  8'h74;        memory[11673] <=  8'h6b;        memory[11674] <=  8'h73;        memory[11675] <=  8'h68;        memory[11676] <=  8'h63;        memory[11677] <=  8'h66;        memory[11678] <=  8'h69;        memory[11679] <=  8'h77;        memory[11680] <=  8'h68;        memory[11681] <=  8'h61;        memory[11682] <=  8'h74;        memory[11683] <=  8'h61;        memory[11684] <=  8'h6e;        memory[11685] <=  8'h61;        memory[11686] <=  8'h62;        memory[11687] <=  8'h61;        memory[11688] <=  8'h63;        memory[11689] <=  8'h61;        memory[11690] <=  8'h74;        memory[11691] <=  8'h61;        memory[11692] <=  8'h62;        memory[11693] <=  8'h61;        memory[11694] <=  8'h72;        memory[11695] <=  8'h63;        memory[11696] <=  8'h61;        memory[11697] <=  8'h68;        memory[11698] <=  8'h64;        memory[11699] <=  8'h75;        memory[11700] <=  8'h63;        memory[11701] <=  8'h74;        memory[11702] <=  8'h61;        memory[11703] <=  8'h64;        memory[11704] <=  8'h61;        memory[11705] <=  8'h61;        memory[11706] <=  8'h63;        memory[11707] <=  8'h61;        memory[11708] <=  8'h72;        memory[11709] <=  8'h62;        memory[11710] <=  8'h61;        memory[11711] <=  8'h72;        memory[11712] <=  8'h74;        memory[11713] <=  8'h78;        memory[11714] <=  8'h61;        memory[11715] <=  8'h74;        memory[11716] <=  8'h6b;        memory[11717] <=  8'h73;        memory[11718] <=  8'h68;        memory[11719] <=  8'h63;        memory[11720] <=  8'h66;        memory[11721] <=  8'h69;        memory[11722] <=  8'h77;        memory[11723] <=  8'h68;        memory[11724] <=  8'h61;        memory[11725] <=  8'h74;        memory[11726] <=  8'h61;        memory[11727] <=  8'h6e;        memory[11728] <=  8'h61;        memory[11729] <=  8'h62;        memory[11730] <=  8'h61;        memory[11731] <=  8'h63;        memory[11732] <=  8'h61;        memory[11733] <=  8'h74;        memory[11734] <=  8'h61;        memory[11735] <=  8'h62;        memory[11736] <=  8'h61;        memory[11737] <=  8'h72;        memory[11738] <=  8'h63;        memory[11739] <=  8'h61;        memory[11740] <=  8'h68;        memory[11741] <=  8'h64;        memory[11742] <=  8'h75;        memory[11743] <=  8'h63;        memory[11744] <=  8'h74;        memory[11745] <=  8'h61;        memory[11746] <=  8'h64;        memory[11747] <=  8'h61;        memory[11748] <=  8'h61;        memory[11749] <=  8'h63;        memory[11750] <=  8'h61;        memory[11751] <=  8'h72;        memory[11752] <=  8'h62;        memory[11753] <=  8'h61;        memory[11754] <=  8'h72;        memory[11755] <=  8'h74;        memory[11756] <=  8'h78;        memory[11757] <=  8'h61;        memory[11758] <=  8'h74;        memory[11759] <=  8'h6b;        memory[11760] <=  8'h73;        memory[11761] <=  8'h68;        memory[11762] <=  8'h63;        memory[11763] <=  8'h66;        memory[11764] <=  8'h69;        memory[11765] <=  8'h77;        memory[11766] <=  8'h68;        memory[11767] <=  8'h61;        memory[11768] <=  8'h74;        memory[11769] <=  8'h61;        memory[11770] <=  8'h6e;        memory[11771] <=  8'h61;        memory[11772] <=  8'h62;        memory[11773] <=  8'h61;        memory[11774] <=  8'h63;        memory[11775] <=  8'h61;        memory[11776] <=  8'h74;        memory[11777] <=  8'h61;        memory[11778] <=  8'h62;        memory[11779] <=  8'h61;        memory[11780] <=  8'h72;        memory[11781] <=  8'h63;        memory[11782] <=  8'h61;        memory[11783] <=  8'h68;        memory[11784] <=  8'h64;        memory[11785] <=  8'h75;        memory[11786] <=  8'h63;        memory[11787] <=  8'h74;        memory[11788] <=  8'h61;        memory[11789] <=  8'h64;        memory[11790] <=  8'h61;        memory[11791] <=  8'h61;        memory[11792] <=  8'h63;        memory[11793] <=  8'h61;        memory[11794] <=  8'h72;        memory[11795] <=  8'h62;        memory[11796] <=  8'h61;        memory[11797] <=  8'h72;        memory[11798] <=  8'h74;        memory[11799] <=  8'h78;        memory[11800] <=  8'h61;        memory[11801] <=  8'h74;        memory[11802] <=  8'h6b;        memory[11803] <=  8'h73;        memory[11804] <=  8'h68;        memory[11805] <=  8'h63;        memory[11806] <=  8'h66;        memory[11807] <=  8'h69;        memory[11808] <=  8'h77;        memory[11809] <=  8'h68;        memory[11810] <=  8'h61;        memory[11811] <=  8'h74;        memory[11812] <=  8'h61;        memory[11813] <=  8'h6e;        memory[11814] <=  8'h61;        memory[11815] <=  8'h62;        memory[11816] <=  8'h61;        memory[11817] <=  8'h63;        memory[11818] <=  8'h61;        memory[11819] <=  8'h74;        memory[11820] <=  8'h61;        memory[11821] <=  8'h62;        memory[11822] <=  8'h61;        memory[11823] <=  8'h72;        memory[11824] <=  8'h63;        memory[11825] <=  8'h61;        memory[11826] <=  8'h68;        memory[11827] <=  8'h64;        memory[11828] <=  8'h75;        memory[11829] <=  8'h63;        memory[11830] <=  8'h74;        memory[11831] <=  8'h61;        memory[11832] <=  8'h64;        memory[11833] <=  8'h61;        memory[11834] <=  8'h61;        memory[11835] <=  8'h63;        memory[11836] <=  8'h61;        memory[11837] <=  8'h72;        memory[11838] <=  8'h62;        memory[11839] <=  8'h61;        memory[11840] <=  8'h72;        memory[11841] <=  8'h74;        memory[11842] <=  8'h78;        memory[11843] <=  8'h61;        memory[11844] <=  8'h74;        memory[11845] <=  8'h6b;        memory[11846] <=  8'h73;        memory[11847] <=  8'h68;        memory[11848] <=  8'h63;        memory[11849] <=  8'h66;        memory[11850] <=  8'h69;        memory[11851] <=  8'h77;        memory[11852] <=  8'h68;        memory[11853] <=  8'h61;        memory[11854] <=  8'h74;        memory[11855] <=  8'h61;        memory[11856] <=  8'h6e;        memory[11857] <=  8'h61;        memory[11858] <=  8'h62;        memory[11859] <=  8'h61;        memory[11860] <=  8'h63;        memory[11861] <=  8'h61;        memory[11862] <=  8'h74;        memory[11863] <=  8'h61;        memory[11864] <=  8'h62;        memory[11865] <=  8'h61;        memory[11866] <=  8'h72;        memory[11867] <=  8'h63;        memory[11868] <=  8'h61;        memory[11869] <=  8'h68;        memory[11870] <=  8'h64;        memory[11871] <=  8'h75;        memory[11872] <=  8'h63;        memory[11873] <=  8'h74;        memory[11874] <=  8'h61;        memory[11875] <=  8'h64;        memory[11876] <=  8'h61;        memory[11877] <=  8'h61;        memory[11878] <=  8'h63;        memory[11879] <=  8'h61;        memory[11880] <=  8'h72;        memory[11881] <=  8'h62;        memory[11882] <=  8'h61;        memory[11883] <=  8'h72;        memory[11884] <=  8'h74;        memory[11885] <=  8'h78;        memory[11886] <=  8'h61;        memory[11887] <=  8'h74;        memory[11888] <=  8'h6b;        memory[11889] <=  8'h73;        memory[11890] <=  8'h68;        memory[11891] <=  8'h63;        memory[11892] <=  8'h66;        memory[11893] <=  8'h69;        memory[11894] <=  8'h77;        memory[11895] <=  8'h68;        memory[11896] <=  8'h61;        memory[11897] <=  8'h74;        memory[11898] <=  8'h61;        memory[11899] <=  8'h6e;        memory[11900] <=  8'h61;        memory[11901] <=  8'h62;        memory[11902] <=  8'h61;        memory[11903] <=  8'h63;        memory[11904] <=  8'h61;        memory[11905] <=  8'h74;        memory[11906] <=  8'h61;        memory[11907] <=  8'h62;        memory[11908] <=  8'h61;        memory[11909] <=  8'h72;        memory[11910] <=  8'h63;        memory[11911] <=  8'h61;        memory[11912] <=  8'h68;        memory[11913] <=  8'h64;        memory[11914] <=  8'h75;        memory[11915] <=  8'h63;        memory[11916] <=  8'h74;        memory[11917] <=  8'h61;        memory[11918] <=  8'h64;        memory[11919] <=  8'h61;        memory[11920] <=  8'h61;        memory[11921] <=  8'h63;        memory[11922] <=  8'h61;        memory[11923] <=  8'h72;        memory[11924] <=  8'h62;        memory[11925] <=  8'h61;        memory[11926] <=  8'h72;        memory[11927] <=  8'h74;        memory[11928] <=  8'h78;        memory[11929] <=  8'h61;        memory[11930] <=  8'h74;        memory[11931] <=  8'h6b;        memory[11932] <=  8'h73;        memory[11933] <=  8'h68;        memory[11934] <=  8'h63;        memory[11935] <=  8'h66;        memory[11936] <=  8'h69;        memory[11937] <=  8'h77;        memory[11938] <=  8'h68;        memory[11939] <=  8'h61;        memory[11940] <=  8'h74;        memory[11941] <=  8'h61;        memory[11942] <=  8'h6e;        memory[11943] <=  8'h61;        memory[11944] <=  8'h62;        memory[11945] <=  8'h61;        memory[11946] <=  8'h63;        memory[11947] <=  8'h61;        memory[11948] <=  8'h74;        memory[11949] <=  8'h61;        memory[11950] <=  8'h62;        memory[11951] <=  8'h61;        memory[11952] <=  8'h72;        memory[11953] <=  8'h63;        memory[11954] <=  8'h61;        memory[11955] <=  8'h68;        memory[11956] <=  8'h64;        memory[11957] <=  8'h75;        memory[11958] <=  8'h63;        memory[11959] <=  8'h74;        memory[11960] <=  8'h61;        memory[11961] <=  8'h64;        memory[11962] <=  8'h61;        memory[11963] <=  8'h61;        memory[11964] <=  8'h63;        memory[11965] <=  8'h61;        memory[11966] <=  8'h72;        memory[11967] <=  8'h62;        memory[11968] <=  8'h61;        memory[11969] <=  8'h72;        memory[11970] <=  8'h74;        memory[11971] <=  8'h78;        memory[11972] <=  8'h61;        memory[11973] <=  8'h74;        memory[11974] <=  8'h6b;        memory[11975] <=  8'h73;        memory[11976] <=  8'h68;        memory[11977] <=  8'h63;        memory[11978] <=  8'h66;        memory[11979] <=  8'h69;        memory[11980] <=  8'h77;        memory[11981] <=  8'h68;        memory[11982] <=  8'h61;        memory[11983] <=  8'h74;        memory[11984] <=  8'h61;        memory[11985] <=  8'h6e;        memory[11986] <=  8'h61;        memory[11987] <=  8'h62;        memory[11988] <=  8'h61;        memory[11989] <=  8'h63;        memory[11990] <=  8'h61;        memory[11991] <=  8'h74;        memory[11992] <=  8'h61;        memory[11993] <=  8'h62;        memory[11994] <=  8'h61;        memory[11995] <=  8'h72;        memory[11996] <=  8'h63;        memory[11997] <=  8'h61;        memory[11998] <=  8'h68;        memory[11999] <=  8'h64;        memory[12000] <=  8'h75;        memory[12001] <=  8'h63;        memory[12002] <=  8'h74;        memory[12003] <=  8'h61;        memory[12004] <=  8'h64;        memory[12005] <=  8'h61;        memory[12006] <=  8'h61;        memory[12007] <=  8'h63;        memory[12008] <=  8'h61;        memory[12009] <=  8'h72;        memory[12010] <=  8'h62;        memory[12011] <=  8'h61;        memory[12012] <=  8'h72;        memory[12013] <=  8'h74;        memory[12014] <=  8'h78;        memory[12015] <=  8'h61;        memory[12016] <=  8'h74;        memory[12017] <=  8'h6b;        memory[12018] <=  8'h73;        memory[12019] <=  8'h68;        memory[12020] <=  8'h63;        memory[12021] <=  8'h66;        memory[12022] <=  8'h69;        memory[12023] <=  8'h77;        memory[12024] <=  8'h68;        memory[12025] <=  8'h61;        memory[12026] <=  8'h74;        memory[12027] <=  8'h61;        memory[12028] <=  8'h6e;        memory[12029] <=  8'h61;        memory[12030] <=  8'h62;        memory[12031] <=  8'h61;        memory[12032] <=  8'h63;        memory[12033] <=  8'h61;        memory[12034] <=  8'h74;        memory[12035] <=  8'h61;        memory[12036] <=  8'h62;        memory[12037] <=  8'h61;        memory[12038] <=  8'h72;        memory[12039] <=  8'h63;        memory[12040] <=  8'h61;        memory[12041] <=  8'h68;        memory[12042] <=  8'h64;        memory[12043] <=  8'h75;        memory[12044] <=  8'h63;        memory[12045] <=  8'h74;        memory[12046] <=  8'h61;        memory[12047] <=  8'h64;        memory[12048] <=  8'h61;        memory[12049] <=  8'h61;        memory[12050] <=  8'h63;        memory[12051] <=  8'h61;        memory[12052] <=  8'h72;        memory[12053] <=  8'h62;        memory[12054] <=  8'h61;        memory[12055] <=  8'h72;        memory[12056] <=  8'h74;        memory[12057] <=  8'h74;        memory[12058] <=  8'h62;        memory[12059] <=  8'h61;        memory[12060] <=  8'h72;        memory[12061] <=  8'h74;        memory[12062] <=  8'h78;        memory[12063] <=  8'h61;        memory[12064] <=  8'h74;        memory[12065] <=  8'h6b;        memory[12066] <=  8'h73;        memory[12067] <=  8'h68;        memory[12068] <=  8'h63;        memory[12069] <=  8'h66;        memory[12070] <=  8'h69;        memory[12071] <=  8'h77;        memory[12072] <=  8'h68;        memory[12073] <=  8'h61;        memory[12074] <=  8'h74;        memory[12075] <=  8'h61;        memory[12076] <=  8'h6e;        memory[12077] <=  8'h61;        memory[12078] <=  8'h62;        memory[12079] <=  8'h61;        memory[12080] <=  8'h63;        memory[12081] <=  8'h61;        memory[12082] <=  8'h74;        memory[12083] <=  8'h61;        memory[12084] <=  8'h62;        memory[12085] <=  8'h61;        memory[12086] <=  8'h72;        memory[12087] <=  8'h63;        memory[12088] <=  8'h61;        memory[12089] <=  8'h68;        memory[12090] <=  8'h64;        memory[12091] <=  8'h75;        memory[12092] <=  8'h63;        memory[12093] <=  8'h74;        memory[12094] <=  8'h61;        memory[12095] <=  8'h64;        memory[12096] <=  8'h61;        memory[12097] <=  8'h61;        memory[12098] <=  8'h63;        memory[12099] <=  8'h61;        memory[12100] <=  8'h72;        memory[12101] <=  8'h63;        memory[12102] <=  8'h74;        memory[12103] <=  8'h72;        memory[12104] <=  8'h63;        memory[12105] <=  8'h61;        memory[12106] <=  8'h74;        memory[12107] <=  8'h72;        memory[12108] <=  8'h63;        memory[12109] <=  8'h61;        memory[12110] <=  8'h74;        memory[12111] <=  8'h63;        memory[12112] <=  8'h62;        memory[12113] <=  8'h61;        memory[12114] <=  8'h74;        memory[12115] <=  8'h62;        memory[12116] <=  8'h72;        memory[12117] <=  8'h63;        memory[12118] <=  8'h61;        memory[12119] <=  8'h72;        memory[12120] <=  8'h62;        memory[12121] <=  8'h78;        memory[12122] <=  8'h74;        memory[12123] <=  8'h61;        memory[12124] <=  8'h72;        memory[12125] <=  8'h64;        memory[12126] <=  8'h66;        memory[12127] <=  8'h73;        memory[12128] <=  8'h67;        memory[12129] <=  8'h76;        memory[12130] <=  8'h68;        memory[12131] <=  8'h62;        memory[12132] <=  8'h6b;        memory[12133] <=  8'h6a;        memory[12134] <=  8'h6e;        memory[12135] <=  8'h6d;        memory[12136] <=  8'h62;        memory[12137] <=  8'h76;        memory[12138] <=  8'h78;        memory[12139] <=  8'h63;        memory[12140] <=  8'h73;        memory[12141] <=  8'h66;        memory[12142] <=  8'h72;        memory[12143] <=  8'h74;        memory[12144] <=  8'h79;        memory[12145] <=  8'h75;        memory[12146] <=  8'h6a;        memory[12147] <=  8'h6e;        memory[12148] <=  8'h62;        memory[12149] <=  8'h76;        memory[12150] <=  8'h63;        memory[12151] <=  8'h64;        memory[12152] <=  8'h74;        memory[12153] <=  8'h79;        memory[12154] <=  8'h75;        memory[12155] <=  8'h69;        memory[12156] <=  8'h6b;        memory[12157] <=  8'h6d;        memory[12158] <=  8'h6e;        memory[12159] <=  8'h62;        memory[12160] <=  8'h76;        memory[12161] <=  8'h63;        memory[12162] <=  8'h78;        memory[12163] <=  8'h73;        memory[12164] <=  8'h64;        memory[12165] <=  8'h72;        memory[12166] <=  8'h74;        memory[12167] <=  8'h79;        memory[12168] <=  8'h75;        memory[12169] <=  8'h69;        memory[12170] <=  8'h6b;        memory[12171] <=  8'h6d;        memory[12172] <=  8'h6e;        memory[12173] <=  8'h62;        memory[12174] <=  8'h76;        memory[12175] <=  8'h63;        memory[12176] <=  8'h73;        memory[12177] <=  8'h77;        memory[12178] <=  8'h33;        memory[12179] <=  8'h34;        memory[12180] <=  8'h35;        memory[12181] <=  8'h36;        memory[12182] <=  8'h37;        memory[12183] <=  8'h38;        memory[12184] <=  8'h69;        memory[12185] <=  8'h6b;        memory[12186] <=  8'h6d;        memory[12187] <=  8'h6e;        memory[12188] <=  8'h62;        memory[12189] <=  8'h76;        memory[12190] <=  8'h63;        memory[12191] <=  8'h64;        memory[12192] <=  8'h65;        memory[12193] <=  8'h72;        memory[12194] <=  8'h36;        memory[12195] <=  8'h37;        memory[12196] <=  8'h38;        memory[12197] <=  8'h69;        memory[12198] <=  8'h6f;        memory[12199] <=  8'h6b;        memory[12200] <=  8'h6a;        memory[12201] <=  8'h6e;        memory[12202] <=  8'h62;        memory[12203] <=  8'h76;        memory[12204] <=  8'h63;        memory[12205] <=  8'h64;        memory[12206] <=  8'h72;        memory[12207] <=  8'h74;        memory[12208] <=  8'h79;        memory[12209] <=  8'h75;        memory[12210] <=  8'h73;        memory[12211] <=  8'h6a;        memory[12212] <=  8'h63;        memory[12213] <=  8'h6e;        memory[12214] <=  8'h62;        memory[12215] <=  8'h64;        memory[12216] <=  8'h66;        memory[12217] <=  8'h73;        memory[12218] <=  8'h74;        memory[12219] <=  8'h79;        memory[12220] <=  8'h75;        memory[12221] <=  8'h61;        memory[12222] <=  8'h69;        memory[12223] <=  8'h6b;        memory[12224] <=  8'h78;        memory[12225] <=  8'h6d;        memory[12226] <=  8'h6e;        memory[12227] <=  8'h73;        memory[12228] <=  8'h6a;        memory[12229] <=  8'h6f;        memory[12230] <=  8'h64;        memory[12231] <=  8'h6c;        memory[12232] <=  8'h63;        memory[12233] <=  8'h78;        memory[12234] <=  8'h2c;        memory[12235] <=  8'h6d;        memory[12236] <=  8'h73;        memory[12237] <=  8'h6b;        memory[12238] <=  8'h64;        memory[12239] <=  8'h6c;        memory[12240] <=  8'h70;        memory[12241] <=  8'h5b;        memory[12242] <=  8'h3b;        memory[12243] <=  8'h73;        memory[12244] <=  8'h6c;        memory[12245] <=  8'h64;        memory[12246] <=  8'h70;        memory[12247] <=  8'h76;        memory[12248] <=  8'h63;        memory[12249] <=  8'h5b;        memory[12250] <=  8'h78;        memory[12251] <=  8'h76;        memory[12252] <=  8'h63;        memory[12253] <=  8'h5b;        memory[12254] <=  8'h78;        memory[12255] <=  8'h70;        memory[12256] <=  8'h6f;        memory[12257] <=  8'h20;        memory[12258] <=  8'h62;        memory[12259] <=  8'h61;        memory[12260] <=  8'h72;        memory[12261] <=  8'h74;        memory[12262] <=  8'h74;        memory[12263] <=  8'h62;        memory[12264] <=  8'h61;        memory[12265] <=  8'h72;        memory[12266] <=  8'h74;        memory[12267] <=  8'h78;        memory[12268] <=  8'h61;        memory[12269] <=  8'h74;        memory[12270] <=  8'h6b;        memory[12271] <=  8'h73;        memory[12272] <=  8'h68;        memory[12273] <=  8'h63;        memory[12274] <=  8'h66;        memory[12275] <=  8'h69;        memory[12276] <=  8'h77;        memory[12277] <=  8'h68;        memory[12278] <=  8'h61;        memory[12279] <=  8'h69;        memory[12280] <=  8'h6a;        memory[12281] <=  8'h78;        memory[12282] <=  8'h5d;        memory[12283] <=  8'h65;        memory[12284] <=  8'h6b;        memory[12285] <=  8'h6f;        memory[12286] <=  8'h39;        memory[12287] <=  8'h64;        memory[12288] <=  8'h75;        memory[12289] <=  8'h38;        memory[12290] <=  8'h79;        memory[12291] <=  8'h20;        memory[12292] <=  8'h37;        memory[12293] <=  8'h63;        memory[12294] <=  8'h67;        memory[12295] <=  8'h78;        memory[12296] <=  8'h63;        memory[12297] <=  8'h75;        memory[12298] <=  8'h68;        memory[12299] <=  8'h69;        memory[12300] <=  8'h6a;        memory[12301] <=  8'h77;        memory[12302] <=  8'h69;        memory[12303] <=  8'h64;        memory[12304] <=  8'h66;        memory[12305] <=  8'h68;        memory[12306] <=  8'h75;        memory[12307] <=  8'h76;        memory[12308] <=  8'h64;        memory[12309] <=  8'h62;        memory[12310] <=  8'h66;        memory[12311] <=  8'h6a;        memory[12312] <=  8'h6e;        memory[12313] <=  8'h6b;        memory[12314] <=  8'h6a;        memory[12315] <=  8'h65;        memory[12316] <=  8'h38;        memory[12317] <=  8'h66;        memory[12318] <=  8'h37;        memory[12319] <=  8'h67;        memory[12320] <=  8'h79;        memory[12321] <=  8'h76;        memory[12322] <=  8'h63;        memory[12323] <=  8'h68;        memory[12324] <=  8'h69;        memory[12325] <=  8'h6a;        memory[12326] <=  8'h33;        memory[12327] <=  8'h65;        memory[12328] <=  8'h67;        memory[12329] <=  8'h79;        memory[12330] <=  8'h72;        memory[12331] <=  8'h64;        memory[12332] <=  8'h62;        memory[12333] <=  8'h6e;        memory[12334] <=  8'h63;        memory[12335] <=  8'h7a;        memory[12336] <=  8'h6a;        memory[12337] <=  8'h6f;        memory[12338] <=  8'h66;        memory[12339] <=  8'h78;        memory[12340] <=  8'h6a;        memory[12341] <=  8'h69;        memory[12342] <=  8'h63;        memory[12343] <=  8'h68;        memory[12344] <=  8'h62;        memory[12345] <=  8'h6e;        memory[12346] <=  8'h6d;        memory[12347] <=  8'h63;        memory[12348] <=  8'h73;        memory[12349] <=  8'h6c;        memory[12350] <=  8'h6b;        memory[12351] <=  8'h6a;        memory[12352] <=  8'h69;        memory[12353] <=  8'h68;        memory[12354] <=  8'h76;        memory[12355] <=  8'h75;        memory[12356] <=  8'h69;        memory[12357] <=  8'h64;        memory[12358] <=  8'h68;        memory[12359] <=  8'h75;        memory[12360] <=  8'h67;        memory[12361] <=  8'h79;        memory[12362] <=  8'h62;        memory[12363] <=  8'h68;        memory[12364] <=  8'h65;        memory[12365] <=  8'h6a;        memory[12366] <=  8'h72;        memory[12367] <=  8'h6b;        memory[12368] <=  8'h6a;        memory[12369] <=  8'h6f;        memory[12370] <=  8'h64;        memory[12371] <=  8'h67;        memory[12372] <=  8'h69;        memory[12373] <=  8'h75;        memory[12374] <=  8'h69;        memory[12375] <=  8'h67;        memory[12376] <=  8'h76;        memory[12377] <=  8'h79;        memory[12378] <=  8'h75;        memory[12379] <=  8'h67;        memory[12380] <=  8'h78;        memory[12381] <=  8'h68;        memory[12382] <=  8'h63;        memory[12383] <=  8'h20;        memory[12384] <=  8'h20;        memory[12385] <=  8'h20;        memory[12386] <=  8'h78;        memory[12387] <=  8'h76;        memory[12388] <=  8'h20;        memory[12389] <=  8'h63;        memory[12390] <=  8'h78;        memory[12391] <=  8'h67;        memory[12392] <=  8'h79;        memory[12393] <=  8'h63;        memory[12394] <=  8'h75;        memory[12395] <=  8'h68;        memory[12396] <=  8'h6a;        memory[12397] <=  8'h6b;        memory[12398] <=  8'h61;        memory[12399] <=  8'h6c;        memory[12400] <=  8'h78;        memory[12401] <=  8'h76;        memory[12402] <=  8'h70;        memory[12403] <=  8'h6f;        memory[12404] <=  8'h69;        memory[12405] <=  8'h6a;        memory[12406] <=  8'h69;        memory[12407] <=  8'h68;        memory[12408] <=  8'h6a;        memory[12409] <=  8'h62;        memory[12410] <=  8'h77;        memory[12411] <=  8'h65;        memory[12412] <=  8'h6e;        memory[12413] <=  8'h61;        memory[12414] <=  8'h66;        memory[12415] <=  8'h6d;        memory[12416] <=  8'h64;        memory[12417] <=  8'h6b;        memory[12418] <=  8'h6d;        memory[12419] <=  8'h76;        memory[12420] <=  8'h6c;        memory[12421] <=  8'h63;        memory[12422] <=  8'h6f;        memory[12423] <=  8'h64;        memory[12424] <=  8'h69;        memory[12425] <=  8'h75;        memory[12426] <=  8'h68;        memory[12427] <=  8'h73;        memory[12428] <=  8'h66;        memory[12429] <=  8'h65;        memory[12430] <=  8'h62;        memory[12431] <=  8'h6e;        memory[12432] <=  8'h64;        memory[12433] <=  8'h73;        memory[12434] <=  8'h63;        memory[12435] <=  8'h6b;        memory[12436] <=  8'h20;        memory[12437] <=  8'h78;        memory[12438] <=  8'h6a;        memory[12439] <=  8'h78;        memory[12440] <=  8'h63;        memory[12441] <=  8'h73;        memory[12442] <=  8'h64;        memory[12443] <=  8'h66;        memory[12444] <=  8'h6b;        memory[12445] <=  8'h64;        memory[12446] <=  8'h6e;        memory[12447] <=  8'h6d;        memory[12448] <=  8'h64;        memory[12449] <=  8'h73;        memory[12450] <=  8'h63;        memory[12451] <=  8'h6b;        memory[12452] <=  8'h78;        memory[12453] <=  8'h6c;        memory[12454] <=  8'h6f;        memory[12455] <=  8'h66;        memory[12456] <=  8'h6a;        memory[12457] <=  8'h69;        memory[12458] <=  8'h61;        memory[12459] <=  8'h62;        memory[12460] <=  8'h6e;        memory[12461] <=  8'h20;        memory[12462] <=  8'h78;        memory[12463] <=  8'h6b;        memory[12464] <=  8'h6d;        memory[12465] <=  8'h20;        memory[12466] <=  8'h6f;        memory[12467] <=  8'h63;        memory[12468] <=  8'h76;        memory[12469] <=  8'h73;        memory[12470] <=  8'h64;        memory[12471] <=  8'h69;        memory[12472] <=  8'h66;        memory[12473] <=  8'h68;        memory[12474] <=  8'h65;        memory[12475] <=  8'h71;        memory[12476] <=  8'h6a;        memory[12477] <=  8'h77;        memory[12478] <=  8'h62;        memory[12479] <=  8'h65;        memory[12480] <=  8'h6e;        memory[12481] <=  8'h20;        memory[12482] <=  8'h6d;        memory[12483] <=  8'h64;        memory[12484] <=  8'h73;        memory[12485] <=  8'h6c;        memory[12486] <=  8'h76;        memory[12487] <=  8'h6b;        memory[12488] <=  8'h63;        memory[12489] <=  8'h78;        memory[12490] <=  8'h20;        memory[12491] <=  8'h6f;        memory[12492] <=  8'h78;        memory[12493] <=  8'h69;        memory[12494] <=  8'h63;        memory[12495] <=  8'h6a;        memory[12496] <=  8'h76;        memory[12497] <=  8'h64;        memory[12498] <=  8'h66;        memory[12499] <=  8'h65;        memory[12500] <=  8'h71;        memory[12501] <=  8'h6e;        memory[12502] <=  8'h20;        memory[12503] <=  8'h64;        memory[12504] <=  8'h6d;        memory[12505] <=  8'h73;        memory[12506] <=  8'h6c;        memory[12507] <=  8'h63;        memory[12508] <=  8'h78;        memory[12509] <=  8'h6b;        memory[12510] <=  8'h20;        memory[12511] <=  8'h6f;        memory[12512] <=  8'h78;        memory[12513] <=  8'h63;        memory[12514] <=  8'h76;        memory[12515] <=  8'h6a;        memory[12516] <=  8'h64;        memory[12517] <=  8'h62;        memory[12518] <=  8'h71;        memory[12519] <=  8'h77;        memory[12520] <=  8'h65;        memory[12521] <=  8'h6e;        memory[12522] <=  8'h6d;        memory[12523] <=  8'h64;        memory[12524] <=  8'h6c;        memory[12525] <=  8'h73;        memory[12526] <=  8'h2c;        memory[12527] <=  8'h76;        memory[12528] <=  8'h63;        memory[12529] <=  8'h78;        memory[12530] <=  8'h20;        memory[12531] <=  8'h63;        memory[12532] <=  8'h6f;        memory[12533] <=  8'h69;        memory[12534] <=  8'h76;        memory[12535] <=  8'h68;        memory[12536] <=  8'h73;        memory[12537] <=  8'h64;        memory[12538] <=  8'h62;        memory[12539] <=  8'h71;        memory[12540] <=  8'h77;        memory[12541] <=  8'h65;        memory[12542] <=  8'h6e;        memory[12543] <=  8'h64;        memory[12544] <=  8'h6b;        memory[12545] <=  8'h73;        memory[12546] <=  8'h76;        memory[12547] <=  8'h6f;        memory[12548] <=  8'h63;        memory[12549] <=  8'h20;        memory[12550] <=  8'h76;        memory[12551] <=  8'h69;        memory[12552] <=  8'h75;        memory[12553] <=  8'h69;        memory[12554] <=  8'h68;        memory[12555] <=  8'h63;        memory[12556] <=  8'h78;        memory[12557] <=  8'h69;        memory[12558] <=  8'h6f;        memory[12559] <=  8'h76;        memory[12560] <=  8'h73;        memory[12561] <=  8'h64;        memory[12562] <=  8'h61;        memory[12563] <=  8'h64;        memory[12564] <=  8'h6e;        memory[12565] <=  8'h77;        memory[12566] <=  8'h71;        memory[12567] <=  8'h6b;        memory[12568] <=  8'h6c;        memory[12569] <=  8'h73;        memory[12570] <=  8'h76;        memory[12571] <=  8'h6e;        memory[12572] <=  8'h62;        memory[12573] <=  8'h20;        memory[12574] <=  8'h64;        memory[12575] <=  8'h66;        memory[12576] <=  8'h6a;        memory[12577] <=  8'h6b;        memory[12578] <=  8'h71;        memory[12579] <=  8'h64;        memory[12580] <=  8'h77;        memory[12581] <=  8'h65;        memory[12582] <=  8'h6e;        memory[12583] <=  8'h62;        memory[12584] <=  8'h20;        memory[12585] <=  8'h64;        memory[12586] <=  8'h73;        memory[12587] <=  8'h76;        memory[12588] <=  8'h68;        memory[12589] <=  8'h64;        memory[12590] <=  8'h61;        memory[12591] <=  8'h71;        memory[12592] <=  8'h77;        memory[12593] <=  8'h6a;        memory[12594] <=  8'h65;        memory[12595] <=  8'h6e;        memory[12596] <=  8'h64;        memory[12597] <=  8'h20;        memory[12598] <=  8'h61;        memory[12599] <=  8'h63;        memory[12600] <=  8'h62;        memory[12601] <=  8'h68;        memory[12602] <=  8'h64;        memory[12603] <=  8'h61;        memory[12604] <=  8'h77;        memory[12605] <=  8'h71;        memory[12606] <=  8'h6e;        memory[12607] <=  8'h20;        memory[12608] <=  8'h62;        memory[12609] <=  8'h73;        memory[12610] <=  8'h76;        memory[12611] <=  8'h61;        memory[12612] <=  8'h67;        memory[12613] <=  8'h76;        memory[12614] <=  8'h68;        memory[12615] <=  8'h67;        memory[12616] <=  8'h61;        memory[12617] <=  8'h73;        memory[12618] <=  8'h6a;        memory[12619] <=  8'h6b;        memory[12620] <=  8'h63;        memory[12621] <=  8'h78;        memory[12622] <=  8'h76;        memory[12623] <=  8'h6e;        memory[12624] <=  8'h73;        memory[12625] <=  8'h64;        memory[12626] <=  8'h20;        memory[12627] <=  8'h66;        memory[12628] <=  8'h62;        memory[12629] <=  8'h64;        memory[12630] <=  8'h61;        memory[12631] <=  8'h73;        memory[12632] <=  8'h76;        memory[12633] <=  8'h67;        memory[12634] <=  8'h63;        memory[12635] <=  8'h79;        memory[12636] <=  8'h7a;        memory[12637] <=  8'h78;        memory[12638] <=  8'h79;        memory[12639] <=  8'h75;        memory[12640] <=  8'h20;        memory[12641] <=  8'h69;        memory[12642] <=  8'h6a;        memory[12643] <=  8'h64;        memory[12644] <=  8'h66;        memory[12645] <=  8'h6b;        memory[12646] <=  8'h61;        memory[12647] <=  8'h64;        memory[12648] <=  8'h63;        memory[12649] <=  8'h78;        memory[12650] <=  8'h68;        memory[12651] <=  8'h20;        memory[12652] <=  8'h67;        memory[12653] <=  8'h61;        memory[12654] <=  8'h68;        memory[12655] <=  8'h75;        memory[12656] <=  8'h64;        memory[12657] <=  8'h73;        memory[12658] <=  8'h69;        memory[12659] <=  8'h6a;        memory[12660] <=  8'h61;        memory[12661] <=  8'h6b;        memory[12662] <=  8'h63;        memory[12663] <=  8'h62;        memory[12664] <=  8'h61;        memory[12665] <=  8'h72;        memory[12666] <=  8'h73;        memory[12667] <=  8'h68;        memory[12668] <=  8'h64;        memory[12669] <=  8'h66;        memory[12670] <=  8'h67;        memory[12671] <=  8'h73;        memory[12672] <=  8'h68;        memory[12673] <=  8'h64;        memory[12674] <=  8'h66;        memory[12675] <=  8'h68;        memory[12676] <=  8'h64;        memory[12677] <=  8'h6a;        memory[12678] <=  8'h68;        memory[12679] <=  8'h62;        memory[12680] <=  8'h67;        memory[12681] <=  8'h63;        memory[12682] <=  8'h61;        memory[12683] <=  8'h66;        memory[12684] <=  8'h73;        memory[12685] <=  8'h79;        memory[12686] <=  8'h67;        memory[12687] <=  8'h6b;        memory[12688] <=  8'h75;        memory[12689] <=  8'h64;        memory[12690] <=  8'h68;        memory[12691] <=  8'h62;        memory[12692] <=  8'h77;        memory[12693] <=  8'h76;        memory[12694] <=  8'h67;        memory[12695] <=  8'h61;        memory[12696] <=  8'h66;        memory[12697] <=  8'h64;        memory[12698] <=  8'h74;        memory[12699] <=  8'h75;        memory[12700] <=  8'h66;        memory[12701] <=  8'h79;        memory[12702] <=  8'h67;        memory[12703] <=  8'h69;        memory[12704] <=  8'h75;        memory[12705] <=  8'h68;        memory[12706] <=  8'h6c;        memory[12707] <=  8'h6a;        memory[12708] <=  8'h62;        memory[12709] <=  8'h6b;        memory[12710] <=  8'h68;        memory[12711] <=  8'h76;        memory[12712] <=  8'h67;        memory[12713] <=  8'h63;        memory[12714] <=  8'h66;        memory[12715] <=  8'h78;        memory[12716] <=  8'h64;        memory[12717] <=  8'h74;        memory[12718] <=  8'h75;        memory[12719] <=  8'h79;        memory[12720] <=  8'h69;        memory[12721] <=  8'h75;        memory[12722] <=  8'h68;        memory[12723] <=  8'h6c;        memory[12724] <=  8'h6a;        memory[12725] <=  8'h6b;        memory[12726] <=  8'h67;        memory[12727] <=  8'h6a;        memory[12728] <=  8'h63;        memory[12729] <=  8'h66;        memory[12730] <=  8'h68;        memory[12731] <=  8'h64;        memory[12732] <=  8'h67;        memory[12733] <=  8'h72;        memory[12734] <=  8'h79;        memory[12735] <=  8'h74;        memory[12736] <=  8'h66;        memory[12737] <=  8'h75;        memory[12738] <=  8'h79;        memory[12739] <=  8'h69;        memory[12740] <=  8'h68;        memory[12741] <=  8'h6c;        memory[12742] <=  8'h62;        memory[12743] <=  8'h6d;        memory[12744] <=  8'h76;        memory[12745] <=  8'h6e;        memory[12746] <=  8'h63;        memory[12747] <=  8'h66;        memory[12748] <=  8'h68;        memory[12749] <=  8'h64;        memory[12750] <=  8'h74;        memory[12751] <=  8'h75;        memory[12752] <=  8'h67;        memory[12753] <=  8'h79;        memory[12754] <=  8'h69;        memory[12755] <=  8'h68;        memory[12756] <=  8'h75;        memory[12757] <=  8'h6a;        memory[12758] <=  8'h6c;        memory[12759] <=  8'h62;        memory[12760] <=  8'h6d;        memory[12761] <=  8'h76;        memory[12762] <=  8'h6e;        memory[12763] <=  8'h63;        memory[12764] <=  8'h66;        memory[12765] <=  8'h68;        memory[12766] <=  8'h67;        memory[12767] <=  8'h79;        memory[12768] <=  8'h68;        memory[12769] <=  8'h75;        memory[12770] <=  8'h6a;        memory[12771] <=  8'h6e;        memory[12772] <=  8'h2c;        memory[12773] <=  8'h62;        memory[12774] <=  8'h6e;        memory[12775] <=  8'h6d;        memory[12776] <=  8'h76;        memory[12777] <=  8'h6e;        memory[12778] <=  8'h63;        memory[12779] <=  8'h66;        memory[12780] <=  8'h68;        memory[12781] <=  8'h74;        memory[12782] <=  8'h79;        memory[12783] <=  8'h69;        memory[12784] <=  8'h75;        memory[12785] <=  8'h6c;        memory[12786] <=  8'h6a;        memory[12787] <=  8'h62;        memory[12788] <=  8'h6d;        memory[12789] <=  8'h76;        memory[12790] <=  8'h6e;        memory[12791] <=  8'h63;        memory[12792] <=  8'h66;        memory[12793] <=  8'h74;        memory[12794] <=  8'h75;        memory[12795] <=  8'h79;        memory[12796] <=  8'h69;        memory[12797] <=  8'h68;        memory[12798] <=  8'h6b;        memory[12799] <=  8'h62;        memory[12800] <=  8'h76;        memory[12801] <=  8'h63;        memory[12802] <=  8'h66;        memory[12803] <=  8'h67;        memory[12804] <=  8'h74;        memory[12805] <=  8'h75;        memory[12806] <=  8'h79;        memory[12807] <=  8'h69;        memory[12808] <=  8'h75;        memory[12809] <=  8'h68;        memory[12810] <=  8'h6a;        memory[12811] <=  8'h6b;        memory[12812] <=  8'h62;        memory[12813] <=  8'h76;        memory[12814] <=  8'h63;        memory[12815] <=  8'h66;        memory[12816] <=  8'h74;        memory[12817] <=  8'h75;        memory[12818] <=  8'h79;        memory[12819] <=  8'h69;        memory[12820] <=  8'h75;        memory[12821] <=  8'h6a;        memory[12822] <=  8'h6b;        memory[12823] <=  8'h6e;        memory[12824] <=  8'h62;        memory[12825] <=  8'h76;        memory[12826] <=  8'h67;        memory[12827] <=  8'h66;        memory[12828] <=  8'h74;        memory[12829] <=  8'h79;        memory[12830] <=  8'h75;        memory[12831] <=  8'h75;        memory[12832] <=  8'h69;        memory[12833] <=  8'h6a;        memory[12834] <=  8'h6b;        memory[12835] <=  8'h68;        memory[12836] <=  8'h62;        memory[12837] <=  8'h6a;        memory[12838] <=  8'h67;        memory[12839] <=  8'h68;        memory[12840] <=  8'h66;        memory[12841] <=  8'h79;        memory[12842] <=  8'h74;        memory[12843] <=  8'h79;        memory[12844] <=  8'h69;        memory[12845] <=  8'h75;        memory[12846] <=  8'h64;        memory[12847] <=  8'h6a;        memory[12848] <=  8'h6b;        memory[12849] <=  8'h68;        memory[12850] <=  8'h63;        memory[12851] <=  8'h7a;        memory[12852] <=  8'h67;        memory[12853] <=  8'h68;        memory[12854] <=  8'h74;        memory[12855] <=  8'h75;        memory[12856] <=  8'h79;        memory[12857] <=  8'h69;        memory[12858] <=  8'h61;        memory[12859] <=  8'h73;        memory[12860] <=  8'h75;        memory[12861] <=  8'h6a;        memory[12862] <=  8'h6b;        memory[12863] <=  8'h62;        memory[12864] <=  8'h6e;        memory[12865] <=  8'h61;        memory[12866] <=  8'h76;        memory[12867] <=  8'h63;        memory[12868] <=  8'h66;        memory[12869] <=  8'h68;        memory[12870] <=  8'h75;        memory[12871] <=  8'h61;        memory[12872] <=  8'h73;        memory[12873] <=  8'h79;        memory[12874] <=  8'h64;        memory[12875] <=  8'h75;        memory[12876] <=  8'h69;        memory[12877] <=  8'h6a;        memory[12878] <=  8'h61;        memory[12879] <=  8'h6b;        memory[12880] <=  8'h62;        memory[12881] <=  8'h63;        memory[12882] <=  8'h78;        memory[12883] <=  8'h68;        memory[12884] <=  8'h67;        memory[12885] <=  8'h79;        memory[12886] <=  8'h75;        memory[12887] <=  8'h7a;        memory[12888] <=  8'h63;        memory[12889] <=  8'h61;        memory[12890] <=  8'h73;        memory[12891] <=  8'h69;        memory[12892] <=  8'h75;        memory[12893] <=  8'h6f;        memory[12894] <=  8'h69;        memory[12895] <=  8'h6a;        memory[12896] <=  8'h61;        memory[12897] <=  8'h6c;        memory[12898] <=  8'h63;        memory[12899] <=  8'h78;        memory[12900] <=  8'h62;        memory[12901] <=  8'h63;        memory[12902] <=  8'h20;        memory[12903] <=  8'h6e;        memory[12904] <=  8'h76;        memory[12905] <=  8'h63;        memory[12906] <=  8'h61;        memory[12907] <=  8'h64;        memory[12908] <=  8'h73;        memory[12909] <=  8'h67;        memory[12910] <=  8'h79;        memory[12911] <=  8'h68;        memory[12912] <=  8'h75;        memory[12913] <=  8'h61;        memory[12914] <=  8'h6a;        memory[12915] <=  8'h6b;        memory[12916] <=  8'h78;        memory[12917] <=  8'h62;        memory[12918] <=  8'h20;        memory[12919] <=  8'h6e;        memory[12920] <=  8'h76;        memory[12921] <=  8'h63;        memory[12922] <=  8'h61;        memory[12923] <=  8'h73;        memory[12924] <=  8'h67;        memory[12925] <=  8'h68;        memory[12926] <=  8'h75;        memory[12927] <=  8'h6a;        memory[12928] <=  8'h6c;        memory[12929] <=  8'h6b;        memory[12930] <=  8'h63;        memory[12931] <=  8'h78;        memory[12932] <=  8'h20;        memory[12933] <=  8'h6a;        memory[12934] <=  8'h6b;        memory[12935] <=  8'h68;        memory[12936] <=  8'h61;        memory[12937] <=  8'h73;        memory[12938] <=  8'h76;        memory[12939] <=  8'h64;        memory[12940] <=  8'h6e;        memory[12941] <=  8'h20;        memory[12942] <=  8'h62;        memory[12943] <=  8'h6e;        memory[12944] <=  8'h6d;        memory[12945] <=  8'h6b;        memory[12946] <=  8'h77;        memory[12947] <=  8'h64;        memory[12948] <=  8'h6f;        memory[12949] <=  8'h77;        memory[12950] <=  8'h69;        memory[12951] <=  8'h6f;        memory[12952] <=  8'h75;        memory[12953] <=  8'h69;        memory[12954] <=  8'h68;        memory[12955] <=  8'h62;        memory[12956] <=  8'h6e;        memory[12957] <=  8'h6b;        memory[12958] <=  8'h77;        memory[12959] <=  8'h69;        memory[12960] <=  8'h6f;        memory[12961] <=  8'h75;        memory[12962] <=  8'h71;        memory[12963] <=  8'h69;        memory[12964] <=  8'h79;        memory[12965] <=  8'h67;        memory[12966] <=  8'h6a;        memory[12967] <=  8'h64;        memory[12968] <=  8'h61;        memory[12969] <=  8'h76;        memory[12970] <=  8'h62;        memory[12971] <=  8'h6e;        memory[12972] <=  8'h6b;        memory[12973] <=  8'h6f;        memory[12974] <=  8'h70;        memory[12975] <=  8'h64;        memory[12976] <=  8'h76;        memory[12977] <=  8'h69;        memory[12978] <=  8'h6f;        memory[12979] <=  8'h75;        memory[12980] <=  8'h69;        memory[12981] <=  8'h48;        memory[12982] <=  8'h42;        memory[12983] <=  8'h6b;        memory[12984] <=  8'h64;        memory[12985] <=  8'h6e;        memory[12986] <=  8'h6c;        memory[12987] <=  8'h71;        memory[12988] <=  8'h6b;        memory[12989] <=  8'h6d;        memory[12990] <=  8'h6a;        memory[12991] <=  8'h70;        memory[12992] <=  8'h69;        memory[12993] <=  8'h6f;        memory[12994] <=  8'h68;        memory[12995] <=  8'h65;        memory[12996] <=  8'h66;        memory[12997] <=  8'h75;        memory[12998] <=  8'h67;        memory[12999] <=  8'h69;        memory[13000] <=  8'h73;        memory[13001] <=  8'h61;        memory[13002] <=  8'h62;        memory[13003] <=  8'h64;        memory[13004] <=  8'h6b;        memory[13005] <=  8'h6a;        memory[13006] <=  8'h6b;        memory[13007] <=  8'h6c;        memory[13008] <=  8'h6a;        memory[13009] <=  8'h69;        memory[13010] <=  8'h73;        memory[13011] <=  8'h6f;        memory[13012] <=  8'h71;        memory[13013] <=  8'h68;        memory[13014] <=  8'h77;        memory[13015] <=  8'h67;        memory[13016] <=  8'h69;        memory[13017] <=  8'h79;        memory[13018] <=  8'h6a;        memory[13019] <=  8'h64;        memory[13020] <=  8'h76;        memory[13021] <=  8'h62;        memory[13022] <=  8'h6e;        memory[13023] <=  8'h61;        memory[13024] <=  8'h73;        memory[13025] <=  8'h66;        memory[13026] <=  8'h6c;        memory[13027] <=  8'h6b;        memory[13028] <=  8'h64;        memory[13029] <=  8'h6a;        memory[13030] <=  8'h68;        memory[13031] <=  8'h63;        memory[13032] <=  8'h67;        memory[13033] <=  8'h6a;        memory[13034] <=  8'h76;        memory[13035] <=  8'h73;        memory[13036] <=  8'h64;        memory[13037] <=  8'h62;        memory[13038] <=  8'h62;        memory[13039] <=  8'h61;        memory[13040] <=  8'h72;        memory[13041] <=  8'h62;        memory[13042] <=  8'h62;        memory[13043] <=  8'h73;        memory[13044] <=  8'h62;        memory[13045] <=  8'h67;        memory[13046] <=  8'h73;        memory[13047] <=  8'h66;        memory[13048] <=  8'h67;        memory[13049] <=  8'h61;        memory[13050] <=  8'h68;        memory[13051] <=  8'h66;        memory[13052] <=  8'h73;        memory[13053] <=  8'h68;        memory[13054] <=  8'h61;        memory[13055] <=  8'h66;        memory[13056] <=  8'h73;        memory[13057] <=  8'h66;        memory[13058] <=  8'h68;        memory[13059] <=  8'h61;        memory[13060] <=  8'h69;        memory[13061] <=  8'h64;        memory[13062] <=  8'h75;        memory[13063] <=  8'h67;        memory[13064] <=  8'h64;        memory[13065] <=  8'h77;        memory[13066] <=  8'h62;        memory[13067] <=  8'h61;        memory[13068] <=  8'h62;        memory[13069] <=  8'h72;        memory[13070] <=  8'h62;        memory[13071] <=  8'h61;        memory[13072] <=  8'h62;        memory[13073] <=  8'h62;        memory[13074] <=  8'h74;        memory[13075] <=  8'h62;        memory[13076] <=  8'h62;        memory[13077] <=  8'h62;        memory[13078] <=  8'h62;        memory[13079] <=  8'h62;        memory[13080] <=  8'h62;        memory[13081] <=  8'h62;        memory[13082] <=  8'h62;        memory[13083] <=  8'h61;        memory[13084] <=  8'h62;        memory[13085] <=  8'h62;        memory[13086] <=  8'h72;        memory[13087] <=  8'h74;        memory[13088] <=  8'h62;        memory[13089] <=  8'h62;        memory[13090] <=  8'h61;        memory[13091] <=  8'h62;        memory[13092] <=  8'h72;        memory[13093] <=  8'h62;        memory[13094] <=  8'h74;        memory[13095] <=  8'h62;        memory[13096] <=  8'h62;        memory[13097] <=  8'h62;        memory[13098] <=  8'h63;        memory[13099] <=  8'h61;        memory[13100] <=  8'h72;        memory[13101] <=  8'h74;        memory[13102] <=  8'h73;        memory[13103] <=  8'h62;        memory[13104] <=  8'h61;        memory[13105] <=  8'h72;        memory[13106] <=  8'h74;        memory[13107] <=  8'h74;        memory[13108] <=  8'h62;        memory[13109] <=  8'h61;        memory[13110] <=  8'h72;        memory[13111] <=  8'h74;        memory[13112] <=  8'h78;        memory[13113] <=  8'h61;        memory[13114] <=  8'h74;        memory[13115] <=  8'h6b;        memory[13116] <=  8'h73;        memory[13117] <=  8'h68;        memory[13118] <=  8'h63;        memory[13119] <=  8'h66;        memory[13120] <=  8'h69;        memory[13121] <=  8'h77;        memory[13122] <=  8'h68;        memory[13123] <=  8'h61;        memory[13124] <=  8'h74;        memory[13125] <=  8'h61;        memory[13126] <=  8'h6e;        memory[13127] <=  8'h61;        memory[13128] <=  8'h62;        memory[13129] <=  8'h61;        memory[13130] <=  8'h63;        memory[13131] <=  8'h61;        memory[13132] <=  8'h74;        memory[13133] <=  8'h61;        memory[13134] <=  8'h62;        memory[13135] <=  8'h61;        memory[13136] <=  8'h72;        memory[13137] <=  8'h63;        memory[13138] <=  8'h61;        memory[13139] <=  8'h68;        memory[13140] <=  8'h64;        memory[13141] <=  8'h75;        memory[13142] <=  8'h63;        memory[13143] <=  8'h74;        memory[13144] <=  8'h61;        memory[13145] <=  8'h64;        memory[13146] <=  8'h61;        memory[13147] <=  8'h61;        memory[13148] <=  8'h63;        memory[13149] <=  8'h61;        memory[13150] <=  8'h72;        memory[13151] <=  8'h63;        memory[13152] <=  8'h74;        memory[13153] <=  8'h72;        memory[13154] <=  8'h63;        memory[13155] <=  8'h61;        memory[13156] <=  8'h74;        memory[13157] <=  8'h72;        memory[13158] <=  8'h63;        memory[13159] <=  8'h61;        memory[13160] <=  8'h74;        memory[13161] <=  8'h63;        memory[13162] <=  8'h62;        memory[13163] <=  8'h61;        memory[13164] <=  8'h74;        memory[13165] <=  8'h62;        memory[13166] <=  8'h72;        memory[13167] <=  8'h63;        memory[13168] <=  8'h61;        memory[13169] <=  8'h74;        memory[13170] <=  8'h72;        memory[13171] <=  8'h6e;        memory[13172] <=  8'h62;        memory[13173] <=  8'h61;        memory[13174] <=  8'h63;        memory[13175] <=  8'h61;        memory[13176] <=  8'h74;        memory[13177] <=  8'h79;        memory[13178] <=  8'h73;        memory[13179] <=  8'h6e;        memory[13180] <=  8'h63;        memory[13181] <=  8'h74;        memory[13182] <=  8'h61;        memory[13183] <=  8'h6e;        memory[13184] <=  8'h62;        memory[13185] <=  8'h61;        memory[13186] <=  8'h63;        memory[13187] <=  8'h72;        memory[13188] <=  8'h6e;        memory[13189] <=  8'h74;        memory[13190] <=  8'h61;        memory[13191] <=  8'h62;        memory[13192] <=  8'h74;        memory[13193] <=  8'h6e;        memory[13194] <=  8'h61;        memory[13195] <=  8'h72;        memory[13196] <=  8'h62;        memory[13197] <=  8'h78;        memory[13198] <=  8'h74;        memory[13199] <=  8'h61;        memory[13200] <=  8'h72;        memory[13201] <=  8'h62;        memory[13202] <=  8'h61;        memory[13203] <=  8'h72;        memory[13204] <=  8'h74;        memory[13205] <=  8'h74;        memory[13206] <=  8'h62;        memory[13207] <=  8'h61;        memory[13208] <=  8'h72;        memory[13209] <=  8'h74;        memory[13210] <=  8'h78;        memory[13211] <=  8'h61;        memory[13212] <=  8'h74;        memory[13213] <=  8'h6b;        memory[13214] <=  8'h73;        memory[13215] <=  8'h68;        memory[13216] <=  8'h63;        memory[13217] <=  8'h66;        memory[13218] <=  8'h69;        memory[13219] <=  8'h77;        memory[13220] <=  8'h68;        memory[13221] <=  8'h61;        memory[13222] <=  8'h74;        memory[13223] <=  8'h61;        memory[13224] <=  8'h6e;        memory[13225] <=  8'h61;        memory[13226] <=  8'h62;        memory[13227] <=  8'h61;        memory[13228] <=  8'h63;        memory[13229] <=  8'h61;        memory[13230] <=  8'h74;        memory[13231] <=  8'h61;        memory[13232] <=  8'h62;        memory[13233] <=  8'h61;        memory[13234] <=  8'h72;        memory[13235] <=  8'h63;        memory[13236] <=  8'h61;        memory[13237] <=  8'h68;        memory[13238] <=  8'h64;        memory[13239] <=  8'h75;        memory[13240] <=  8'h63;        memory[13241] <=  8'h74;        memory[13242] <=  8'h61;        memory[13243] <=  8'h64;        memory[13244] <=  8'h61;        memory[13245] <=  8'h61;        memory[13246] <=  8'h63;        memory[13247] <=  8'h61;        memory[13248] <=  8'h72;        memory[13249] <=  8'h63;        memory[13250] <=  8'h74;        memory[13251] <=  8'h72;        memory[13252] <=  8'h63;        memory[13253] <=  8'h61;        memory[13254] <=  8'h74;        memory[13255] <=  8'h72;        memory[13256] <=  8'h63;        memory[13257] <=  8'h61;        memory[13258] <=  8'h74;        memory[13259] <=  8'h63;        memory[13260] <=  8'h62;        memory[13261] <=  8'h61;        memory[13262] <=  8'h74;        memory[13263] <=  8'h62;        memory[13264] <=  8'h72;        memory[13265] <=  8'h63;        memory[13266] <=  8'h61;        memory[13267] <=  8'h74;        memory[13268] <=  8'h72;        memory[13269] <=  8'h6e;        memory[13270] <=  8'h62;        memory[13271] <=  8'h61;        memory[13272] <=  8'h63;        memory[13273] <=  8'h61;        memory[13274] <=  8'h74;        memory[13275] <=  8'h79;        memory[13276] <=  8'h73;        memory[13277] <=  8'h6e;        memory[13278] <=  8'h63;        memory[13279] <=  8'h74;        memory[13280] <=  8'h61;        memory[13281] <=  8'h6e;        memory[13282] <=  8'h62;        memory[13283] <=  8'h61;        memory[13284] <=  8'h63;        memory[13285] <=  8'h72;        memory[13286] <=  8'h6e;        memory[13287] <=  8'h74;        memory[13288] <=  8'h61;        memory[13289] <=  8'h62;        memory[13290] <=  8'h74;        memory[13291] <=  8'h6e;        memory[13292] <=  8'h61;        memory[13293] <=  8'h72;        memory[13294] <=  8'h62;        memory[13295] <=  8'h78;        memory[13296] <=  8'h74;        memory[13297] <=  8'h61;        memory[13298] <=  8'h72;        memory[13299] <=  8'h62;        memory[13300] <=  8'h61;        memory[13301] <=  8'h72;        memory[13302] <=  8'h74;        memory[13303] <=  8'h74;        memory[13304] <=  8'h62;        memory[13305] <=  8'h61;        memory[13306] <=  8'h72;        memory[13307] <=  8'h74;        memory[13308] <=  8'h78;        memory[13309] <=  8'h61;        memory[13310] <=  8'h74;        memory[13311] <=  8'h6b;        memory[13312] <=  8'h73;        memory[13313] <=  8'h68;        memory[13314] <=  8'h63;        memory[13315] <=  8'h66;        memory[13316] <=  8'h69;        memory[13317] <=  8'h77;        memory[13318] <=  8'h68;        memory[13319] <=  8'h61;        memory[13320] <=  8'h74;        memory[13321] <=  8'h61;        memory[13322] <=  8'h6e;        memory[13323] <=  8'h61;        memory[13324] <=  8'h62;        memory[13325] <=  8'h61;        memory[13326] <=  8'h63;        memory[13327] <=  8'h61;        memory[13328] <=  8'h74;        memory[13329] <=  8'h61;        memory[13330] <=  8'h62;        memory[13331] <=  8'h61;        memory[13332] <=  8'h72;        memory[13333] <=  8'h63;        memory[13334] <=  8'h61;        memory[13335] <=  8'h68;        memory[13336] <=  8'h64;        memory[13337] <=  8'h75;        memory[13338] <=  8'h63;        memory[13339] <=  8'h74;        memory[13340] <=  8'h61;        memory[13341] <=  8'h64;        memory[13342] <=  8'h61;        memory[13343] <=  8'h61;        memory[13344] <=  8'h63;        memory[13345] <=  8'h61;        memory[13346] <=  8'h72;        memory[13347] <=  8'h63;        memory[13348] <=  8'h74;        memory[13349] <=  8'h72;        memory[13350] <=  8'h63;        memory[13351] <=  8'h61;        memory[13352] <=  8'h74;        memory[13353] <=  8'h72;        memory[13354] <=  8'h63;        memory[13355] <=  8'h61;        memory[13356] <=  8'h74;        memory[13357] <=  8'h63;        memory[13358] <=  8'h62;        memory[13359] <=  8'h61;        memory[13360] <=  8'h74;        memory[13361] <=  8'h62;        memory[13362] <=  8'h72;        memory[13363] <=  8'h63;        memory[13364] <=  8'h61;        memory[13365] <=  8'h74;        memory[13366] <=  8'h72;        memory[13367] <=  8'h6e;        memory[13368] <=  8'h62;        memory[13369] <=  8'h61;        memory[13370] <=  8'h63;        memory[13371] <=  8'h61;        memory[13372] <=  8'h74;        memory[13373] <=  8'h79;        memory[13374] <=  8'h73;        memory[13375] <=  8'h6e;        memory[13376] <=  8'h63;        memory[13377] <=  8'h74;        memory[13378] <=  8'h61;        memory[13379] <=  8'h6e;        memory[13380] <=  8'h62;        memory[13381] <=  8'h61;        memory[13382] <=  8'h63;        memory[13383] <=  8'h72;        memory[13384] <=  8'h6e;        memory[13385] <=  8'h74;        memory[13386] <=  8'h61;        memory[13387] <=  8'h62;        memory[13388] <=  8'h74;        memory[13389] <=  8'h6e;        memory[13390] <=  8'h61;        memory[13391] <=  8'h72;        memory[13392] <=  8'h62;        memory[13393] <=  8'h78;        memory[13394] <=  8'h74;        memory[13395] <=  8'h61;        memory[13396] <=  8'h72;        memory[13397] <=  8'h5d;        memory[13398] <=  8'h5d;        memory[13399] <=  8'h65;        memory[13400] <=  8'h66;        memory[13401] <=  8'h77;        memory[13402] <=  8'h65;        memory[13403] <=  8'h5d;        memory[13404] <=  8'h65;        memory[13405] <=  8'h67;        memory[13406] <=  8'h73;        memory[13407] <=  8'h67;        memory[13408] <=  8'h66;        memory[13409] <=  8'h62;        memory[13410] <=  8'h61;        memory[13411] <=  8'h72;        memory[13412] <=  8'h74;        memory[13413] <=  8'h74;        memory[13414] <=  8'h62;        memory[13415] <=  8'h61;        memory[13416] <=  8'h72;        memory[13417] <=  8'h74;        memory[13418] <=  8'h78;        memory[13419] <=  8'h61;        memory[13420] <=  8'h74;        memory[13421] <=  8'h6b;        memory[13422] <=  8'h73;        memory[13423] <=  8'h68;        memory[13424] <=  8'h63;        memory[13425] <=  8'h66;        memory[13426] <=  8'h69;        memory[13427] <=  8'h77;        memory[13428] <=  8'h68;        memory[13429] <=  8'h61;        memory[13430] <=  8'h74;        memory[13431] <=  8'h61;        memory[13432] <=  8'h6e;        memory[13433] <=  8'h61;        memory[13434] <=  8'h62;        memory[13435] <=  8'h61;        memory[13436] <=  8'h63;        memory[13437] <=  8'h61;        memory[13438] <=  8'h74;        memory[13439] <=  8'h61;        memory[13440] <=  8'h62;        memory[13441] <=  8'h61;        memory[13442] <=  8'h72;        memory[13443] <=  8'h63;        memory[13444] <=  8'h61;        memory[13445] <=  8'h68;        memory[13446] <=  8'h64;        memory[13447] <=  8'h75;        memory[13448] <=  8'h63;        memory[13449] <=  8'h74;        memory[13450] <=  8'h61;        memory[13451] <=  8'h64;        memory[13452] <=  8'h61;        memory[13453] <=  8'h61;        memory[13454] <=  8'h63;        memory[13455] <=  8'h61;        memory[13456] <=  8'h72;        memory[13457] <=  8'h63;        memory[13458] <=  8'h74;        memory[13459] <=  8'h72;        memory[13460] <=  8'h63;        memory[13461] <=  8'h61;        memory[13462] <=  8'h74;        memory[13463] <=  8'h72;        memory[13464] <=  8'h63;        memory[13465] <=  8'h61;        memory[13466] <=  8'h74;        memory[13467] <=  8'h63;        memory[13468] <=  8'h62;        memory[13469] <=  8'h61;        memory[13470] <=  8'h74;        memory[13471] <=  8'h62;        memory[13472] <=  8'h72;        memory[13473] <=  8'h63;        memory[13474] <=  8'h61;        memory[13475] <=  8'h74;        memory[13476] <=  8'h72;        memory[13477] <=  8'h6e;        memory[13478] <=  8'h62;        memory[13479] <=  8'h61;        memory[13480] <=  8'h63;        memory[13481] <=  8'h61;        memory[13482] <=  8'h74;        memory[13483] <=  8'h79;        memory[13484] <=  8'h73;        memory[13485] <=  8'h6e;        memory[13486] <=  8'h63;        memory[13487] <=  8'h74;        memory[13488] <=  8'h61;        memory[13489] <=  8'h6e;        memory[13490] <=  8'h62;        memory[13491] <=  8'h61;        memory[13492] <=  8'h63;        memory[13493] <=  8'h72;        memory[13494] <=  8'h6e;        memory[13495] <=  8'h74;        memory[13496] <=  8'h61;        memory[13497] <=  8'h62;        memory[13498] <=  8'h74;        memory[13499] <=  8'h6e;        memory[13500] <=  8'h61;        memory[13501] <=  8'h72;        memory[13502] <=  8'h62;        memory[13503] <=  8'h78;        memory[13504] <=  8'h74;        memory[13505] <=  8'h61;        memory[13506] <=  8'h72;        memory[13507] <=  8'h62;        memory[13508] <=  8'h61;        memory[13509] <=  8'h72;        memory[13510] <=  8'h74;        memory[13511] <=  8'h74;        memory[13512] <=  8'h62;        memory[13513] <=  8'h61;        memory[13514] <=  8'h72;        memory[13515] <=  8'h74;        memory[13516] <=  8'h78;        memory[13517] <=  8'h61;        memory[13518] <=  8'h74;        memory[13519] <=  8'h6b;        memory[13520] <=  8'h73;        memory[13521] <=  8'h68;        memory[13522] <=  8'h63;        memory[13523] <=  8'h66;        memory[13524] <=  8'h69;        memory[13525] <=  8'h77;        memory[13526] <=  8'h68;        memory[13527] <=  8'h61;        memory[13528] <=  8'h74;        memory[13529] <=  8'h61;        memory[13530] <=  8'h6e;        memory[13531] <=  8'h61;        memory[13532] <=  8'h62;        memory[13533] <=  8'h61;        memory[13534] <=  8'h63;        memory[13535] <=  8'h61;        memory[13536] <=  8'h74;        memory[13537] <=  8'h61;        memory[13538] <=  8'h62;        memory[13539] <=  8'h61;        memory[13540] <=  8'h72;        memory[13541] <=  8'h63;        memory[13542] <=  8'h61;        memory[13543] <=  8'h68;        memory[13544] <=  8'h64;        memory[13545] <=  8'h75;        memory[13546] <=  8'h63;        memory[13547] <=  8'h74;        memory[13548] <=  8'h61;        memory[13549] <=  8'h64;        memory[13550] <=  8'h61;        memory[13551] <=  8'h61;        memory[13552] <=  8'h63;        memory[13553] <=  8'h61;        memory[13554] <=  8'h72;        memory[13555] <=  8'h63;        memory[13556] <=  8'h74;        memory[13557] <=  8'h72;        memory[13558] <=  8'h63;        memory[13559] <=  8'h61;        memory[13560] <=  8'h74;        memory[13561] <=  8'h72;        memory[13562] <=  8'h63;        memory[13563] <=  8'h61;        memory[13564] <=  8'h74;        memory[13565] <=  8'h63;        memory[13566] <=  8'h62;        memory[13567] <=  8'h61;        memory[13568] <=  8'h74;        memory[13569] <=  8'h62;        memory[13570] <=  8'h72;        memory[13571] <=  8'h63;        memory[13572] <=  8'h61;        memory[13573] <=  8'h74;        memory[13574] <=  8'h72;        memory[13575] <=  8'h6e;        memory[13576] <=  8'h62;        memory[13577] <=  8'h61;        memory[13578] <=  8'h63;        memory[13579] <=  8'h61;        memory[13580] <=  8'h74;        memory[13581] <=  8'h79;        memory[13582] <=  8'h73;        memory[13583] <=  8'h6e;        memory[13584] <=  8'h63;        memory[13585] <=  8'h74;        memory[13586] <=  8'h61;        memory[13587] <=  8'h6e;        memory[13588] <=  8'h62;        memory[13589] <=  8'h61;        memory[13590] <=  8'h63;        memory[13591] <=  8'h72;        memory[13592] <=  8'h6e;        memory[13593] <=  8'h74;        memory[13594] <=  8'h61;        memory[13595] <=  8'h62;        memory[13596] <=  8'h74;        memory[13597] <=  8'h6e;        memory[13598] <=  8'h61;        memory[13599] <=  8'h72;        memory[13600] <=  8'h62;        memory[13601] <=  8'h78;        memory[13602] <=  8'h74;        memory[13603] <=  8'h61;        memory[13604] <=  8'h72;        memory[13605] <=  8'h64;        memory[13606] <=  8'h66;        memory[13607] <=  8'h73;        memory[13608] <=  8'h67;        memory[13609] <=  8'h76;        memory[13610] <=  8'h68;        memory[13611] <=  8'h62;        memory[13612] <=  8'h6b;        memory[13613] <=  8'h6a;        memory[13614] <=  8'h6e;        memory[13615] <=  8'h6d;        memory[13616] <=  8'h62;        memory[13617] <=  8'h76;        memory[13618] <=  8'h78;        memory[13619] <=  8'h63;        memory[13620] <=  8'h73;        memory[13621] <=  8'h66;        memory[13622] <=  8'h72;        memory[13623] <=  8'h74;        memory[13624] <=  8'h79;        memory[13625] <=  8'h75;        memory[13626] <=  8'h6a;        memory[13627] <=  8'h6e;        memory[13628] <=  8'h62;        memory[13629] <=  8'h76;        memory[13630] <=  8'h63;        memory[13631] <=  8'h64;        memory[13632] <=  8'h74;        memory[13633] <=  8'h79;        memory[13634] <=  8'h75;        memory[13635] <=  8'h69;        memory[13636] <=  8'h6b;        memory[13637] <=  8'h6d;        memory[13638] <=  8'h6e;        memory[13639] <=  8'h62;        memory[13640] <=  8'h76;        memory[13641] <=  8'h63;        memory[13642] <=  8'h78;        memory[13643] <=  8'h73;        memory[13644] <=  8'h64;        memory[13645] <=  8'h72;        memory[13646] <=  8'h74;        memory[13647] <=  8'h79;        memory[13648] <=  8'h75;        memory[13649] <=  8'h69;        memory[13650] <=  8'h6b;        memory[13651] <=  8'h6d;        memory[13652] <=  8'h6e;        memory[13653] <=  8'h62;        memory[13654] <=  8'h76;        memory[13655] <=  8'h63;        memory[13656] <=  8'h73;        memory[13657] <=  8'h77;        memory[13658] <=  8'h33;        memory[13659] <=  8'h34;        memory[13660] <=  8'h35;        memory[13661] <=  8'h36;        memory[13662] <=  8'h37;        memory[13663] <=  8'h38;        memory[13664] <=  8'h69;        memory[13665] <=  8'h6b;        memory[13666] <=  8'h6d;        memory[13667] <=  8'h6e;        memory[13668] <=  8'h62;        memory[13669] <=  8'h76;        memory[13670] <=  8'h63;        memory[13671] <=  8'h64;        memory[13672] <=  8'h65;        memory[13673] <=  8'h72;        memory[13674] <=  8'h36;        memory[13675] <=  8'h37;        memory[13676] <=  8'h38;        memory[13677] <=  8'h69;        memory[13678] <=  8'h6f;        memory[13679] <=  8'h6b;        memory[13680] <=  8'h6a;        memory[13681] <=  8'h6e;        memory[13682] <=  8'h62;        memory[13683] <=  8'h76;        memory[13684] <=  8'h63;        memory[13685] <=  8'h64;        memory[13686] <=  8'h72;        memory[13687] <=  8'h74;        memory[13688] <=  8'h79;        memory[13689] <=  8'h75;        memory[13690] <=  8'h73;        memory[13691] <=  8'h6a;        memory[13692] <=  8'h63;        memory[13693] <=  8'h6e;        memory[13694] <=  8'h62;        memory[13695] <=  8'h64;        memory[13696] <=  8'h66;        memory[13697] <=  8'h73;        memory[13698] <=  8'h74;        memory[13699] <=  8'h79;        memory[13700] <=  8'h75;        memory[13701] <=  8'h61;        memory[13702] <=  8'h69;        memory[13703] <=  8'h6b;        memory[13704] <=  8'h78;        memory[13705] <=  8'h6d;        memory[13706] <=  8'h6e;        memory[13707] <=  8'h73;        memory[13708] <=  8'h6a;        memory[13709] <=  8'h6f;        memory[13710] <=  8'h64;        memory[13711] <=  8'h6c;        memory[13712] <=  8'h63;        memory[13713] <=  8'h78;        memory[13714] <=  8'h62;        memory[13715] <=  8'h61;        memory[13716] <=  8'h72;        memory[13717] <=  8'h74;        memory[13718] <=  8'h78;        memory[13719] <=  8'h61;        memory[13720] <=  8'h74;        memory[13721] <=  8'h6b;        memory[13722] <=  8'h73;        memory[13723] <=  8'h68;        memory[13724] <=  8'h63;        memory[13725] <=  8'h66;        memory[13726] <=  8'h69;        memory[13727] <=  8'h77;        memory[13728] <=  8'h68;        memory[13729] <=  8'h61;        memory[13730] <=  8'h74;        memory[13731] <=  8'h61;        memory[13732] <=  8'h6e;        memory[13733] <=  8'h61;        memory[13734] <=  8'h62;        memory[13735] <=  8'h61;        memory[13736] <=  8'h63;        memory[13737] <=  8'h61;        memory[13738] <=  8'h74;        memory[13739] <=  8'h61;        memory[13740] <=  8'h62;        memory[13741] <=  8'h61;        memory[13742] <=  8'h72;        memory[13743] <=  8'h63;        memory[13744] <=  8'h61;        memory[13745] <=  8'h68;        memory[13746] <=  8'h64;        memory[13747] <=  8'h75;        memory[13748] <=  8'h63;        memory[13749] <=  8'h74;        memory[13750] <=  8'h61;        memory[13751] <=  8'h64;        memory[13752] <=  8'h61;        memory[13753] <=  8'h61;        memory[13754] <=  8'h63;        memory[13755] <=  8'h61;        memory[13756] <=  8'h72;        memory[13757] <=  8'h62;        memory[13758] <=  8'h61;        memory[13759] <=  8'h72;        memory[13760] <=  8'h74;        memory[13761] <=  8'h78;        memory[13762] <=  8'h61;        memory[13763] <=  8'h74;        memory[13764] <=  8'h6b;        memory[13765] <=  8'h73;        memory[13766] <=  8'h68;        memory[13767] <=  8'h63;        memory[13768] <=  8'h66;        memory[13769] <=  8'h69;        memory[13770] <=  8'h77;        memory[13771] <=  8'h68;        memory[13772] <=  8'h61;        memory[13773] <=  8'h74;        memory[13774] <=  8'h61;        memory[13775] <=  8'h6e;        memory[13776] <=  8'h61;        memory[13777] <=  8'h62;        memory[13778] <=  8'h61;        memory[13779] <=  8'h63;        memory[13780] <=  8'h61;        memory[13781] <=  8'h74;        memory[13782] <=  8'h61;        memory[13783] <=  8'h62;        memory[13784] <=  8'h61;        memory[13785] <=  8'h72;        memory[13786] <=  8'h63;        memory[13787] <=  8'h61;        memory[13788] <=  8'h68;        memory[13789] <=  8'h64;        memory[13790] <=  8'h75;        memory[13791] <=  8'h63;        memory[13792] <=  8'h74;        memory[13793] <=  8'h61;        memory[13794] <=  8'h64;        memory[13795] <=  8'h61;        memory[13796] <=  8'h61;        memory[13797] <=  8'h63;        memory[13798] <=  8'h61;        memory[13799] <=  8'h72;        memory[13800] <=  8'h62;        memory[13801] <=  8'h61;        memory[13802] <=  8'h72;        memory[13803] <=  8'h74;        memory[13804] <=  8'h78;        memory[13805] <=  8'h61;        memory[13806] <=  8'h74;        memory[13807] <=  8'h6b;        memory[13808] <=  8'h73;        memory[13809] <=  8'h68;        memory[13810] <=  8'h63;        memory[13811] <=  8'h66;        memory[13812] <=  8'h69;        memory[13813] <=  8'h77;        memory[13814] <=  8'h68;        memory[13815] <=  8'h61;        memory[13816] <=  8'h74;        memory[13817] <=  8'h61;        memory[13818] <=  8'h6e;        memory[13819] <=  8'h61;        memory[13820] <=  8'h62;        memory[13821] <=  8'h61;        memory[13822] <=  8'h63;        memory[13823] <=  8'h61;        memory[13824] <=  8'h74;        memory[13825] <=  8'h61;        memory[13826] <=  8'h62;        memory[13827] <=  8'h61;        memory[13828] <=  8'h72;        memory[13829] <=  8'h63;        memory[13830] <=  8'h61;        memory[13831] <=  8'h68;        memory[13832] <=  8'h64;        memory[13833] <=  8'h75;        memory[13834] <=  8'h63;        memory[13835] <=  8'h74;        memory[13836] <=  8'h61;        memory[13837] <=  8'h64;        memory[13838] <=  8'h61;        memory[13839] <=  8'h61;        memory[13840] <=  8'h63;        memory[13841] <=  8'h61;        memory[13842] <=  8'h72;        memory[13843] <=  8'h62;        memory[13844] <=  8'h61;        memory[13845] <=  8'h72;        memory[13846] <=  8'h74;        memory[13847] <=  8'h78;        memory[13848] <=  8'h61;        memory[13849] <=  8'h74;        memory[13850] <=  8'h6b;        memory[13851] <=  8'h73;        memory[13852] <=  8'h68;        memory[13853] <=  8'h63;        memory[13854] <=  8'h66;        memory[13855] <=  8'h69;        memory[13856] <=  8'h77;        memory[13857] <=  8'h68;        memory[13858] <=  8'h61;        memory[13859] <=  8'h74;        memory[13860] <=  8'h61;        memory[13861] <=  8'h6e;        memory[13862] <=  8'h61;        memory[13863] <=  8'h62;        memory[13864] <=  8'h61;        memory[13865] <=  8'h63;        memory[13866] <=  8'h61;        memory[13867] <=  8'h74;        memory[13868] <=  8'h61;        memory[13869] <=  8'h62;        memory[13870] <=  8'h61;        memory[13871] <=  8'h72;        memory[13872] <=  8'h63;        memory[13873] <=  8'h61;        memory[13874] <=  8'h68;        memory[13875] <=  8'h64;        memory[13876] <=  8'h75;        memory[13877] <=  8'h63;        memory[13878] <=  8'h74;        memory[13879] <=  8'h61;        memory[13880] <=  8'h64;        memory[13881] <=  8'h61;        memory[13882] <=  8'h61;        memory[13883] <=  8'h63;        memory[13884] <=  8'h61;        memory[13885] <=  8'h72;        memory[13886] <=  8'h62;        memory[13887] <=  8'h61;        memory[13888] <=  8'h72;        memory[13889] <=  8'h74;        memory[13890] <=  8'h78;        memory[13891] <=  8'h61;        memory[13892] <=  8'h74;        memory[13893] <=  8'h6b;        memory[13894] <=  8'h73;        memory[13895] <=  8'h68;        memory[13896] <=  8'h63;        memory[13897] <=  8'h66;        memory[13898] <=  8'h69;        memory[13899] <=  8'h77;        memory[13900] <=  8'h68;        memory[13901] <=  8'h61;        memory[13902] <=  8'h74;        memory[13903] <=  8'h61;        memory[13904] <=  8'h6e;        memory[13905] <=  8'h61;        memory[13906] <=  8'h62;        memory[13907] <=  8'h61;        memory[13908] <=  8'h63;        memory[13909] <=  8'h61;        memory[13910] <=  8'h74;        memory[13911] <=  8'h61;        memory[13912] <=  8'h62;        memory[13913] <=  8'h61;        memory[13914] <=  8'h72;        memory[13915] <=  8'h63;        memory[13916] <=  8'h61;        memory[13917] <=  8'h68;        memory[13918] <=  8'h64;        memory[13919] <=  8'h75;        memory[13920] <=  8'h63;        memory[13921] <=  8'h74;        memory[13922] <=  8'h61;        memory[13923] <=  8'h64;        memory[13924] <=  8'h61;        memory[13925] <=  8'h61;        memory[13926] <=  8'h63;        memory[13927] <=  8'h61;        memory[13928] <=  8'h72;        memory[13929] <=  8'h62;        memory[13930] <=  8'h61;        memory[13931] <=  8'h72;        memory[13932] <=  8'h74;        memory[13933] <=  8'h78;        memory[13934] <=  8'h61;        memory[13935] <=  8'h74;        memory[13936] <=  8'h6b;        memory[13937] <=  8'h73;        memory[13938] <=  8'h68;        memory[13939] <=  8'h63;        memory[13940] <=  8'h66;        memory[13941] <=  8'h69;        memory[13942] <=  8'h77;        memory[13943] <=  8'h68;        memory[13944] <=  8'h61;        memory[13945] <=  8'h74;        memory[13946] <=  8'h61;        memory[13947] <=  8'h6e;        memory[13948] <=  8'h61;        memory[13949] <=  8'h62;        memory[13950] <=  8'h61;        memory[13951] <=  8'h63;        memory[13952] <=  8'h61;        memory[13953] <=  8'h74;        memory[13954] <=  8'h61;        memory[13955] <=  8'h62;        memory[13956] <=  8'h61;        memory[13957] <=  8'h72;        memory[13958] <=  8'h63;        memory[13959] <=  8'h61;        memory[13960] <=  8'h68;        memory[13961] <=  8'h64;        memory[13962] <=  8'h75;        memory[13963] <=  8'h63;        memory[13964] <=  8'h74;        memory[13965] <=  8'h61;        memory[13966] <=  8'h64;        memory[13967] <=  8'h61;        memory[13968] <=  8'h61;        memory[13969] <=  8'h63;        memory[13970] <=  8'h61;        memory[13971] <=  8'h72;        memory[13972] <=  8'h62;        memory[13973] <=  8'h61;        memory[13974] <=  8'h72;        memory[13975] <=  8'h74;        memory[13976] <=  8'h78;        memory[13977] <=  8'h61;        memory[13978] <=  8'h74;        memory[13979] <=  8'h6b;        memory[13980] <=  8'h73;        memory[13981] <=  8'h68;        memory[13982] <=  8'h63;        memory[13983] <=  8'h66;        memory[13984] <=  8'h69;        memory[13985] <=  8'h77;        memory[13986] <=  8'h68;        memory[13987] <=  8'h61;        memory[13988] <=  8'h74;        memory[13989] <=  8'h61;        memory[13990] <=  8'h6e;        memory[13991] <=  8'h61;        memory[13992] <=  8'h62;        memory[13993] <=  8'h61;        memory[13994] <=  8'h63;        memory[13995] <=  8'h61;        memory[13996] <=  8'h74;        memory[13997] <=  8'h61;        memory[13998] <=  8'h62;        memory[13999] <=  8'h61;        memory[14000] <=  8'h72;        memory[14001] <=  8'h63;        memory[14002] <=  8'h61;        memory[14003] <=  8'h68;        memory[14004] <=  8'h64;        memory[14005] <=  8'h75;        memory[14006] <=  8'h63;        memory[14007] <=  8'h74;        memory[14008] <=  8'h61;        memory[14009] <=  8'h64;        memory[14010] <=  8'h61;        memory[14011] <=  8'h61;        memory[14012] <=  8'h63;        memory[14013] <=  8'h61;        memory[14014] <=  8'h72;        memory[14015] <=  8'h62;        memory[14016] <=  8'h61;        memory[14017] <=  8'h72;        memory[14018] <=  8'h74;        memory[14019] <=  8'h78;        memory[14020] <=  8'h61;        memory[14021] <=  8'h74;        memory[14022] <=  8'h6b;        memory[14023] <=  8'h73;        memory[14024] <=  8'h68;        memory[14025] <=  8'h63;        memory[14026] <=  8'h66;        memory[14027] <=  8'h69;        memory[14028] <=  8'h77;        memory[14029] <=  8'h68;        memory[14030] <=  8'h61;        memory[14031] <=  8'h74;        memory[14032] <=  8'h61;        memory[14033] <=  8'h6e;        memory[14034] <=  8'h61;        memory[14035] <=  8'h62;        memory[14036] <=  8'h61;        memory[14037] <=  8'h63;        memory[14038] <=  8'h61;        memory[14039] <=  8'h74;        memory[14040] <=  8'h61;        memory[14041] <=  8'h62;        memory[14042] <=  8'h61;        memory[14043] <=  8'h72;        memory[14044] <=  8'h63;        memory[14045] <=  8'h61;        memory[14046] <=  8'h68;        memory[14047] <=  8'h64;        memory[14048] <=  8'h75;        memory[14049] <=  8'h63;        memory[14050] <=  8'h74;        memory[14051] <=  8'h61;        memory[14052] <=  8'h64;        memory[14053] <=  8'h61;        memory[14054] <=  8'h61;        memory[14055] <=  8'h63;        memory[14056] <=  8'h61;        memory[14057] <=  8'h72;        memory[14058] <=  8'h62;        memory[14059] <=  8'h61;        memory[14060] <=  8'h72;        memory[14061] <=  8'h74;        memory[14062] <=  8'h78;        memory[14063] <=  8'h61;        memory[14064] <=  8'h74;        memory[14065] <=  8'h6b;        memory[14066] <=  8'h73;        memory[14067] <=  8'h68;        memory[14068] <=  8'h63;        memory[14069] <=  8'h66;        memory[14070] <=  8'h69;        memory[14071] <=  8'h77;        memory[14072] <=  8'h68;        memory[14073] <=  8'h61;        memory[14074] <=  8'h74;        memory[14075] <=  8'h61;        memory[14076] <=  8'h6e;        memory[14077] <=  8'h61;        memory[14078] <=  8'h62;        memory[14079] <=  8'h61;        memory[14080] <=  8'h63;        memory[14081] <=  8'h61;        memory[14082] <=  8'h74;        memory[14083] <=  8'h61;        memory[14084] <=  8'h62;        memory[14085] <=  8'h61;        memory[14086] <=  8'h72;        memory[14087] <=  8'h63;        memory[14088] <=  8'h61;        memory[14089] <=  8'h68;        memory[14090] <=  8'h64;        memory[14091] <=  8'h75;        memory[14092] <=  8'h63;        memory[14093] <=  8'h74;        memory[14094] <=  8'h61;        memory[14095] <=  8'h64;        memory[14096] <=  8'h61;        memory[14097] <=  8'h61;        memory[14098] <=  8'h63;        memory[14099] <=  8'h61;        memory[14100] <=  8'h72;        memory[14101] <=  8'h62;        memory[14102] <=  8'h61;        memory[14103] <=  8'h72;        memory[14104] <=  8'h74;        memory[14105] <=  8'h74;        memory[14106] <=  8'h62;        memory[14107] <=  8'h61;        memory[14108] <=  8'h72;        memory[14109] <=  8'h74;        memory[14110] <=  8'h78;        memory[14111] <=  8'h61;        memory[14112] <=  8'h74;        memory[14113] <=  8'h6b;        memory[14114] <=  8'h73;        memory[14115] <=  8'h68;        memory[14116] <=  8'h63;        memory[14117] <=  8'h66;        memory[14118] <=  8'h69;        memory[14119] <=  8'h77;        memory[14120] <=  8'h68;        memory[14121] <=  8'h61;        memory[14122] <=  8'h74;        memory[14123] <=  8'h61;        memory[14124] <=  8'h6e;        memory[14125] <=  8'h61;        memory[14126] <=  8'h62;        memory[14127] <=  8'h61;        memory[14128] <=  8'h63;        memory[14129] <=  8'h61;        memory[14130] <=  8'h74;        memory[14131] <=  8'h61;        memory[14132] <=  8'h62;        memory[14133] <=  8'h61;        memory[14134] <=  8'h72;        memory[14135] <=  8'h63;        memory[14136] <=  8'h61;        memory[14137] <=  8'h68;        memory[14138] <=  8'h64;        memory[14139] <=  8'h75;        memory[14140] <=  8'h63;        memory[14141] <=  8'h74;        memory[14142] <=  8'h61;        memory[14143] <=  8'h64;        memory[14144] <=  8'h61;        memory[14145] <=  8'h61;        memory[14146] <=  8'h63;        memory[14147] <=  8'h61;        memory[14148] <=  8'h72;        memory[14149] <=  8'h63;        memory[14150] <=  8'h74;        memory[14151] <=  8'h72;        memory[14152] <=  8'h63;        memory[14153] <=  8'h61;        memory[14154] <=  8'h74;        memory[14155] <=  8'h72;        memory[14156] <=  8'h63;        memory[14157] <=  8'h61;        memory[14158] <=  8'h74;        memory[14159] <=  8'h63;        memory[14160] <=  8'h62;        memory[14161] <=  8'h61;        memory[14162] <=  8'h74;        memory[14163] <=  8'h62;        memory[14164] <=  8'h72;        memory[14165] <=  8'h63;        memory[14166] <=  8'h61;        memory[14167] <=  8'h72;        memory[14168] <=  8'h62;        memory[14169] <=  8'h78;        memory[14170] <=  8'h74;        memory[14171] <=  8'h61;        memory[14172] <=  8'h72;        memory[14173] <=  8'h64;        memory[14174] <=  8'h66;        memory[14175] <=  8'h73;        memory[14176] <=  8'h67;        memory[14177] <=  8'h76;        memory[14178] <=  8'h68;        memory[14179] <=  8'h62;        memory[14180] <=  8'h6b;        memory[14181] <=  8'h6a;        memory[14182] <=  8'h6e;        memory[14183] <=  8'h6d;        memory[14184] <=  8'h62;        memory[14185] <=  8'h76;        memory[14186] <=  8'h78;        memory[14187] <=  8'h63;        memory[14188] <=  8'h73;        memory[14189] <=  8'h66;        memory[14190] <=  8'h72;        memory[14191] <=  8'h74;        memory[14192] <=  8'h79;        memory[14193] <=  8'h75;        memory[14194] <=  8'h6a;        memory[14195] <=  8'h6e;        memory[14196] <=  8'h62;        memory[14197] <=  8'h76;        memory[14198] <=  8'h63;        memory[14199] <=  8'h64;        memory[14200] <=  8'h74;        memory[14201] <=  8'h79;        memory[14202] <=  8'h75;        memory[14203] <=  8'h69;        memory[14204] <=  8'h6b;        memory[14205] <=  8'h6d;        memory[14206] <=  8'h6e;        memory[14207] <=  8'h62;        memory[14208] <=  8'h76;        memory[14209] <=  8'h63;        memory[14210] <=  8'h78;        memory[14211] <=  8'h73;        memory[14212] <=  8'h64;        memory[14213] <=  8'h72;        memory[14214] <=  8'h74;        memory[14215] <=  8'h79;        memory[14216] <=  8'h75;        memory[14217] <=  8'h69;        memory[14218] <=  8'h6b;        memory[14219] <=  8'h6d;        memory[14220] <=  8'h6e;        memory[14221] <=  8'h62;        memory[14222] <=  8'h76;        memory[14223] <=  8'h63;        memory[14224] <=  8'h73;        memory[14225] <=  8'h77;        memory[14226] <=  8'h33;        memory[14227] <=  8'h34;        memory[14228] <=  8'h35;        memory[14229] <=  8'h36;        memory[14230] <=  8'h37;        memory[14231] <=  8'h38;        memory[14232] <=  8'h69;        memory[14233] <=  8'h6b;        memory[14234] <=  8'h6d;        memory[14235] <=  8'h6e;        memory[14236] <=  8'h62;        memory[14237] <=  8'h76;        memory[14238] <=  8'h63;        memory[14239] <=  8'h64;        memory[14240] <=  8'h65;        memory[14241] <=  8'h72;        memory[14242] <=  8'h36;        memory[14243] <=  8'h37;        memory[14244] <=  8'h38;        memory[14245] <=  8'h69;        memory[14246] <=  8'h6f;        memory[14247] <=  8'h6b;        memory[14248] <=  8'h6a;        memory[14249] <=  8'h6e;        memory[14250] <=  8'h62;        memory[14251] <=  8'h76;        memory[14252] <=  8'h63;        memory[14253] <=  8'h64;        memory[14254] <=  8'h72;        memory[14255] <=  8'h74;        memory[14256] <=  8'h79;        memory[14257] <=  8'h75;        memory[14258] <=  8'h73;        memory[14259] <=  8'h6a;        memory[14260] <=  8'h63;        memory[14261] <=  8'h6e;        memory[14262] <=  8'h62;        memory[14263] <=  8'h64;        memory[14264] <=  8'h66;        memory[14265] <=  8'h73;        memory[14266] <=  8'h74;        memory[14267] <=  8'h79;        memory[14268] <=  8'h75;        memory[14269] <=  8'h61;        memory[14270] <=  8'h69;        memory[14271] <=  8'h6b;        memory[14272] <=  8'h78;        memory[14273] <=  8'h6d;        memory[14274] <=  8'h6e;        memory[14275] <=  8'h73;        memory[14276] <=  8'h6a;        memory[14277] <=  8'h6f;        memory[14278] <=  8'h64;        memory[14279] <=  8'h6c;        memory[14280] <=  8'h63;        memory[14281] <=  8'h78;        memory[14282] <=  8'h2c;        memory[14283] <=  8'h6d;        memory[14284] <=  8'h73;        memory[14285] <=  8'h6b;        memory[14286] <=  8'h64;        memory[14287] <=  8'h6c;        memory[14288] <=  8'h70;        memory[14289] <=  8'h5b;        memory[14290] <=  8'h3b;        memory[14291] <=  8'h73;        memory[14292] <=  8'h6c;        memory[14293] <=  8'h64;        memory[14294] <=  8'h70;        memory[14295] <=  8'h76;        memory[14296] <=  8'h63;        memory[14297] <=  8'h5b;        memory[14298] <=  8'h78;        memory[14299] <=  8'h76;        memory[14300] <=  8'h63;        memory[14301] <=  8'h5b;        memory[14302] <=  8'h78;        memory[14303] <=  8'h70;        memory[14304] <=  8'h6f;        memory[14305] <=  8'h20;        memory[14306] <=  8'h62;        memory[14307] <=  8'h61;        memory[14308] <=  8'h72;        memory[14309] <=  8'h74;        memory[14310] <=  8'h74;        memory[14311] <=  8'h62;        memory[14312] <=  8'h61;        memory[14313] <=  8'h72;        memory[14314] <=  8'h74;        memory[14315] <=  8'h78;        memory[14316] <=  8'h61;        memory[14317] <=  8'h74;        memory[14318] <=  8'h6b;        memory[14319] <=  8'h73;        memory[14320] <=  8'h68;        memory[14321] <=  8'h63;        memory[14322] <=  8'h66;        memory[14323] <=  8'h69;        memory[14324] <=  8'h77;        memory[14325] <=  8'h68;        memory[14326] <=  8'h61;        memory[14327] <=  8'h69;        memory[14328] <=  8'h6a;        memory[14329] <=  8'h78;        memory[14330] <=  8'h5d;        memory[14331] <=  8'h65;        memory[14332] <=  8'h6b;        memory[14333] <=  8'h6f;        memory[14334] <=  8'h39;        memory[14335] <=  8'h64;        memory[14336] <=  8'h75;        memory[14337] <=  8'h38;        memory[14338] <=  8'h79;        memory[14339] <=  8'h20;        memory[14340] <=  8'h37;        memory[14341] <=  8'h63;        memory[14342] <=  8'h67;        memory[14343] <=  8'h78;        memory[14344] <=  8'h63;        memory[14345] <=  8'h75;        memory[14346] <=  8'h68;        memory[14347] <=  8'h69;        memory[14348] <=  8'h6a;        memory[14349] <=  8'h77;        memory[14350] <=  8'h69;        memory[14351] <=  8'h64;        memory[14352] <=  8'h66;        memory[14353] <=  8'h68;        memory[14354] <=  8'h75;        memory[14355] <=  8'h76;        memory[14356] <=  8'h64;        memory[14357] <=  8'h62;        memory[14358] <=  8'h66;        memory[14359] <=  8'h6a;        memory[14360] <=  8'h6e;        memory[14361] <=  8'h6b;        memory[14362] <=  8'h6a;        memory[14363] <=  8'h65;        memory[14364] <=  8'h38;        memory[14365] <=  8'h66;        memory[14366] <=  8'h37;        memory[14367] <=  8'h67;        memory[14368] <=  8'h79;        memory[14369] <=  8'h76;        memory[14370] <=  8'h63;        memory[14371] <=  8'h68;        memory[14372] <=  8'h69;        memory[14373] <=  8'h6a;        memory[14374] <=  8'h33;        memory[14375] <=  8'h65;        memory[14376] <=  8'h67;        memory[14377] <=  8'h79;        memory[14378] <=  8'h72;        memory[14379] <=  8'h64;        memory[14380] <=  8'h62;        memory[14381] <=  8'h6e;        memory[14382] <=  8'h63;        memory[14383] <=  8'h7a;        memory[14384] <=  8'h6a;        memory[14385] <=  8'h6f;        memory[14386] <=  8'h66;        memory[14387] <=  8'h78;        memory[14388] <=  8'h6a;        memory[14389] <=  8'h69;        memory[14390] <=  8'h63;        memory[14391] <=  8'h68;        memory[14392] <=  8'h62;        memory[14393] <=  8'h6e;        memory[14394] <=  8'h6d;        memory[14395] <=  8'h63;        memory[14396] <=  8'h73;        memory[14397] <=  8'h6c;        memory[14398] <=  8'h6b;        memory[14399] <=  8'h6a;        memory[14400] <=  8'h69;        memory[14401] <=  8'h68;        memory[14402] <=  8'h76;        memory[14403] <=  8'h75;        memory[14404] <=  8'h69;        memory[14405] <=  8'h64;        memory[14406] <=  8'h68;        memory[14407] <=  8'h75;        memory[14408] <=  8'h67;        memory[14409] <=  8'h79;        memory[14410] <=  8'h62;        memory[14411] <=  8'h68;        memory[14412] <=  8'h65;        memory[14413] <=  8'h6a;        memory[14414] <=  8'h72;        memory[14415] <=  8'h6b;        memory[14416] <=  8'h6a;        memory[14417] <=  8'h6f;        memory[14418] <=  8'h64;        memory[14419] <=  8'h67;        memory[14420] <=  8'h69;        memory[14421] <=  8'h75;        memory[14422] <=  8'h69;        memory[14423] <=  8'h67;        memory[14424] <=  8'h76;        memory[14425] <=  8'h79;        memory[14426] <=  8'h75;        memory[14427] <=  8'h67;        memory[14428] <=  8'h78;        memory[14429] <=  8'h68;        memory[14430] <=  8'h63;        memory[14431] <=  8'h20;        memory[14432] <=  8'h20;        memory[14433] <=  8'h20;        memory[14434] <=  8'h78;        memory[14435] <=  8'h76;        memory[14436] <=  8'h20;        memory[14437] <=  8'h63;        memory[14438] <=  8'h78;        memory[14439] <=  8'h67;        memory[14440] <=  8'h79;        memory[14441] <=  8'h63;        memory[14442] <=  8'h75;        memory[14443] <=  8'h68;        memory[14444] <=  8'h6a;        memory[14445] <=  8'h6b;        memory[14446] <=  8'h61;        memory[14447] <=  8'h6c;        memory[14448] <=  8'h78;        memory[14449] <=  8'h76;        memory[14450] <=  8'h70;        memory[14451] <=  8'h6f;        memory[14452] <=  8'h69;        memory[14453] <=  8'h6a;        memory[14454] <=  8'h69;        memory[14455] <=  8'h68;        memory[14456] <=  8'h6a;        memory[14457] <=  8'h62;        memory[14458] <=  8'h77;        memory[14459] <=  8'h65;        memory[14460] <=  8'h6e;        memory[14461] <=  8'h61;        memory[14462] <=  8'h66;        memory[14463] <=  8'h6d;        memory[14464] <=  8'h64;        memory[14465] <=  8'h6b;        memory[14466] <=  8'h6d;        memory[14467] <=  8'h76;        memory[14468] <=  8'h6c;        memory[14469] <=  8'h63;        memory[14470] <=  8'h6f;        memory[14471] <=  8'h64;        memory[14472] <=  8'h69;        memory[14473] <=  8'h75;        memory[14474] <=  8'h68;        memory[14475] <=  8'h73;        memory[14476] <=  8'h66;        memory[14477] <=  8'h65;        memory[14478] <=  8'h62;        memory[14479] <=  8'h6e;        memory[14480] <=  8'h64;        memory[14481] <=  8'h73;        memory[14482] <=  8'h63;        memory[14483] <=  8'h6b;        memory[14484] <=  8'h20;        memory[14485] <=  8'h78;        memory[14486] <=  8'h6a;        memory[14487] <=  8'h78;        memory[14488] <=  8'h63;        memory[14489] <=  8'h73;        memory[14490] <=  8'h64;        memory[14491] <=  8'h66;        memory[14492] <=  8'h6b;        memory[14493] <=  8'h64;        memory[14494] <=  8'h6e;        memory[14495] <=  8'h6d;        memory[14496] <=  8'h64;        memory[14497] <=  8'h73;        memory[14498] <=  8'h63;        memory[14499] <=  8'h6b;        memory[14500] <=  8'h78;        memory[14501] <=  8'h6c;        memory[14502] <=  8'h6f;        memory[14503] <=  8'h66;        memory[14504] <=  8'h6a;        memory[14505] <=  8'h69;        memory[14506] <=  8'h61;        memory[14507] <=  8'h62;        memory[14508] <=  8'h6e;        memory[14509] <=  8'h20;        memory[14510] <=  8'h78;        memory[14511] <=  8'h6b;        memory[14512] <=  8'h6d;        memory[14513] <=  8'h20;        memory[14514] <=  8'h6f;        memory[14515] <=  8'h63;        memory[14516] <=  8'h76;        memory[14517] <=  8'h73;        memory[14518] <=  8'h64;        memory[14519] <=  8'h69;        memory[14520] <=  8'h66;        memory[14521] <=  8'h68;        memory[14522] <=  8'h65;        memory[14523] <=  8'h71;        memory[14524] <=  8'h6a;        memory[14525] <=  8'h77;        memory[14526] <=  8'h62;        memory[14527] <=  8'h65;        memory[14528] <=  8'h6e;        memory[14529] <=  8'h20;        memory[14530] <=  8'h6d;        memory[14531] <=  8'h64;        memory[14532] <=  8'h73;        memory[14533] <=  8'h6c;        memory[14534] <=  8'h76;        memory[14535] <=  8'h6b;        memory[14536] <=  8'h63;        memory[14537] <=  8'h78;        memory[14538] <=  8'h20;        memory[14539] <=  8'h6f;        memory[14540] <=  8'h78;        memory[14541] <=  8'h69;        memory[14542] <=  8'h63;        memory[14543] <=  8'h6a;        memory[14544] <=  8'h76;        memory[14545] <=  8'h64;        memory[14546] <=  8'h66;        memory[14547] <=  8'h65;        memory[14548] <=  8'h71;        memory[14549] <=  8'h6e;        memory[14550] <=  8'h20;        memory[14551] <=  8'h64;        memory[14552] <=  8'h6d;        memory[14553] <=  8'h73;        memory[14554] <=  8'h6c;        memory[14555] <=  8'h63;        memory[14556] <=  8'h78;        memory[14557] <=  8'h6b;        memory[14558] <=  8'h20;        memory[14559] <=  8'h6f;        memory[14560] <=  8'h78;        memory[14561] <=  8'h63;        memory[14562] <=  8'h76;        memory[14563] <=  8'h6a;        memory[14564] <=  8'h64;        memory[14565] <=  8'h62;        memory[14566] <=  8'h71;        memory[14567] <=  8'h77;        memory[14568] <=  8'h65;        memory[14569] <=  8'h6e;        memory[14570] <=  8'h6d;        memory[14571] <=  8'h64;        memory[14572] <=  8'h6c;        memory[14573] <=  8'h73;        memory[14574] <=  8'h2c;        memory[14575] <=  8'h76;        memory[14576] <=  8'h63;        memory[14577] <=  8'h78;        memory[14578] <=  8'h20;        memory[14579] <=  8'h63;        memory[14580] <=  8'h6f;        memory[14581] <=  8'h69;        memory[14582] <=  8'h76;        memory[14583] <=  8'h68;        memory[14584] <=  8'h73;        memory[14585] <=  8'h64;        memory[14586] <=  8'h62;        memory[14587] <=  8'h71;        memory[14588] <=  8'h77;        memory[14589] <=  8'h65;        memory[14590] <=  8'h6e;        memory[14591] <=  8'h64;        memory[14592] <=  8'h6b;        memory[14593] <=  8'h73;        memory[14594] <=  8'h76;        memory[14595] <=  8'h6f;        memory[14596] <=  8'h63;        memory[14597] <=  8'h20;        memory[14598] <=  8'h76;        memory[14599] <=  8'h69;        memory[14600] <=  8'h75;        memory[14601] <=  8'h69;        memory[14602] <=  8'h68;        memory[14603] <=  8'h63;        memory[14604] <=  8'h78;        memory[14605] <=  8'h69;        memory[14606] <=  8'h6f;        memory[14607] <=  8'h76;        memory[14608] <=  8'h73;        memory[14609] <=  8'h64;        memory[14610] <=  8'h61;        memory[14611] <=  8'h64;        memory[14612] <=  8'h6e;        memory[14613] <=  8'h77;        memory[14614] <=  8'h71;        memory[14615] <=  8'h6b;        memory[14616] <=  8'h6c;        memory[14617] <=  8'h73;        memory[14618] <=  8'h76;        memory[14619] <=  8'h6e;        memory[14620] <=  8'h62;        memory[14621] <=  8'h20;        memory[14622] <=  8'h64;        memory[14623] <=  8'h66;        memory[14624] <=  8'h6a;        memory[14625] <=  8'h6b;        memory[14626] <=  8'h71;        memory[14627] <=  8'h64;        memory[14628] <=  8'h77;        memory[14629] <=  8'h65;        memory[14630] <=  8'h6e;        memory[14631] <=  8'h62;        memory[14632] <=  8'h20;        memory[14633] <=  8'h64;        memory[14634] <=  8'h73;        memory[14635] <=  8'h76;        memory[14636] <=  8'h68;        memory[14637] <=  8'h64;        memory[14638] <=  8'h61;        memory[14639] <=  8'h71;        memory[14640] <=  8'h77;        memory[14641] <=  8'h6a;        memory[14642] <=  8'h65;        memory[14643] <=  8'h6e;        memory[14644] <=  8'h64;        memory[14645] <=  8'h20;        memory[14646] <=  8'h61;        memory[14647] <=  8'h63;        memory[14648] <=  8'h62;        memory[14649] <=  8'h68;        memory[14650] <=  8'h64;        memory[14651] <=  8'h61;        memory[14652] <=  8'h77;        memory[14653] <=  8'h71;        memory[14654] <=  8'h6e;        memory[14655] <=  8'h20;        memory[14656] <=  8'h62;        memory[14657] <=  8'h73;        memory[14658] <=  8'h76;        memory[14659] <=  8'h61;        memory[14660] <=  8'h67;        memory[14661] <=  8'h76;        memory[14662] <=  8'h68;        memory[14663] <=  8'h67;        memory[14664] <=  8'h61;        memory[14665] <=  8'h73;        memory[14666] <=  8'h6a;        memory[14667] <=  8'h6b;        memory[14668] <=  8'h63;        memory[14669] <=  8'h78;        memory[14670] <=  8'h76;        memory[14671] <=  8'h6e;        memory[14672] <=  8'h73;        memory[14673] <=  8'h64;        memory[14674] <=  8'h20;        memory[14675] <=  8'h66;        memory[14676] <=  8'h62;        memory[14677] <=  8'h64;        memory[14678] <=  8'h61;        memory[14679] <=  8'h73;        memory[14680] <=  8'h76;        memory[14681] <=  8'h67;        memory[14682] <=  8'h63;        memory[14683] <=  8'h79;        memory[14684] <=  8'h7a;        memory[14685] <=  8'h78;        memory[14686] <=  8'h79;        memory[14687] <=  8'h75;        memory[14688] <=  8'h20;        memory[14689] <=  8'h69;        memory[14690] <=  8'h6a;        memory[14691] <=  8'h64;        memory[14692] <=  8'h66;        memory[14693] <=  8'h6b;        memory[14694] <=  8'h61;        memory[14695] <=  8'h64;        memory[14696] <=  8'h63;        memory[14697] <=  8'h78;        memory[14698] <=  8'h68;        memory[14699] <=  8'h20;        memory[14700] <=  8'h67;        memory[14701] <=  8'h61;        memory[14702] <=  8'h68;        memory[14703] <=  8'h75;        memory[14704] <=  8'h64;        memory[14705] <=  8'h73;        memory[14706] <=  8'h69;        memory[14707] <=  8'h6a;        memory[14708] <=  8'h61;        memory[14709] <=  8'h6b;        memory[14710] <=  8'h63;        memory[14711] <=  8'h62;        memory[14712] <=  8'h61;        memory[14713] <=  8'h72;        memory[14714] <=  8'h73;        memory[14715] <=  8'h68;        memory[14716] <=  8'h64;        memory[14717] <=  8'h66;        memory[14718] <=  8'h67;        memory[14719] <=  8'h73;        memory[14720] <=  8'h68;        memory[14721] <=  8'h64;        memory[14722] <=  8'h66;        memory[14723] <=  8'h68;        memory[14724] <=  8'h64;        memory[14725] <=  8'h6a;        memory[14726] <=  8'h68;        memory[14727] <=  8'h62;        memory[14728] <=  8'h67;        memory[14729] <=  8'h63;        memory[14730] <=  8'h61;        memory[14731] <=  8'h66;        memory[14732] <=  8'h73;        memory[14733] <=  8'h79;        memory[14734] <=  8'h67;        memory[14735] <=  8'h6b;        memory[14736] <=  8'h75;        memory[14737] <=  8'h64;        memory[14738] <=  8'h68;        memory[14739] <=  8'h62;        memory[14740] <=  8'h77;        memory[14741] <=  8'h76;        memory[14742] <=  8'h67;        memory[14743] <=  8'h61;        memory[14744] <=  8'h66;        memory[14745] <=  8'h64;        memory[14746] <=  8'h74;        memory[14747] <=  8'h75;        memory[14748] <=  8'h66;        memory[14749] <=  8'h79;        memory[14750] <=  8'h67;        memory[14751] <=  8'h69;        memory[14752] <=  8'h75;        memory[14753] <=  8'h68;        memory[14754] <=  8'h6c;        memory[14755] <=  8'h6a;        memory[14756] <=  8'h62;        memory[14757] <=  8'h6b;        memory[14758] <=  8'h68;        memory[14759] <=  8'h76;        memory[14760] <=  8'h67;        memory[14761] <=  8'h63;        memory[14762] <=  8'h66;        memory[14763] <=  8'h78;        memory[14764] <=  8'h64;        memory[14765] <=  8'h74;        memory[14766] <=  8'h75;        memory[14767] <=  8'h79;        memory[14768] <=  8'h69;        memory[14769] <=  8'h75;        memory[14770] <=  8'h68;        memory[14771] <=  8'h6c;        memory[14772] <=  8'h6a;        memory[14773] <=  8'h6b;        memory[14774] <=  8'h67;        memory[14775] <=  8'h6a;        memory[14776] <=  8'h63;        memory[14777] <=  8'h66;        memory[14778] <=  8'h68;        memory[14779] <=  8'h64;        memory[14780] <=  8'h67;        memory[14781] <=  8'h72;        memory[14782] <=  8'h79;        memory[14783] <=  8'h74;        memory[14784] <=  8'h66;        memory[14785] <=  8'h75;        memory[14786] <=  8'h79;        memory[14787] <=  8'h69;        memory[14788] <=  8'h68;        memory[14789] <=  8'h6c;        memory[14790] <=  8'h62;        memory[14791] <=  8'h6d;        memory[14792] <=  8'h76;        memory[14793] <=  8'h6e;        memory[14794] <=  8'h63;        memory[14795] <=  8'h66;        memory[14796] <=  8'h68;        memory[14797] <=  8'h64;        memory[14798] <=  8'h74;        memory[14799] <=  8'h75;        memory[14800] <=  8'h67;        memory[14801] <=  8'h79;        memory[14802] <=  8'h69;        memory[14803] <=  8'h68;        memory[14804] <=  8'h75;        memory[14805] <=  8'h6a;        memory[14806] <=  8'h6c;        memory[14807] <=  8'h62;        memory[14808] <=  8'h6d;        memory[14809] <=  8'h76;        memory[14810] <=  8'h6e;        memory[14811] <=  8'h63;        memory[14812] <=  8'h66;        memory[14813] <=  8'h68;        memory[14814] <=  8'h67;        memory[14815] <=  8'h79;        memory[14816] <=  8'h68;        memory[14817] <=  8'h75;        memory[14818] <=  8'h6a;        memory[14819] <=  8'h6e;        memory[14820] <=  8'h2c;        memory[14821] <=  8'h62;        memory[14822] <=  8'h6e;        memory[14823] <=  8'h6d;        memory[14824] <=  8'h76;        memory[14825] <=  8'h6e;        memory[14826] <=  8'h63;        memory[14827] <=  8'h66;        memory[14828] <=  8'h68;        memory[14829] <=  8'h74;        memory[14830] <=  8'h79;        memory[14831] <=  8'h69;        memory[14832] <=  8'h75;        memory[14833] <=  8'h6c;        memory[14834] <=  8'h6a;        memory[14835] <=  8'h62;        memory[14836] <=  8'h6d;        memory[14837] <=  8'h76;        memory[14838] <=  8'h6e;        memory[14839] <=  8'h63;        memory[14840] <=  8'h66;        memory[14841] <=  8'h74;        memory[14842] <=  8'h75;        memory[14843] <=  8'h79;        memory[14844] <=  8'h69;        memory[14845] <=  8'h68;        memory[14846] <=  8'h6b;        memory[14847] <=  8'h62;        memory[14848] <=  8'h76;        memory[14849] <=  8'h63;        memory[14850] <=  8'h66;        memory[14851] <=  8'h67;        memory[14852] <=  8'h74;        memory[14853] <=  8'h75;        memory[14854] <=  8'h79;        memory[14855] <=  8'h69;        memory[14856] <=  8'h75;        memory[14857] <=  8'h68;        memory[14858] <=  8'h6a;        memory[14859] <=  8'h6b;        memory[14860] <=  8'h62;        memory[14861] <=  8'h76;        memory[14862] <=  8'h63;        memory[14863] <=  8'h66;        memory[14864] <=  8'h74;        memory[14865] <=  8'h75;        memory[14866] <=  8'h79;        memory[14867] <=  8'h69;        memory[14868] <=  8'h75;        memory[14869] <=  8'h6a;        memory[14870] <=  8'h6b;        memory[14871] <=  8'h6e;        memory[14872] <=  8'h62;        memory[14873] <=  8'h76;        memory[14874] <=  8'h67;        memory[14875] <=  8'h66;        memory[14876] <=  8'h74;        memory[14877] <=  8'h79;        memory[14878] <=  8'h75;        memory[14879] <=  8'h75;        memory[14880] <=  8'h69;        memory[14881] <=  8'h6a;        memory[14882] <=  8'h6b;        memory[14883] <=  8'h68;        memory[14884] <=  8'h62;        memory[14885] <=  8'h6a;        memory[14886] <=  8'h67;        memory[14887] <=  8'h68;        memory[14888] <=  8'h66;        memory[14889] <=  8'h79;        memory[14890] <=  8'h74;        memory[14891] <=  8'h79;        memory[14892] <=  8'h69;        memory[14893] <=  8'h75;        memory[14894] <=  8'h64;        memory[14895] <=  8'h6a;        memory[14896] <=  8'h6b;        memory[14897] <=  8'h68;        memory[14898] <=  8'h63;        memory[14899] <=  8'h7a;        memory[14900] <=  8'h67;        memory[14901] <=  8'h68;        memory[14902] <=  8'h74;        memory[14903] <=  8'h75;        memory[14904] <=  8'h79;        memory[14905] <=  8'h69;        memory[14906] <=  8'h61;        memory[14907] <=  8'h73;        memory[14908] <=  8'h75;        memory[14909] <=  8'h6a;        memory[14910] <=  8'h6b;        memory[14911] <=  8'h62;        memory[14912] <=  8'h6e;        memory[14913] <=  8'h61;        memory[14914] <=  8'h76;        memory[14915] <=  8'h63;        memory[14916] <=  8'h66;        memory[14917] <=  8'h68;        memory[14918] <=  8'h75;        memory[14919] <=  8'h61;        memory[14920] <=  8'h73;        memory[14921] <=  8'h79;        memory[14922] <=  8'h64;        memory[14923] <=  8'h75;        memory[14924] <=  8'h69;        memory[14925] <=  8'h6a;        memory[14926] <=  8'h61;        memory[14927] <=  8'h6b;        memory[14928] <=  8'h62;        memory[14929] <=  8'h63;        memory[14930] <=  8'h78;        memory[14931] <=  8'h68;        memory[14932] <=  8'h67;        memory[14933] <=  8'h79;        memory[14934] <=  8'h75;        memory[14935] <=  8'h7a;        memory[14936] <=  8'h63;        memory[14937] <=  8'h61;        memory[14938] <=  8'h73;        memory[14939] <=  8'h69;        memory[14940] <=  8'h75;        memory[14941] <=  8'h6f;        memory[14942] <=  8'h69;        memory[14943] <=  8'h6a;        memory[14944] <=  8'h61;        memory[14945] <=  8'h6c;        memory[14946] <=  8'h63;        memory[14947] <=  8'h78;        memory[14948] <=  8'h62;        memory[14949] <=  8'h63;        memory[14950] <=  8'h20;        memory[14951] <=  8'h6e;        memory[14952] <=  8'h76;        memory[14953] <=  8'h63;        memory[14954] <=  8'h61;        memory[14955] <=  8'h64;        memory[14956] <=  8'h73;        memory[14957] <=  8'h67;        memory[14958] <=  8'h79;        memory[14959] <=  8'h68;        memory[14960] <=  8'h75;        memory[14961] <=  8'h61;        memory[14962] <=  8'h6a;        memory[14963] <=  8'h6b;        memory[14964] <=  8'h78;        memory[14965] <=  8'h62;        memory[14966] <=  8'h20;        memory[14967] <=  8'h6e;        memory[14968] <=  8'h76;        memory[14969] <=  8'h63;        memory[14970] <=  8'h61;        memory[14971] <=  8'h73;        memory[14972] <=  8'h67;        memory[14973] <=  8'h68;        memory[14974] <=  8'h75;        memory[14975] <=  8'h6a;        memory[14976] <=  8'h6c;        memory[14977] <=  8'h6b;        memory[14978] <=  8'h63;        memory[14979] <=  8'h78;        memory[14980] <=  8'h20;        memory[14981] <=  8'h6a;        memory[14982] <=  8'h6b;        memory[14983] <=  8'h68;        memory[14984] <=  8'h61;        memory[14985] <=  8'h73;        memory[14986] <=  8'h76;        memory[14987] <=  8'h64;        memory[14988] <=  8'h6e;        memory[14989] <=  8'h20;        memory[14990] <=  8'h62;        memory[14991] <=  8'h6e;        memory[14992] <=  8'h6d;        memory[14993] <=  8'h6b;        memory[14994] <=  8'h77;        memory[14995] <=  8'h64;        memory[14996] <=  8'h6f;        memory[14997] <=  8'h77;        memory[14998] <=  8'h69;        memory[14999] <=  8'h6f;        memory[15000] <=  8'h75;        memory[15001] <=  8'h69;        memory[15002] <=  8'h68;        memory[15003] <=  8'h62;        memory[15004] <=  8'h6e;        memory[15005] <=  8'h6b;        memory[15006] <=  8'h77;        memory[15007] <=  8'h69;        memory[15008] <=  8'h6f;        memory[15009] <=  8'h75;        memory[15010] <=  8'h71;        memory[15011] <=  8'h69;        memory[15012] <=  8'h79;        memory[15013] <=  8'h67;        memory[15014] <=  8'h6a;        memory[15015] <=  8'h64;        memory[15016] <=  8'h61;        memory[15017] <=  8'h76;        memory[15018] <=  8'h62;        memory[15019] <=  8'h6e;        memory[15020] <=  8'h6b;        memory[15021] <=  8'h6f;        memory[15022] <=  8'h70;        memory[15023] <=  8'h64;        memory[15024] <=  8'h76;        memory[15025] <=  8'h69;        memory[15026] <=  8'h6f;        memory[15027] <=  8'h75;        memory[15028] <=  8'h69;        memory[15029] <=  8'h48;        memory[15030] <=  8'h42;        memory[15031] <=  8'h6b;        memory[15032] <=  8'h64;        memory[15033] <=  8'h6e;        memory[15034] <=  8'h6c;        memory[15035] <=  8'h71;        memory[15036] <=  8'h6b;        memory[15037] <=  8'h6d;        memory[15038] <=  8'h6a;        memory[15039] <=  8'h70;        memory[15040] <=  8'h69;        memory[15041] <=  8'h6f;        memory[15042] <=  8'h68;        memory[15043] <=  8'h65;        memory[15044] <=  8'h66;        memory[15045] <=  8'h75;        memory[15046] <=  8'h67;        memory[15047] <=  8'h69;        memory[15048] <=  8'h73;        memory[15049] <=  8'h61;        memory[15050] <=  8'h62;        memory[15051] <=  8'h64;        memory[15052] <=  8'h6b;        memory[15053] <=  8'h6a;        memory[15054] <=  8'h6b;        memory[15055] <=  8'h6c;        memory[15056] <=  8'h6a;        memory[15057] <=  8'h69;        memory[15058] <=  8'h73;        memory[15059] <=  8'h6f;        memory[15060] <=  8'h71;        memory[15061] <=  8'h68;        memory[15062] <=  8'h77;        memory[15063] <=  8'h67;        memory[15064] <=  8'h69;        memory[15065] <=  8'h79;        memory[15066] <=  8'h6a;        memory[15067] <=  8'h64;        memory[15068] <=  8'h76;        memory[15069] <=  8'h62;        memory[15070] <=  8'h6e;        memory[15071] <=  8'h61;        memory[15072] <=  8'h73;        memory[15073] <=  8'h66;        memory[15074] <=  8'h6c;        memory[15075] <=  8'h6b;        memory[15076] <=  8'h64;        memory[15077] <=  8'h6a;        memory[15078] <=  8'h68;        memory[15079] <=  8'h63;        memory[15080] <=  8'h67;        memory[15081] <=  8'h6a;        memory[15082] <=  8'h76;        memory[15083] <=  8'h73;        memory[15084] <=  8'h64;        memory[15085] <=  8'h62;        memory[15086] <=  8'h62;        memory[15087] <=  8'h61;        memory[15088] <=  8'h72;        memory[15089] <=  8'h62;        memory[15090] <=  8'h62;        memory[15091] <=  8'h73;        memory[15092] <=  8'h62;        memory[15093] <=  8'h67;        memory[15094] <=  8'h73;        memory[15095] <=  8'h66;        memory[15096] <=  8'h67;        memory[15097] <=  8'h61;        memory[15098] <=  8'h68;        memory[15099] <=  8'h66;        memory[15100] <=  8'h73;        memory[15101] <=  8'h68;        memory[15102] <=  8'h61;        memory[15103] <=  8'h66;        memory[15104] <=  8'h73;        memory[15105] <=  8'h66;        memory[15106] <=  8'h68;        memory[15107] <=  8'h61;        memory[15108] <=  8'h69;        memory[15109] <=  8'h64;        memory[15110] <=  8'h75;        memory[15111] <=  8'h67;        memory[15112] <=  8'h64;        memory[15113] <=  8'h77;        memory[15114] <=  8'h62;        memory[15115] <=  8'h61;        memory[15116] <=  8'h62;        memory[15117] <=  8'h72;        memory[15118] <=  8'h62;        memory[15119] <=  8'h61;        memory[15120] <=  8'h62;        memory[15121] <=  8'h62;        memory[15122] <=  8'h74;        memory[15123] <=  8'h62;        memory[15124] <=  8'h62;        memory[15125] <=  8'h62;        memory[15126] <=  8'h62;        memory[15127] <=  8'h62;        memory[15128] <=  8'h62;        memory[15129] <=  8'h62;        memory[15130] <=  8'h62;        memory[15131] <=  8'h61;        memory[15132] <=  8'h62;        memory[15133] <=  8'h62;        memory[15134] <=  8'h72;        memory[15135] <=  8'h74;        memory[15136] <=  8'h62;        memory[15137] <=  8'h62;        memory[15138] <=  8'h61;        memory[15139] <=  8'h62;        memory[15140] <=  8'h72;        memory[15141] <=  8'h62;        memory[15142] <=  8'h74;        memory[15143] <=  8'h62;        memory[15144] <=  8'h62;        memory[15145] <=  8'h62;        memory[15146] <=  8'h63;        memory[15147] <=  8'h61;        memory[15148] <=  8'h72;        memory[15149] <=  8'h74;        memory[15150] <=  8'h73;        memory[15151] <=  8'h62;        memory[15152] <=  8'h61;        memory[15153] <=  8'h72;        memory[15154] <=  8'h74;        memory[15155] <=  8'h74;        memory[15156] <=  8'h62;        memory[15157] <=  8'h61;        memory[15158] <=  8'h72;        memory[15159] <=  8'h74;        memory[15160] <=  8'h78;        memory[15161] <=  8'h61;        memory[15162] <=  8'h74;        memory[15163] <=  8'h6b;        memory[15164] <=  8'h73;        memory[15165] <=  8'h68;        memory[15166] <=  8'h63;        memory[15167] <=  8'h66;        memory[15168] <=  8'h69;        memory[15169] <=  8'h77;        memory[15170] <=  8'h68;        memory[15171] <=  8'h61;        memory[15172] <=  8'h74;        memory[15173] <=  8'h61;        memory[15174] <=  8'h6e;        memory[15175] <=  8'h61;        memory[15176] <=  8'h62;        memory[15177] <=  8'h61;        memory[15178] <=  8'h63;        memory[15179] <=  8'h61;        memory[15180] <=  8'h74;        memory[15181] <=  8'h61;        memory[15182] <=  8'h62;        memory[15183] <=  8'h61;        memory[15184] <=  8'h72;        memory[15185] <=  8'h63;        memory[15186] <=  8'h61;        memory[15187] <=  8'h68;        memory[15188] <=  8'h64;        memory[15189] <=  8'h75;        memory[15190] <=  8'h63;        memory[15191] <=  8'h74;        memory[15192] <=  8'h61;        memory[15193] <=  8'h64;        memory[15194] <=  8'h61;        memory[15195] <=  8'h61;        memory[15196] <=  8'h63;        memory[15197] <=  8'h61;        memory[15198] <=  8'h72;        memory[15199] <=  8'h63;        memory[15200] <=  8'h74;        memory[15201] <=  8'h72;        memory[15202] <=  8'h63;        memory[15203] <=  8'h61;        memory[15204] <=  8'h74;        memory[15205] <=  8'h72;        memory[15206] <=  8'h63;        memory[15207] <=  8'h61;        memory[15208] <=  8'h74;        memory[15209] <=  8'h63;        memory[15210] <=  8'h62;        memory[15211] <=  8'h61;        memory[15212] <=  8'h74;        memory[15213] <=  8'h62;        memory[15214] <=  8'h72;        memory[15215] <=  8'h63;        memory[15216] <=  8'h61;        memory[15217] <=  8'h74;        memory[15218] <=  8'h72;        memory[15219] <=  8'h6e;        memory[15220] <=  8'h62;        memory[15221] <=  8'h61;        memory[15222] <=  8'h63;        memory[15223] <=  8'h61;        memory[15224] <=  8'h74;        memory[15225] <=  8'h79;        memory[15226] <=  8'h73;        memory[15227] <=  8'h6e;        memory[15228] <=  8'h63;        memory[15229] <=  8'h74;        memory[15230] <=  8'h61;        memory[15231] <=  8'h6e;        memory[15232] <=  8'h62;        memory[15233] <=  8'h61;        memory[15234] <=  8'h63;        memory[15235] <=  8'h72;        memory[15236] <=  8'h6e;        memory[15237] <=  8'h74;        memory[15238] <=  8'h61;        memory[15239] <=  8'h62;        memory[15240] <=  8'h74;        memory[15241] <=  8'h6e;        memory[15242] <=  8'h61;        memory[15243] <=  8'h72;        memory[15244] <=  8'h62;        memory[15245] <=  8'h78;        memory[15246] <=  8'h74;        memory[15247] <=  8'h61;        memory[15248] <=  8'h72;        memory[15249] <=  8'h62;        memory[15250] <=  8'h61;        memory[15251] <=  8'h72;        memory[15252] <=  8'h74;        memory[15253] <=  8'h74;        memory[15254] <=  8'h62;        memory[15255] <=  8'h61;        memory[15256] <=  8'h72;        memory[15257] <=  8'h74;        memory[15258] <=  8'h78;        memory[15259] <=  8'h61;        memory[15260] <=  8'h74;        memory[15261] <=  8'h6b;        memory[15262] <=  8'h73;        memory[15263] <=  8'h68;        memory[15264] <=  8'h63;        memory[15265] <=  8'h66;        memory[15266] <=  8'h69;        memory[15267] <=  8'h77;        memory[15268] <=  8'h68;        memory[15269] <=  8'h61;        memory[15270] <=  8'h74;        memory[15271] <=  8'h61;        memory[15272] <=  8'h6e;        memory[15273] <=  8'h61;        memory[15274] <=  8'h62;        memory[15275] <=  8'h61;        memory[15276] <=  8'h63;        memory[15277] <=  8'h61;        memory[15278] <=  8'h74;        memory[15279] <=  8'h61;        memory[15280] <=  8'h62;        memory[15281] <=  8'h61;        memory[15282] <=  8'h72;        memory[15283] <=  8'h63;        memory[15284] <=  8'h61;        memory[15285] <=  8'h68;        memory[15286] <=  8'h64;        memory[15287] <=  8'h75;        memory[15288] <=  8'h63;        memory[15289] <=  8'h74;        memory[15290] <=  8'h61;        memory[15291] <=  8'h64;        memory[15292] <=  8'h61;        memory[15293] <=  8'h61;        memory[15294] <=  8'h63;        memory[15295] <=  8'h61;        memory[15296] <=  8'h72;        memory[15297] <=  8'h63;        memory[15298] <=  8'h74;        memory[15299] <=  8'h72;        memory[15300] <=  8'h63;        memory[15301] <=  8'h61;        memory[15302] <=  8'h74;        memory[15303] <=  8'h72;        memory[15304] <=  8'h63;        memory[15305] <=  8'h61;        memory[15306] <=  8'h74;        memory[15307] <=  8'h63;        memory[15308] <=  8'h62;        memory[15309] <=  8'h61;        memory[15310] <=  8'h74;        memory[15311] <=  8'h62;        memory[15312] <=  8'h72;        memory[15313] <=  8'h63;        memory[15314] <=  8'h61;        memory[15315] <=  8'h74;        memory[15316] <=  8'h72;        memory[15317] <=  8'h6e;        memory[15318] <=  8'h62;        memory[15319] <=  8'h61;        memory[15320] <=  8'h63;        memory[15321] <=  8'h61;        memory[15322] <=  8'h74;        memory[15323] <=  8'h79;        memory[15324] <=  8'h73;        memory[15325] <=  8'h6e;        memory[15326] <=  8'h63;        memory[15327] <=  8'h74;        memory[15328] <=  8'h61;        memory[15329] <=  8'h6e;        memory[15330] <=  8'h62;        memory[15331] <=  8'h61;        memory[15332] <=  8'h63;        memory[15333] <=  8'h72;        memory[15334] <=  8'h6e;        memory[15335] <=  8'h74;        memory[15336] <=  8'h61;        memory[15337] <=  8'h62;        memory[15338] <=  8'h74;        memory[15339] <=  8'h6e;        memory[15340] <=  8'h61;        memory[15341] <=  8'h72;        memory[15342] <=  8'h62;        memory[15343] <=  8'h78;        memory[15344] <=  8'h74;        memory[15345] <=  8'h61;        memory[15346] <=  8'h72;        memory[15347] <=  8'h62;        memory[15348] <=  8'h61;        memory[15349] <=  8'h72;        memory[15350] <=  8'h74;        memory[15351] <=  8'h74;        memory[15352] <=  8'h62;        memory[15353] <=  8'h61;        memory[15354] <=  8'h72;        memory[15355] <=  8'h74;        memory[15356] <=  8'h78;        memory[15357] <=  8'h61;        memory[15358] <=  8'h74;        memory[15359] <=  8'h6b;        memory[15360] <=  8'h73;        memory[15361] <=  8'h68;        memory[15362] <=  8'h63;        memory[15363] <=  8'h66;        memory[15364] <=  8'h69;        memory[15365] <=  8'h77;        memory[15366] <=  8'h68;        memory[15367] <=  8'h61;        memory[15368] <=  8'h74;        memory[15369] <=  8'h61;        memory[15370] <=  8'h6e;        memory[15371] <=  8'h61;        memory[15372] <=  8'h62;        memory[15373] <=  8'h61;        memory[15374] <=  8'h63;        memory[15375] <=  8'h61;        memory[15376] <=  8'h74;        memory[15377] <=  8'h61;        memory[15378] <=  8'h62;        memory[15379] <=  8'h61;        memory[15380] <=  8'h72;        memory[15381] <=  8'h63;        memory[15382] <=  8'h61;        memory[15383] <=  8'h68;        memory[15384] <=  8'h64;        memory[15385] <=  8'h75;        memory[15386] <=  8'h63;        memory[15387] <=  8'h74;        memory[15388] <=  8'h61;        memory[15389] <=  8'h64;        memory[15390] <=  8'h61;        memory[15391] <=  8'h61;        memory[15392] <=  8'h63;        memory[15393] <=  8'h61;        memory[15394] <=  8'h72;        memory[15395] <=  8'h63;        memory[15396] <=  8'h74;        memory[15397] <=  8'h72;        memory[15398] <=  8'h63;        memory[15399] <=  8'h61;        memory[15400] <=  8'h74;        memory[15401] <=  8'h72;        memory[15402] <=  8'h63;        memory[15403] <=  8'h61;        memory[15404] <=  8'h74;        memory[15405] <=  8'h63;        memory[15406] <=  8'h62;        memory[15407] <=  8'h61;        memory[15408] <=  8'h74;        memory[15409] <=  8'h62;        memory[15410] <=  8'h72;        memory[15411] <=  8'h63;        memory[15412] <=  8'h61;        memory[15413] <=  8'h74;        memory[15414] <=  8'h72;        memory[15415] <=  8'h6e;        memory[15416] <=  8'h62;        memory[15417] <=  8'h61;        memory[15418] <=  8'h63;        memory[15419] <=  8'h61;        memory[15420] <=  8'h74;        memory[15421] <=  8'h79;        memory[15422] <=  8'h73;        memory[15423] <=  8'h6e;        memory[15424] <=  8'h63;        memory[15425] <=  8'h74;        memory[15426] <=  8'h61;        memory[15427] <=  8'h6e;        memory[15428] <=  8'h62;        memory[15429] <=  8'h61;        memory[15430] <=  8'h63;        memory[15431] <=  8'h72;        memory[15432] <=  8'h6e;        memory[15433] <=  8'h74;        memory[15434] <=  8'h61;        memory[15435] <=  8'h62;        memory[15436] <=  8'h74;        memory[15437] <=  8'h6e;        memory[15438] <=  8'h61;        memory[15439] <=  8'h72;        memory[15440] <=  8'h62;        memory[15441] <=  8'h78;        memory[15442] <=  8'h74;        memory[15443] <=  8'h61;        memory[15444] <=  8'h72;        memory[15445] <=  8'h5d;        memory[15446] <=  8'h5d;        memory[15447] <=  8'h65;        memory[15448] <=  8'h66;        memory[15449] <=  8'h77;        memory[15450] <=  8'h65;        memory[15451] <=  8'h5d;        memory[15452] <=  8'h65;        memory[15453] <=  8'h67;        memory[15454] <=  8'h73;        memory[15455] <=  8'h67;        memory[15456] <=  8'h66;        memory[15457] <=  8'h62;        memory[15458] <=  8'h61;        memory[15459] <=  8'h72;        memory[15460] <=  8'h74;        memory[15461] <=  8'h74;        memory[15462] <=  8'h62;        memory[15463] <=  8'h61;        memory[15464] <=  8'h72;        memory[15465] <=  8'h74;        memory[15466] <=  8'h78;        memory[15467] <=  8'h61;        memory[15468] <=  8'h74;        memory[15469] <=  8'h6b;        memory[15470] <=  8'h73;        memory[15471] <=  8'h68;        memory[15472] <=  8'h63;        memory[15473] <=  8'h66;        memory[15474] <=  8'h69;        memory[15475] <=  8'h77;        memory[15476] <=  8'h68;        memory[15477] <=  8'h61;        memory[15478] <=  8'h74;        memory[15479] <=  8'h61;        memory[15480] <=  8'h6e;        memory[15481] <=  8'h61;        memory[15482] <=  8'h62;        memory[15483] <=  8'h61;        memory[15484] <=  8'h63;        memory[15485] <=  8'h61;        memory[15486] <=  8'h74;        memory[15487] <=  8'h61;        memory[15488] <=  8'h62;        memory[15489] <=  8'h61;        memory[15490] <=  8'h72;        memory[15491] <=  8'h63;        memory[15492] <=  8'h61;        memory[15493] <=  8'h68;        memory[15494] <=  8'h64;        memory[15495] <=  8'h75;        memory[15496] <=  8'h63;        memory[15497] <=  8'h74;        memory[15498] <=  8'h61;        memory[15499] <=  8'h64;        memory[15500] <=  8'h61;        memory[15501] <=  8'h61;        memory[15502] <=  8'h63;        memory[15503] <=  8'h61;        memory[15504] <=  8'h72;        memory[15505] <=  8'h63;        memory[15506] <=  8'h74;        memory[15507] <=  8'h72;        memory[15508] <=  8'h63;        memory[15509] <=  8'h61;        memory[15510] <=  8'h74;        memory[15511] <=  8'h72;        memory[15512] <=  8'h63;        memory[15513] <=  8'h61;        memory[15514] <=  8'h74;        memory[15515] <=  8'h63;        memory[15516] <=  8'h62;        memory[15517] <=  8'h61;        memory[15518] <=  8'h74;        memory[15519] <=  8'h62;        memory[15520] <=  8'h72;        memory[15521] <=  8'h63;        memory[15522] <=  8'h61;        memory[15523] <=  8'h74;        memory[15524] <=  8'h72;        memory[15525] <=  8'h6e;        memory[15526] <=  8'h62;        memory[15527] <=  8'h61;        memory[15528] <=  8'h63;        memory[15529] <=  8'h61;        memory[15530] <=  8'h74;        memory[15531] <=  8'h79;        memory[15532] <=  8'h73;        memory[15533] <=  8'h6e;        memory[15534] <=  8'h63;        memory[15535] <=  8'h74;        memory[15536] <=  8'h61;        memory[15537] <=  8'h6e;        memory[15538] <=  8'h62;        memory[15539] <=  8'h61;        memory[15540] <=  8'h63;        memory[15541] <=  8'h72;        memory[15542] <=  8'h6e;        memory[15543] <=  8'h74;        memory[15544] <=  8'h61;        memory[15545] <=  8'h62;        memory[15546] <=  8'h74;        memory[15547] <=  8'h6e;        memory[15548] <=  8'h61;        memory[15549] <=  8'h72;        memory[15550] <=  8'h62;        memory[15551] <=  8'h78;        memory[15552] <=  8'h74;        memory[15553] <=  8'h61;        memory[15554] <=  8'h72;        memory[15555] <=  8'h62;        memory[15556] <=  8'h61;        memory[15557] <=  8'h72;        memory[15558] <=  8'h74;        memory[15559] <=  8'h74;        memory[15560] <=  8'h62;        memory[15561] <=  8'h61;        memory[15562] <=  8'h72;        memory[15563] <=  8'h74;        memory[15564] <=  8'h78;        memory[15565] <=  8'h61;        memory[15566] <=  8'h74;        memory[15567] <=  8'h6b;        memory[15568] <=  8'h73;        memory[15569] <=  8'h68;        memory[15570] <=  8'h63;        memory[15571] <=  8'h66;        memory[15572] <=  8'h69;        memory[15573] <=  8'h77;        memory[15574] <=  8'h68;        memory[15575] <=  8'h61;        memory[15576] <=  8'h74;        memory[15577] <=  8'h61;        memory[15578] <=  8'h6e;        memory[15579] <=  8'h61;        memory[15580] <=  8'h62;        memory[15581] <=  8'h61;        memory[15582] <=  8'h63;        memory[15583] <=  8'h61;        memory[15584] <=  8'h74;        memory[15585] <=  8'h61;        memory[15586] <=  8'h62;        memory[15587] <=  8'h61;        memory[15588] <=  8'h72;        memory[15589] <=  8'h63;        memory[15590] <=  8'h61;        memory[15591] <=  8'h68;        memory[15592] <=  8'h64;        memory[15593] <=  8'h75;        memory[15594] <=  8'h63;        memory[15595] <=  8'h74;        memory[15596] <=  8'h61;        memory[15597] <=  8'h64;        memory[15598] <=  8'h61;        memory[15599] <=  8'h61;        memory[15600] <=  8'h63;        memory[15601] <=  8'h61;        memory[15602] <=  8'h72;        memory[15603] <=  8'h63;        memory[15604] <=  8'h74;        memory[15605] <=  8'h72;        memory[15606] <=  8'h63;        memory[15607] <=  8'h61;        memory[15608] <=  8'h74;        memory[15609] <=  8'h72;        memory[15610] <=  8'h63;        memory[15611] <=  8'h61;        memory[15612] <=  8'h74;        memory[15613] <=  8'h63;        memory[15614] <=  8'h62;        memory[15615] <=  8'h61;        memory[15616] <=  8'h74;        memory[15617] <=  8'h62;        memory[15618] <=  8'h72;        memory[15619] <=  8'h63;        memory[15620] <=  8'h61;        memory[15621] <=  8'h74;        memory[15622] <=  8'h72;        memory[15623] <=  8'h6e;        memory[15624] <=  8'h62;        memory[15625] <=  8'h61;        memory[15626] <=  8'h63;        memory[15627] <=  8'h61;        memory[15628] <=  8'h74;        memory[15629] <=  8'h79;        memory[15630] <=  8'h73;        memory[15631] <=  8'h6e;        memory[15632] <=  8'h63;        memory[15633] <=  8'h74;        memory[15634] <=  8'h61;        memory[15635] <=  8'h6e;        memory[15636] <=  8'h62;        memory[15637] <=  8'h61;        memory[15638] <=  8'h63;        memory[15639] <=  8'h72;        memory[15640] <=  8'h6e;        memory[15641] <=  8'h74;        memory[15642] <=  8'h61;        memory[15643] <=  8'h62;        memory[15644] <=  8'h74;        memory[15645] <=  8'h6e;        memory[15646] <=  8'h61;        memory[15647] <=  8'h72;        memory[15648] <=  8'h62;        memory[15649] <=  8'h78;        memory[15650] <=  8'h74;        memory[15651] <=  8'h61;        memory[15652] <=  8'h72;        memory[15653] <=  8'h64;        memory[15654] <=  8'h66;        memory[15655] <=  8'h73;        memory[15656] <=  8'h67;        memory[15657] <=  8'h76;        memory[15658] <=  8'h68;        memory[15659] <=  8'h62;        memory[15660] <=  8'h6b;        memory[15661] <=  8'h6a;        memory[15662] <=  8'h6e;        memory[15663] <=  8'h6d;        memory[15664] <=  8'h62;        memory[15665] <=  8'h76;        memory[15666] <=  8'h78;        memory[15667] <=  8'h63;        memory[15668] <=  8'h73;        memory[15669] <=  8'h66;        memory[15670] <=  8'h72;        memory[15671] <=  8'h74;        memory[15672] <=  8'h79;        memory[15673] <=  8'h75;        memory[15674] <=  8'h6a;        memory[15675] <=  8'h6e;        memory[15676] <=  8'h62;        memory[15677] <=  8'h76;        memory[15678] <=  8'h63;        memory[15679] <=  8'h64;        memory[15680] <=  8'h74;        memory[15681] <=  8'h79;        memory[15682] <=  8'h75;        memory[15683] <=  8'h69;        memory[15684] <=  8'h6b;        memory[15685] <=  8'h6d;        memory[15686] <=  8'h6e;        memory[15687] <=  8'h62;        memory[15688] <=  8'h76;        memory[15689] <=  8'h63;        memory[15690] <=  8'h78;        memory[15691] <=  8'h73;        memory[15692] <=  8'h64;        memory[15693] <=  8'h72;        memory[15694] <=  8'h74;        memory[15695] <=  8'h79;        memory[15696] <=  8'h75;        memory[15697] <=  8'h69;        memory[15698] <=  8'h6b;        memory[15699] <=  8'h6d;        memory[15700] <=  8'h6e;        memory[15701] <=  8'h62;        memory[15702] <=  8'h76;        memory[15703] <=  8'h63;        memory[15704] <=  8'h73;        memory[15705] <=  8'h77;        memory[15706] <=  8'h33;        memory[15707] <=  8'h34;        memory[15708] <=  8'h35;        memory[15709] <=  8'h36;        memory[15710] <=  8'h37;        memory[15711] <=  8'h38;        memory[15712] <=  8'h69;        memory[15713] <=  8'h6b;        memory[15714] <=  8'h6d;        memory[15715] <=  8'h6e;        memory[15716] <=  8'h62;        memory[15717] <=  8'h76;        memory[15718] <=  8'h63;        memory[15719] <=  8'h64;        memory[15720] <=  8'h65;        memory[15721] <=  8'h72;        memory[15722] <=  8'h36;        memory[15723] <=  8'h37;        memory[15724] <=  8'h38;        memory[15725] <=  8'h69;        memory[15726] <=  8'h6f;        memory[15727] <=  8'h6b;        memory[15728] <=  8'h6a;        memory[15729] <=  8'h6e;        memory[15730] <=  8'h62;        memory[15731] <=  8'h76;        memory[15732] <=  8'h63;        memory[15733] <=  8'h64;        memory[15734] <=  8'h72;        memory[15735] <=  8'h74;        memory[15736] <=  8'h79;        memory[15737] <=  8'h75;        memory[15738] <=  8'h73;        memory[15739] <=  8'h6a;        memory[15740] <=  8'h63;        memory[15741] <=  8'h6e;        memory[15742] <=  8'h62;        memory[15743] <=  8'h64;        memory[15744] <=  8'h66;        memory[15745] <=  8'h73;        memory[15746] <=  8'h74;        memory[15747] <=  8'h79;        memory[15748] <=  8'h75;        memory[15749] <=  8'h61;        memory[15750] <=  8'h69;        memory[15751] <=  8'h6b;        memory[15752] <=  8'h78;        memory[15753] <=  8'h6d;        memory[15754] <=  8'h6e;        memory[15755] <=  8'h73;        memory[15756] <=  8'h6a;        memory[15757] <=  8'h6f;        memory[15758] <=  8'h64;        memory[15759] <=  8'h6c;        memory[15760] <=  8'h63;        memory[15761] <=  8'h78;        memory[15762] <=  8'h62;        memory[15763] <=  8'h61;        memory[15764] <=  8'h72;        memory[15765] <=  8'h74;        memory[15766] <=  8'h78;        memory[15767] <=  8'h61;        memory[15768] <=  8'h74;        memory[15769] <=  8'h6b;        memory[15770] <=  8'h73;        memory[15771] <=  8'h68;        memory[15772] <=  8'h63;        memory[15773] <=  8'h66;        memory[15774] <=  8'h69;        memory[15775] <=  8'h77;        memory[15776] <=  8'h68;        memory[15777] <=  8'h61;        memory[15778] <=  8'h74;        memory[15779] <=  8'h61;        memory[15780] <=  8'h6e;        memory[15781] <=  8'h61;        memory[15782] <=  8'h62;        memory[15783] <=  8'h61;        memory[15784] <=  8'h63;        memory[15785] <=  8'h61;        memory[15786] <=  8'h74;        memory[15787] <=  8'h61;        memory[15788] <=  8'h62;        memory[15789] <=  8'h61;        memory[15790] <=  8'h72;        memory[15791] <=  8'h63;        memory[15792] <=  8'h61;        memory[15793] <=  8'h68;        memory[15794] <=  8'h64;        memory[15795] <=  8'h75;        memory[15796] <=  8'h63;        memory[15797] <=  8'h74;        memory[15798] <=  8'h61;        memory[15799] <=  8'h64;        memory[15800] <=  8'h61;        memory[15801] <=  8'h61;        memory[15802] <=  8'h63;        memory[15803] <=  8'h61;        memory[15804] <=  8'h72;        memory[15805] <=  8'h62;        memory[15806] <=  8'h61;        memory[15807] <=  8'h72;        memory[15808] <=  8'h74;        memory[15809] <=  8'h78;        memory[15810] <=  8'h61;        memory[15811] <=  8'h74;        memory[15812] <=  8'h6b;        memory[15813] <=  8'h73;        memory[15814] <=  8'h68;        memory[15815] <=  8'h63;        memory[15816] <=  8'h66;        memory[15817] <=  8'h69;        memory[15818] <=  8'h77;        memory[15819] <=  8'h68;        memory[15820] <=  8'h61;        memory[15821] <=  8'h74;        memory[15822] <=  8'h61;        memory[15823] <=  8'h6e;        memory[15824] <=  8'h61;        memory[15825] <=  8'h62;        memory[15826] <=  8'h61;        memory[15827] <=  8'h63;        memory[15828] <=  8'h61;        memory[15829] <=  8'h74;        memory[15830] <=  8'h61;        memory[15831] <=  8'h62;        memory[15832] <=  8'h61;        memory[15833] <=  8'h72;        memory[15834] <=  8'h63;        memory[15835] <=  8'h61;        memory[15836] <=  8'h68;        memory[15837] <=  8'h64;        memory[15838] <=  8'h75;        memory[15839] <=  8'h63;        memory[15840] <=  8'h74;        memory[15841] <=  8'h61;        memory[15842] <=  8'h64;        memory[15843] <=  8'h61;        memory[15844] <=  8'h61;        memory[15845] <=  8'h63;        memory[15846] <=  8'h61;        memory[15847] <=  8'h72;        memory[15848] <=  8'h62;        memory[15849] <=  8'h61;        memory[15850] <=  8'h72;        memory[15851] <=  8'h74;        memory[15852] <=  8'h78;        memory[15853] <=  8'h61;        memory[15854] <=  8'h74;        memory[15855] <=  8'h6b;        memory[15856] <=  8'h73;        memory[15857] <=  8'h68;        memory[15858] <=  8'h63;        memory[15859] <=  8'h66;        memory[15860] <=  8'h69;        memory[15861] <=  8'h77;        memory[15862] <=  8'h68;        memory[15863] <=  8'h61;        memory[15864] <=  8'h74;        memory[15865] <=  8'h61;        memory[15866] <=  8'h6e;        memory[15867] <=  8'h61;        memory[15868] <=  8'h62;        memory[15869] <=  8'h61;        memory[15870] <=  8'h63;        memory[15871] <=  8'h61;        memory[15872] <=  8'h74;        memory[15873] <=  8'h61;        memory[15874] <=  8'h62;        memory[15875] <=  8'h61;        memory[15876] <=  8'h72;        memory[15877] <=  8'h63;        memory[15878] <=  8'h61;        memory[15879] <=  8'h68;        memory[15880] <=  8'h64;        memory[15881] <=  8'h75;        memory[15882] <=  8'h63;        memory[15883] <=  8'h74;        memory[15884] <=  8'h61;        memory[15885] <=  8'h64;        memory[15886] <=  8'h61;        memory[15887] <=  8'h61;        memory[15888] <=  8'h63;        memory[15889] <=  8'h61;        memory[15890] <=  8'h72;        memory[15891] <=  8'h62;        memory[15892] <=  8'h61;        memory[15893] <=  8'h72;        memory[15894] <=  8'h74;        memory[15895] <=  8'h78;        memory[15896] <=  8'h61;        memory[15897] <=  8'h74;        memory[15898] <=  8'h6b;        memory[15899] <=  8'h73;        memory[15900] <=  8'h68;        memory[15901] <=  8'h63;        memory[15902] <=  8'h66;        memory[15903] <=  8'h69;        memory[15904] <=  8'h77;        memory[15905] <=  8'h68;        memory[15906] <=  8'h61;        memory[15907] <=  8'h74;        memory[15908] <=  8'h61;        memory[15909] <=  8'h6e;        memory[15910] <=  8'h61;        memory[15911] <=  8'h62;        memory[15912] <=  8'h61;        memory[15913] <=  8'h63;        memory[15914] <=  8'h61;        memory[15915] <=  8'h74;        memory[15916] <=  8'h61;        memory[15917] <=  8'h62;        memory[15918] <=  8'h61;        memory[15919] <=  8'h72;        memory[15920] <=  8'h63;        memory[15921] <=  8'h61;        memory[15922] <=  8'h68;        memory[15923] <=  8'h64;        memory[15924] <=  8'h75;        memory[15925] <=  8'h63;        memory[15926] <=  8'h74;        memory[15927] <=  8'h61;        memory[15928] <=  8'h64;        memory[15929] <=  8'h61;        memory[15930] <=  8'h61;        memory[15931] <=  8'h63;        memory[15932] <=  8'h61;        memory[15933] <=  8'h72;        memory[15934] <=  8'h62;        memory[15935] <=  8'h61;        memory[15936] <=  8'h72;        memory[15937] <=  8'h74;        memory[15938] <=  8'h78;        memory[15939] <=  8'h61;        memory[15940] <=  8'h74;        memory[15941] <=  8'h6b;        memory[15942] <=  8'h73;        memory[15943] <=  8'h68;        memory[15944] <=  8'h63;        memory[15945] <=  8'h66;        memory[15946] <=  8'h69;        memory[15947] <=  8'h77;        memory[15948] <=  8'h68;        memory[15949] <=  8'h61;        memory[15950] <=  8'h74;        memory[15951] <=  8'h61;        memory[15952] <=  8'h6e;        memory[15953] <=  8'h61;        memory[15954] <=  8'h62;        memory[15955] <=  8'h61;        memory[15956] <=  8'h63;        memory[15957] <=  8'h61;        memory[15958] <=  8'h74;        memory[15959] <=  8'h61;        memory[15960] <=  8'h62;        memory[15961] <=  8'h61;        memory[15962] <=  8'h72;        memory[15963] <=  8'h63;        memory[15964] <=  8'h61;        memory[15965] <=  8'h68;        memory[15966] <=  8'h64;        memory[15967] <=  8'h75;        memory[15968] <=  8'h63;        memory[15969] <=  8'h74;        memory[15970] <=  8'h61;        memory[15971] <=  8'h64;        memory[15972] <=  8'h61;        memory[15973] <=  8'h61;        memory[15974] <=  8'h63;        memory[15975] <=  8'h61;        memory[15976] <=  8'h72;        memory[15977] <=  8'h62;        memory[15978] <=  8'h61;        memory[15979] <=  8'h72;        memory[15980] <=  8'h74;        memory[15981] <=  8'h78;        memory[15982] <=  8'h61;        memory[15983] <=  8'h74;        memory[15984] <=  8'h6b;        memory[15985] <=  8'h73;        memory[15986] <=  8'h68;        memory[15987] <=  8'h63;        memory[15988] <=  8'h66;        memory[15989] <=  8'h69;        memory[15990] <=  8'h77;        memory[15991] <=  8'h68;        memory[15992] <=  8'h61;        memory[15993] <=  8'h74;        memory[15994] <=  8'h61;        memory[15995] <=  8'h6e;        memory[15996] <=  8'h61;        memory[15997] <=  8'h62;        memory[15998] <=  8'h61;        memory[15999] <=  8'h63;        memory[16000] <=  8'h61;        memory[16001] <=  8'h74;        memory[16002] <=  8'h61;        memory[16003] <=  8'h62;        memory[16004] <=  8'h61;        memory[16005] <=  8'h72;        memory[16006] <=  8'h63;        memory[16007] <=  8'h61;        memory[16008] <=  8'h68;        memory[16009] <=  8'h64;        memory[16010] <=  8'h75;        memory[16011] <=  8'h63;        memory[16012] <=  8'h74;        memory[16013] <=  8'h61;        memory[16014] <=  8'h64;        memory[16015] <=  8'h61;        memory[16016] <=  8'h61;        memory[16017] <=  8'h63;        memory[16018] <=  8'h61;        memory[16019] <=  8'h72;        memory[16020] <=  8'h62;        memory[16021] <=  8'h61;        memory[16022] <=  8'h72;        memory[16023] <=  8'h74;        memory[16024] <=  8'h78;        memory[16025] <=  8'h61;        memory[16026] <=  8'h74;        memory[16027] <=  8'h6b;        memory[16028] <=  8'h73;        memory[16029] <=  8'h68;        memory[16030] <=  8'h63;        memory[16031] <=  8'h66;        memory[16032] <=  8'h69;        memory[16033] <=  8'h77;        memory[16034] <=  8'h68;        memory[16035] <=  8'h61;        memory[16036] <=  8'h74;        memory[16037] <=  8'h61;        memory[16038] <=  8'h6e;        memory[16039] <=  8'h61;        memory[16040] <=  8'h62;        memory[16041] <=  8'h61;        memory[16042] <=  8'h63;        memory[16043] <=  8'h61;        memory[16044] <=  8'h74;        memory[16045] <=  8'h61;        memory[16046] <=  8'h62;        memory[16047] <=  8'h61;        memory[16048] <=  8'h72;        memory[16049] <=  8'h63;        memory[16050] <=  8'h61;        memory[16051] <=  8'h68;        memory[16052] <=  8'h64;        memory[16053] <=  8'h75;        memory[16054] <=  8'h63;        memory[16055] <=  8'h74;        memory[16056] <=  8'h61;        memory[16057] <=  8'h64;        memory[16058] <=  8'h61;        memory[16059] <=  8'h61;        memory[16060] <=  8'h63;        memory[16061] <=  8'h61;        memory[16062] <=  8'h72;        memory[16063] <=  8'h62;        memory[16064] <=  8'h61;        memory[16065] <=  8'h72;        memory[16066] <=  8'h74;        memory[16067] <=  8'h78;        memory[16068] <=  8'h61;        memory[16069] <=  8'h74;        memory[16070] <=  8'h6b;        memory[16071] <=  8'h73;        memory[16072] <=  8'h68;        memory[16073] <=  8'h63;        memory[16074] <=  8'h66;        memory[16075] <=  8'h69;        memory[16076] <=  8'h77;        memory[16077] <=  8'h68;        memory[16078] <=  8'h61;        memory[16079] <=  8'h74;        memory[16080] <=  8'h61;        memory[16081] <=  8'h6e;        memory[16082] <=  8'h61;        memory[16083] <=  8'h62;        memory[16084] <=  8'h61;        memory[16085] <=  8'h63;        memory[16086] <=  8'h61;        memory[16087] <=  8'h74;        memory[16088] <=  8'h61;        memory[16089] <=  8'h62;        memory[16090] <=  8'h61;        memory[16091] <=  8'h72;        memory[16092] <=  8'h63;        memory[16093] <=  8'h61;        memory[16094] <=  8'h68;        memory[16095] <=  8'h64;        memory[16096] <=  8'h75;        memory[16097] <=  8'h63;        memory[16098] <=  8'h74;        memory[16099] <=  8'h61;        memory[16100] <=  8'h64;        memory[16101] <=  8'h61;        memory[16102] <=  8'h61;        memory[16103] <=  8'h63;        memory[16104] <=  8'h61;        memory[16105] <=  8'h72;        memory[16106] <=  8'h62;        memory[16107] <=  8'h61;        memory[16108] <=  8'h72;        memory[16109] <=  8'h74;        memory[16110] <=  8'h78;        memory[16111] <=  8'h61;        memory[16112] <=  8'h74;        memory[16113] <=  8'h6b;        memory[16114] <=  8'h73;        memory[16115] <=  8'h68;        memory[16116] <=  8'h63;        memory[16117] <=  8'h66;        memory[16118] <=  8'h69;        memory[16119] <=  8'h77;        memory[16120] <=  8'h68;        memory[16121] <=  8'h61;        memory[16122] <=  8'h74;        memory[16123] <=  8'h61;        memory[16124] <=  8'h6e;        memory[16125] <=  8'h61;        memory[16126] <=  8'h62;        memory[16127] <=  8'h61;        memory[16128] <=  8'h63;        memory[16129] <=  8'h61;        memory[16130] <=  8'h74;        memory[16131] <=  8'h61;        memory[16132] <=  8'h62;        memory[16133] <=  8'h61;        memory[16134] <=  8'h72;        memory[16135] <=  8'h63;        memory[16136] <=  8'h61;        memory[16137] <=  8'h68;        memory[16138] <=  8'h64;        memory[16139] <=  8'h75;        memory[16140] <=  8'h63;        memory[16141] <=  8'h74;        memory[16142] <=  8'h61;        memory[16143] <=  8'h64;        memory[16144] <=  8'h61;        memory[16145] <=  8'h61;        memory[16146] <=  8'h63;        memory[16147] <=  8'h61;        memory[16148] <=  8'h72;        memory[16149] <=  8'h62;        memory[16150] <=  8'h61;        memory[16151] <=  8'h72;        memory[16152] <=  8'h74;        memory[16153] <=  8'h74;        memory[16154] <=  8'h62;        memory[16155] <=  8'h61;        memory[16156] <=  8'h72;        memory[16157] <=  8'h74;        memory[16158] <=  8'h78;        memory[16159] <=  8'h61;        memory[16160] <=  8'h74;        memory[16161] <=  8'h6b;        memory[16162] <=  8'h73;        memory[16163] <=  8'h68;        memory[16164] <=  8'h63;        memory[16165] <=  8'h66;        memory[16166] <=  8'h69;        memory[16167] <=  8'h77;        memory[16168] <=  8'h68;        memory[16169] <=  8'h61;        memory[16170] <=  8'h74;        memory[16171] <=  8'h61;        memory[16172] <=  8'h6e;        memory[16173] <=  8'h61;        memory[16174] <=  8'h62;        memory[16175] <=  8'h61;        memory[16176] <=  8'h63;        memory[16177] <=  8'h61;        memory[16178] <=  8'h74;        memory[16179] <=  8'h61;        memory[16180] <=  8'h62;        memory[16181] <=  8'h61;        memory[16182] <=  8'h72;        memory[16183] <=  8'h63;        memory[16184] <=  8'h61;        memory[16185] <=  8'h68;        memory[16186] <=  8'h64;        memory[16187] <=  8'h75;        memory[16188] <=  8'h63;        memory[16189] <=  8'h74;        memory[16190] <=  8'h61;        memory[16191] <=  8'h64;        memory[16192] <=  8'h61;        memory[16193] <=  8'h61;        memory[16194] <=  8'h63;        memory[16195] <=  8'h61;        memory[16196] <=  8'h72;        memory[16197] <=  8'h63;        memory[16198] <=  8'h74;        memory[16199] <=  8'h72;        memory[16200] <=  8'h63;        memory[16201] <=  8'h61;        memory[16202] <=  8'h74;        memory[16203] <=  8'h72;        memory[16204] <=  8'h63;        memory[16205] <=  8'h61;        memory[16206] <=  8'h74;        memory[16207] <=  8'h63;        memory[16208] <=  8'h62;        memory[16209] <=  8'h61;        memory[16210] <=  8'h74;        memory[16211] <=  8'h62;        memory[16212] <=  8'h72;        memory[16213] <=  8'h63;        memory[16214] <=  8'h61;        memory[16215] <=  8'h72;        memory[16216] <=  8'h62;        memory[16217] <=  8'h78;        memory[16218] <=  8'h74;        memory[16219] <=  8'h61;        memory[16220] <=  8'h72;        memory[16221] <=  8'h64;        memory[16222] <=  8'h66;        memory[16223] <=  8'h73;        memory[16224] <=  8'h67;        memory[16225] <=  8'h76;        memory[16226] <=  8'h68;        memory[16227] <=  8'h62;        memory[16228] <=  8'h6b;        memory[16229] <=  8'h6a;        memory[16230] <=  8'h6e;        memory[16231] <=  8'h6d;        memory[16232] <=  8'h62;        memory[16233] <=  8'h76;        memory[16234] <=  8'h78;        memory[16235] <=  8'h63;        memory[16236] <=  8'h73;        memory[16237] <=  8'h66;        memory[16238] <=  8'h72;        memory[16239] <=  8'h74;        memory[16240] <=  8'h79;        memory[16241] <=  8'h75;        memory[16242] <=  8'h6a;        memory[16243] <=  8'h6e;        memory[16244] <=  8'h62;        memory[16245] <=  8'h76;        memory[16246] <=  8'h63;        memory[16247] <=  8'h64;        memory[16248] <=  8'h74;        memory[16249] <=  8'h79;        memory[16250] <=  8'h75;        memory[16251] <=  8'h69;        memory[16252] <=  8'h6b;        memory[16253] <=  8'h6d;        memory[16254] <=  8'h6e;        memory[16255] <=  8'h62;        memory[16256] <=  8'h76;        memory[16257] <=  8'h63;        memory[16258] <=  8'h78;        memory[16259] <=  8'h73;        memory[16260] <=  8'h64;        memory[16261] <=  8'h72;        memory[16262] <=  8'h74;        memory[16263] <=  8'h79;        memory[16264] <=  8'h75;        memory[16265] <=  8'h69;        memory[16266] <=  8'h6b;        memory[16267] <=  8'h6d;        memory[16268] <=  8'h6e;        memory[16269] <=  8'h62;        memory[16270] <=  8'h76;        memory[16271] <=  8'h63;        memory[16272] <=  8'h73;        memory[16273] <=  8'h77;        memory[16274] <=  8'h33;        memory[16275] <=  8'h34;        memory[16276] <=  8'h35;        memory[16277] <=  8'h36;        memory[16278] <=  8'h37;        memory[16279] <=  8'h38;        memory[16280] <=  8'h69;        memory[16281] <=  8'h6b;        memory[16282] <=  8'h6d;        memory[16283] <=  8'h6e;        memory[16284] <=  8'h62;        memory[16285] <=  8'h76;        memory[16286] <=  8'h63;        memory[16287] <=  8'h64;        memory[16288] <=  8'h65;        memory[16289] <=  8'h72;        memory[16290] <=  8'h36;        memory[16291] <=  8'h37;        memory[16292] <=  8'h38;        memory[16293] <=  8'h69;        memory[16294] <=  8'h6f;        memory[16295] <=  8'h6b;        memory[16296] <=  8'h6a;        memory[16297] <=  8'h6e;        memory[16298] <=  8'h62;        memory[16299] <=  8'h76;        memory[16300] <=  8'h63;        memory[16301] <=  8'h64;        memory[16302] <=  8'h72;        memory[16303] <=  8'h74;        memory[16304] <=  8'h79;        memory[16305] <=  8'h75;        memory[16306] <=  8'h73;        memory[16307] <=  8'h6a;        memory[16308] <=  8'h63;        memory[16309] <=  8'h6e;        memory[16310] <=  8'h62;        memory[16311] <=  8'h64;        memory[16312] <=  8'h66;        memory[16313] <=  8'h73;        memory[16314] <=  8'h74;        memory[16315] <=  8'h79;        memory[16316] <=  8'h75;        memory[16317] <=  8'h61;        memory[16318] <=  8'h69;        memory[16319] <=  8'h6b;        memory[16320] <=  8'h78;        memory[16321] <=  8'h6d;        memory[16322] <=  8'h6e;        memory[16323] <=  8'h73;        memory[16324] <=  8'h6a;        memory[16325] <=  8'h6f;        memory[16326] <=  8'h64;        memory[16327] <=  8'h6c;        memory[16328] <=  8'h63;        memory[16329] <=  8'h78;        memory[16330] <=  8'h2c;        memory[16331] <=  8'h6d;        memory[16332] <=  8'h73;        memory[16333] <=  8'h6b;        memory[16334] <=  8'h64;        memory[16335] <=  8'h6c;        memory[16336] <=  8'h70;        memory[16337] <=  8'h5b;        memory[16338] <=  8'h3b;        memory[16339] <=  8'h73;        memory[16340] <=  8'h6c;        memory[16341] <=  8'h64;        memory[16342] <=  8'h70;        memory[16343] <=  8'h76;        memory[16344] <=  8'h63;        memory[16345] <=  8'h5b;        memory[16346] <=  8'h78;        memory[16347] <=  8'h76;        memory[16348] <=  8'h63;        memory[16349] <=  8'h5b;        memory[16350] <=  8'h78;        memory[16351] <=  8'h70;        memory[16352] <=  8'h6f;        memory[16353] <=  8'h20;        memory[16354] <=  8'h62;        memory[16355] <=  8'h61;        memory[16356] <=  8'h72;        memory[16357] <=  8'h74;        memory[16358] <=  8'h74;        memory[16359] <=  8'h62;        memory[16360] <=  8'h61;        memory[16361] <=  8'h72;        memory[16362] <=  8'h74;        memory[16363] <=  8'h78;        memory[16364] <=  8'h61;        memory[16365] <=  8'h74;        memory[16366] <=  8'h6b;        memory[16367] <=  8'h73;        memory[16368] <=  8'h68;        memory[16369] <=  8'h63;        memory[16370] <=  8'h66;        memory[16371] <=  8'h69;        memory[16372] <=  8'h77;        memory[16373] <=  8'h68;        memory[16374] <=  8'h61;        memory[16375] <=  8'h69;        memory[16376] <=  8'h6a;        memory[16377] <=  8'h78;        memory[16378] <=  8'h5d;        memory[16379] <=  8'h65;        memory[16380] <=  8'h6b;        memory[16381] <=  8'h6f;        memory[16382] <=  8'h39;        memory[16383] <=  8'h64;        memory[16384] <=  8'h75;        memory[16385] <=  8'h38;        memory[16386] <=  8'h79;        memory[16387] <=  8'h20;        memory[16388] <=  8'h37;        memory[16389] <=  8'h63;        memory[16390] <=  8'h67;        memory[16391] <=  8'h78;        memory[16392] <=  8'h63;        memory[16393] <=  8'h75;        memory[16394] <=  8'h68;        memory[16395] <=  8'h69;        memory[16396] <=  8'h6a;        memory[16397] <=  8'h77;        memory[16398] <=  8'h69;        memory[16399] <=  8'h64;        memory[16400] <=  8'h66;        memory[16401] <=  8'h68;        memory[16402] <=  8'h75;        memory[16403] <=  8'h76;        memory[16404] <=  8'h64;        memory[16405] <=  8'h62;        memory[16406] <=  8'h66;        memory[16407] <=  8'h6a;        memory[16408] <=  8'h6e;        memory[16409] <=  8'h6b;        memory[16410] <=  8'h6a;        memory[16411] <=  8'h65;        memory[16412] <=  8'h38;        memory[16413] <=  8'h66;        memory[16414] <=  8'h37;        memory[16415] <=  8'h67;        memory[16416] <=  8'h79;        memory[16417] <=  8'h76;        memory[16418] <=  8'h63;        memory[16419] <=  8'h68;        memory[16420] <=  8'h69;        memory[16421] <=  8'h6a;        memory[16422] <=  8'h33;        memory[16423] <=  8'h65;        memory[16424] <=  8'h67;        memory[16425] <=  8'h79;        memory[16426] <=  8'h72;        memory[16427] <=  8'h64;        memory[16428] <=  8'h62;        memory[16429] <=  8'h6e;        memory[16430] <=  8'h63;        memory[16431] <=  8'h7a;        memory[16432] <=  8'h6a;        memory[16433] <=  8'h6f;        memory[16434] <=  8'h66;        memory[16435] <=  8'h78;        memory[16436] <=  8'h6a;        memory[16437] <=  8'h69;        memory[16438] <=  8'h63;        memory[16439] <=  8'h68;        memory[16440] <=  8'h62;        memory[16441] <=  8'h6e;        memory[16442] <=  8'h6d;        memory[16443] <=  8'h63;        memory[16444] <=  8'h73;        memory[16445] <=  8'h6c;        memory[16446] <=  8'h6b;        memory[16447] <=  8'h6a;        memory[16448] <=  8'h69;        memory[16449] <=  8'h68;        memory[16450] <=  8'h76;        memory[16451] <=  8'h75;        memory[16452] <=  8'h69;        memory[16453] <=  8'h64;        memory[16454] <=  8'h68;        memory[16455] <=  8'h75;        memory[16456] <=  8'h67;        memory[16457] <=  8'h79;        memory[16458] <=  8'h62;        memory[16459] <=  8'h68;        memory[16460] <=  8'h65;        memory[16461] <=  8'h6a;        memory[16462] <=  8'h72;        memory[16463] <=  8'h6b;        memory[16464] <=  8'h6a;        memory[16465] <=  8'h6f;        memory[16466] <=  8'h64;        memory[16467] <=  8'h67;        memory[16468] <=  8'h69;        memory[16469] <=  8'h75;        memory[16470] <=  8'h69;        memory[16471] <=  8'h67;        memory[16472] <=  8'h76;        memory[16473] <=  8'h79;        memory[16474] <=  8'h75;        memory[16475] <=  8'h67;        memory[16476] <=  8'h78;        memory[16477] <=  8'h68;        memory[16478] <=  8'h63;        memory[16479] <=  8'h20;        memory[16480] <=  8'h20;        memory[16481] <=  8'h20;        memory[16482] <=  8'h78;        memory[16483] <=  8'h76;        memory[16484] <=  8'h20;        memory[16485] <=  8'h63;        memory[16486] <=  8'h78;        memory[16487] <=  8'h67;        memory[16488] <=  8'h79;        memory[16489] <=  8'h63;        memory[16490] <=  8'h75;        memory[16491] <=  8'h68;        memory[16492] <=  8'h6a;        memory[16493] <=  8'h6b;        memory[16494] <=  8'h61;        memory[16495] <=  8'h6c;        memory[16496] <=  8'h78;        memory[16497] <=  8'h76;        memory[16498] <=  8'h70;        memory[16499] <=  8'h6f;        memory[16500] <=  8'h69;        memory[16501] <=  8'h6a;        memory[16502] <=  8'h69;        memory[16503] <=  8'h68;        memory[16504] <=  8'h6a;        memory[16505] <=  8'h62;        memory[16506] <=  8'h77;        memory[16507] <=  8'h65;        memory[16508] <=  8'h6e;        memory[16509] <=  8'h61;        memory[16510] <=  8'h66;        memory[16511] <=  8'h6d;        memory[16512] <=  8'h64;        memory[16513] <=  8'h6b;        memory[16514] <=  8'h6d;        memory[16515] <=  8'h76;        memory[16516] <=  8'h6c;        memory[16517] <=  8'h63;        memory[16518] <=  8'h6f;        memory[16519] <=  8'h64;        memory[16520] <=  8'h69;        memory[16521] <=  8'h75;        memory[16522] <=  8'h68;        memory[16523] <=  8'h73;        memory[16524] <=  8'h66;        memory[16525] <=  8'h65;        memory[16526] <=  8'h62;        memory[16527] <=  8'h6e;        memory[16528] <=  8'h64;        memory[16529] <=  8'h73;        memory[16530] <=  8'h63;        memory[16531] <=  8'h6b;        memory[16532] <=  8'h20;        memory[16533] <=  8'h78;        memory[16534] <=  8'h6a;        memory[16535] <=  8'h78;        memory[16536] <=  8'h63;        memory[16537] <=  8'h73;        memory[16538] <=  8'h64;        memory[16539] <=  8'h66;        memory[16540] <=  8'h6b;        memory[16541] <=  8'h64;        memory[16542] <=  8'h6e;        memory[16543] <=  8'h6d;        memory[16544] <=  8'h64;        memory[16545] <=  8'h73;        memory[16546] <=  8'h63;        memory[16547] <=  8'h6b;        memory[16548] <=  8'h78;        memory[16549] <=  8'h6c;        memory[16550] <=  8'h6f;        memory[16551] <=  8'h66;        memory[16552] <=  8'h6a;        memory[16553] <=  8'h69;        memory[16554] <=  8'h61;        memory[16555] <=  8'h62;        memory[16556] <=  8'h6e;        memory[16557] <=  8'h20;        memory[16558] <=  8'h78;        memory[16559] <=  8'h6b;        memory[16560] <=  8'h6d;        memory[16561] <=  8'h20;        memory[16562] <=  8'h6f;        memory[16563] <=  8'h63;        memory[16564] <=  8'h76;        memory[16565] <=  8'h73;        memory[16566] <=  8'h64;        memory[16567] <=  8'h69;        memory[16568] <=  8'h66;        memory[16569] <=  8'h68;        memory[16570] <=  8'h65;        memory[16571] <=  8'h71;        memory[16572] <=  8'h6a;        memory[16573] <=  8'h77;        memory[16574] <=  8'h62;        memory[16575] <=  8'h65;        memory[16576] <=  8'h6e;        memory[16577] <=  8'h20;        memory[16578] <=  8'h6d;        memory[16579] <=  8'h64;        memory[16580] <=  8'h73;        memory[16581] <=  8'h6c;        memory[16582] <=  8'h76;        memory[16583] <=  8'h6b;        memory[16584] <=  8'h63;        memory[16585] <=  8'h78;        memory[16586] <=  8'h20;        memory[16587] <=  8'h6f;        memory[16588] <=  8'h78;        memory[16589] <=  8'h69;        memory[16590] <=  8'h63;        memory[16591] <=  8'h6a;        memory[16592] <=  8'h76;        memory[16593] <=  8'h64;        memory[16594] <=  8'h66;        memory[16595] <=  8'h65;        memory[16596] <=  8'h71;        memory[16597] <=  8'h6e;        memory[16598] <=  8'h20;        memory[16599] <=  8'h64;        memory[16600] <=  8'h6d;        memory[16601] <=  8'h73;        memory[16602] <=  8'h6c;        memory[16603] <=  8'h63;        memory[16604] <=  8'h78;        memory[16605] <=  8'h6b;        memory[16606] <=  8'h20;        memory[16607] <=  8'h6f;        memory[16608] <=  8'h78;        memory[16609] <=  8'h63;        memory[16610] <=  8'h76;        memory[16611] <=  8'h6a;        memory[16612] <=  8'h64;        memory[16613] <=  8'h62;        memory[16614] <=  8'h71;        memory[16615] <=  8'h77;        memory[16616] <=  8'h65;        memory[16617] <=  8'h6e;        memory[16618] <=  8'h6d;        memory[16619] <=  8'h64;        memory[16620] <=  8'h6c;        memory[16621] <=  8'h73;        memory[16622] <=  8'h2c;        memory[16623] <=  8'h76;        memory[16624] <=  8'h63;        memory[16625] <=  8'h78;        memory[16626] <=  8'h20;        memory[16627] <=  8'h63;        memory[16628] <=  8'h6f;        memory[16629] <=  8'h69;        memory[16630] <=  8'h76;        memory[16631] <=  8'h68;        memory[16632] <=  8'h73;        memory[16633] <=  8'h64;        memory[16634] <=  8'h62;        memory[16635] <=  8'h71;        memory[16636] <=  8'h77;        memory[16637] <=  8'h65;        memory[16638] <=  8'h6e;        memory[16639] <=  8'h64;        memory[16640] <=  8'h6b;        memory[16641] <=  8'h73;        memory[16642] <=  8'h76;        memory[16643] <=  8'h6f;        memory[16644] <=  8'h63;        memory[16645] <=  8'h20;        memory[16646] <=  8'h76;        memory[16647] <=  8'h69;        memory[16648] <=  8'h75;        memory[16649] <=  8'h69;        memory[16650] <=  8'h68;        memory[16651] <=  8'h63;        memory[16652] <=  8'h78;        memory[16653] <=  8'h69;        memory[16654] <=  8'h6f;        memory[16655] <=  8'h76;        memory[16656] <=  8'h73;        memory[16657] <=  8'h64;        memory[16658] <=  8'h61;        memory[16659] <=  8'h64;        memory[16660] <=  8'h6e;        memory[16661] <=  8'h77;        memory[16662] <=  8'h71;        memory[16663] <=  8'h6b;        memory[16664] <=  8'h6c;        memory[16665] <=  8'h73;        memory[16666] <=  8'h76;        memory[16667] <=  8'h6e;        memory[16668] <=  8'h62;        memory[16669] <=  8'h20;        memory[16670] <=  8'h64;        memory[16671] <=  8'h66;        memory[16672] <=  8'h6a;        memory[16673] <=  8'h6b;        memory[16674] <=  8'h71;        memory[16675] <=  8'h64;        memory[16676] <=  8'h77;        memory[16677] <=  8'h65;        memory[16678] <=  8'h6e;        memory[16679] <=  8'h62;        memory[16680] <=  8'h20;        memory[16681] <=  8'h64;        memory[16682] <=  8'h73;        memory[16683] <=  8'h76;        memory[16684] <=  8'h68;        memory[16685] <=  8'h64;        memory[16686] <=  8'h61;        memory[16687] <=  8'h71;        memory[16688] <=  8'h77;        memory[16689] <=  8'h6a;        memory[16690] <=  8'h65;        memory[16691] <=  8'h6e;        memory[16692] <=  8'h64;        memory[16693] <=  8'h20;        memory[16694] <=  8'h61;        memory[16695] <=  8'h63;        memory[16696] <=  8'h62;        memory[16697] <=  8'h68;        memory[16698] <=  8'h64;        memory[16699] <=  8'h61;        memory[16700] <=  8'h77;        memory[16701] <=  8'h71;        memory[16702] <=  8'h6e;        memory[16703] <=  8'h20;        memory[16704] <=  8'h62;        memory[16705] <=  8'h73;        memory[16706] <=  8'h76;        memory[16707] <=  8'h61;        memory[16708] <=  8'h67;        memory[16709] <=  8'h76;        memory[16710] <=  8'h68;        memory[16711] <=  8'h67;        memory[16712] <=  8'h61;        memory[16713] <=  8'h73;        memory[16714] <=  8'h6a;        memory[16715] <=  8'h6b;        memory[16716] <=  8'h63;        memory[16717] <=  8'h78;        memory[16718] <=  8'h76;        memory[16719] <=  8'h6e;        memory[16720] <=  8'h73;        memory[16721] <=  8'h64;        memory[16722] <=  8'h20;        memory[16723] <=  8'h66;        memory[16724] <=  8'h62;        memory[16725] <=  8'h64;        memory[16726] <=  8'h61;        memory[16727] <=  8'h73;        memory[16728] <=  8'h76;        memory[16729] <=  8'h67;        memory[16730] <=  8'h63;        memory[16731] <=  8'h79;        memory[16732] <=  8'h7a;        memory[16733] <=  8'h78;        memory[16734] <=  8'h79;        memory[16735] <=  8'h75;        memory[16736] <=  8'h20;        memory[16737] <=  8'h69;        memory[16738] <=  8'h6a;        memory[16739] <=  8'h64;        memory[16740] <=  8'h66;        memory[16741] <=  8'h6b;        memory[16742] <=  8'h61;        memory[16743] <=  8'h64;        memory[16744] <=  8'h63;        memory[16745] <=  8'h78;        memory[16746] <=  8'h68;        memory[16747] <=  8'h20;        memory[16748] <=  8'h67;        memory[16749] <=  8'h61;        memory[16750] <=  8'h68;        memory[16751] <=  8'h75;        memory[16752] <=  8'h64;        memory[16753] <=  8'h73;        memory[16754] <=  8'h69;        memory[16755] <=  8'h6a;        memory[16756] <=  8'h61;        memory[16757] <=  8'h6b;        memory[16758] <=  8'h63;        memory[16759] <=  8'h62;        memory[16760] <=  8'h61;        memory[16761] <=  8'h72;        memory[16762] <=  8'h73;        memory[16763] <=  8'h68;        memory[16764] <=  8'h64;        memory[16765] <=  8'h66;        memory[16766] <=  8'h67;        memory[16767] <=  8'h73;        memory[16768] <=  8'h68;        memory[16769] <=  8'h64;        memory[16770] <=  8'h66;        memory[16771] <=  8'h68;        memory[16772] <=  8'h64;        memory[16773] <=  8'h6a;        memory[16774] <=  8'h68;        memory[16775] <=  8'h62;        memory[16776] <=  8'h67;        memory[16777] <=  8'h63;        memory[16778] <=  8'h61;        memory[16779] <=  8'h66;        memory[16780] <=  8'h73;        memory[16781] <=  8'h79;        memory[16782] <=  8'h67;        memory[16783] <=  8'h6b;        memory[16784] <=  8'h75;        memory[16785] <=  8'h64;        memory[16786] <=  8'h68;        memory[16787] <=  8'h62;        memory[16788] <=  8'h77;        memory[16789] <=  8'h76;        memory[16790] <=  8'h67;        memory[16791] <=  8'h61;        memory[16792] <=  8'h66;        memory[16793] <=  8'h64;        memory[16794] <=  8'h74;        memory[16795] <=  8'h75;        memory[16796] <=  8'h66;        memory[16797] <=  8'h79;        memory[16798] <=  8'h67;        memory[16799] <=  8'h69;        memory[16800] <=  8'h75;        memory[16801] <=  8'h68;        memory[16802] <=  8'h6c;        memory[16803] <=  8'h6a;        memory[16804] <=  8'h62;        memory[16805] <=  8'h6b;        memory[16806] <=  8'h68;        memory[16807] <=  8'h76;        memory[16808] <=  8'h67;        memory[16809] <=  8'h63;        memory[16810] <=  8'h66;        memory[16811] <=  8'h78;        memory[16812] <=  8'h64;        memory[16813] <=  8'h74;        memory[16814] <=  8'h75;        memory[16815] <=  8'h79;        memory[16816] <=  8'h69;        memory[16817] <=  8'h75;        memory[16818] <=  8'h68;        memory[16819] <=  8'h6c;        memory[16820] <=  8'h6a;        memory[16821] <=  8'h6b;        memory[16822] <=  8'h67;        memory[16823] <=  8'h6a;        memory[16824] <=  8'h63;        memory[16825] <=  8'h66;        memory[16826] <=  8'h68;        memory[16827] <=  8'h64;        memory[16828] <=  8'h67;        memory[16829] <=  8'h72;        memory[16830] <=  8'h79;        memory[16831] <=  8'h74;        memory[16832] <=  8'h66;        memory[16833] <=  8'h75;        memory[16834] <=  8'h79;        memory[16835] <=  8'h69;        memory[16836] <=  8'h68;        memory[16837] <=  8'h6c;        memory[16838] <=  8'h62;        memory[16839] <=  8'h6d;        memory[16840] <=  8'h76;        memory[16841] <=  8'h6e;        memory[16842] <=  8'h63;        memory[16843] <=  8'h66;        memory[16844] <=  8'h68;        memory[16845] <=  8'h64;        memory[16846] <=  8'h74;        memory[16847] <=  8'h75;        memory[16848] <=  8'h67;        memory[16849] <=  8'h79;        memory[16850] <=  8'h69;        memory[16851] <=  8'h68;        memory[16852] <=  8'h75;        memory[16853] <=  8'h6a;        memory[16854] <=  8'h6c;        memory[16855] <=  8'h62;        memory[16856] <=  8'h6d;        memory[16857] <=  8'h76;        memory[16858] <=  8'h6e;        memory[16859] <=  8'h63;        memory[16860] <=  8'h66;        memory[16861] <=  8'h68;        memory[16862] <=  8'h67;        memory[16863] <=  8'h79;        memory[16864] <=  8'h68;        memory[16865] <=  8'h75;        memory[16866] <=  8'h6a;        memory[16867] <=  8'h6e;        memory[16868] <=  8'h2c;        memory[16869] <=  8'h62;        memory[16870] <=  8'h6e;        memory[16871] <=  8'h6d;        memory[16872] <=  8'h76;        memory[16873] <=  8'h6e;        memory[16874] <=  8'h63;        memory[16875] <=  8'h66;        memory[16876] <=  8'h68;        memory[16877] <=  8'h74;        memory[16878] <=  8'h79;        memory[16879] <=  8'h69;        memory[16880] <=  8'h75;        memory[16881] <=  8'h6c;        memory[16882] <=  8'h6a;        memory[16883] <=  8'h62;        memory[16884] <=  8'h6d;        memory[16885] <=  8'h76;        memory[16886] <=  8'h6e;        memory[16887] <=  8'h63;        memory[16888] <=  8'h66;        memory[16889] <=  8'h74;        memory[16890] <=  8'h75;        memory[16891] <=  8'h79;        memory[16892] <=  8'h69;        memory[16893] <=  8'h68;        memory[16894] <=  8'h6b;        memory[16895] <=  8'h62;        memory[16896] <=  8'h76;        memory[16897] <=  8'h63;        memory[16898] <=  8'h66;        memory[16899] <=  8'h67;        memory[16900] <=  8'h74;        memory[16901] <=  8'h75;        memory[16902] <=  8'h79;        memory[16903] <=  8'h69;        memory[16904] <=  8'h75;        memory[16905] <=  8'h68;        memory[16906] <=  8'h6a;        memory[16907] <=  8'h6b;        memory[16908] <=  8'h62;        memory[16909] <=  8'h76;        memory[16910] <=  8'h63;        memory[16911] <=  8'h66;        memory[16912] <=  8'h74;        memory[16913] <=  8'h75;        memory[16914] <=  8'h79;        memory[16915] <=  8'h69;        memory[16916] <=  8'h75;        memory[16917] <=  8'h6a;        memory[16918] <=  8'h6b;        memory[16919] <=  8'h6e;        memory[16920] <=  8'h62;        memory[16921] <=  8'h76;        memory[16922] <=  8'h67;        memory[16923] <=  8'h66;        memory[16924] <=  8'h74;        memory[16925] <=  8'h79;        memory[16926] <=  8'h75;        memory[16927] <=  8'h75;        memory[16928] <=  8'h69;        memory[16929] <=  8'h6a;        memory[16930] <=  8'h6b;        memory[16931] <=  8'h68;        memory[16932] <=  8'h62;        memory[16933] <=  8'h6a;        memory[16934] <=  8'h67;        memory[16935] <=  8'h68;        memory[16936] <=  8'h66;        memory[16937] <=  8'h79;        memory[16938] <=  8'h74;        memory[16939] <=  8'h79;        memory[16940] <=  8'h69;        memory[16941] <=  8'h75;        memory[16942] <=  8'h64;        memory[16943] <=  8'h6a;        memory[16944] <=  8'h6b;        memory[16945] <=  8'h68;        memory[16946] <=  8'h63;        memory[16947] <=  8'h7a;        memory[16948] <=  8'h67;        memory[16949] <=  8'h68;        memory[16950] <=  8'h74;        memory[16951] <=  8'h75;        memory[16952] <=  8'h79;        memory[16953] <=  8'h69;        memory[16954] <=  8'h61;        memory[16955] <=  8'h73;        memory[16956] <=  8'h75;        memory[16957] <=  8'h6a;        memory[16958] <=  8'h6b;        memory[16959] <=  8'h62;        memory[16960] <=  8'h6e;        memory[16961] <=  8'h61;        memory[16962] <=  8'h76;        memory[16963] <=  8'h63;        memory[16964] <=  8'h66;        memory[16965] <=  8'h68;        memory[16966] <=  8'h75;        memory[16967] <=  8'h61;        memory[16968] <=  8'h73;        memory[16969] <=  8'h79;        memory[16970] <=  8'h64;        memory[16971] <=  8'h75;        memory[16972] <=  8'h69;        memory[16973] <=  8'h6a;        memory[16974] <=  8'h61;        memory[16975] <=  8'h6b;        memory[16976] <=  8'h62;        memory[16977] <=  8'h63;        memory[16978] <=  8'h78;        memory[16979] <=  8'h68;        memory[16980] <=  8'h67;        memory[16981] <=  8'h79;        memory[16982] <=  8'h75;        memory[16983] <=  8'h7a;        memory[16984] <=  8'h63;        memory[16985] <=  8'h61;        memory[16986] <=  8'h73;        memory[16987] <=  8'h69;        memory[16988] <=  8'h75;        memory[16989] <=  8'h6f;        memory[16990] <=  8'h69;        memory[16991] <=  8'h6a;        memory[16992] <=  8'h61;        memory[16993] <=  8'h6c;        memory[16994] <=  8'h63;        memory[16995] <=  8'h78;        memory[16996] <=  8'h62;        memory[16997] <=  8'h63;        memory[16998] <=  8'h20;        memory[16999] <=  8'h6e;        memory[17000] <=  8'h76;        memory[17001] <=  8'h63;        memory[17002] <=  8'h61;        memory[17003] <=  8'h64;        memory[17004] <=  8'h73;        memory[17005] <=  8'h67;        memory[17006] <=  8'h79;        memory[17007] <=  8'h68;        memory[17008] <=  8'h75;        memory[17009] <=  8'h61;        memory[17010] <=  8'h6a;        memory[17011] <=  8'h6b;        memory[17012] <=  8'h78;        memory[17013] <=  8'h62;        memory[17014] <=  8'h20;        memory[17015] <=  8'h6e;        memory[17016] <=  8'h76;        memory[17017] <=  8'h63;        memory[17018] <=  8'h61;        memory[17019] <=  8'h73;        memory[17020] <=  8'h67;        memory[17021] <=  8'h68;        memory[17022] <=  8'h75;        memory[17023] <=  8'h6a;        memory[17024] <=  8'h6c;        memory[17025] <=  8'h6b;        memory[17026] <=  8'h63;        memory[17027] <=  8'h78;        memory[17028] <=  8'h20;        memory[17029] <=  8'h6a;        memory[17030] <=  8'h6b;        memory[17031] <=  8'h68;        memory[17032] <=  8'h61;        memory[17033] <=  8'h73;        memory[17034] <=  8'h76;        memory[17035] <=  8'h64;        memory[17036] <=  8'h6e;        memory[17037] <=  8'h20;        memory[17038] <=  8'h62;        memory[17039] <=  8'h6e;        memory[17040] <=  8'h6d;        memory[17041] <=  8'h6b;        memory[17042] <=  8'h77;        memory[17043] <=  8'h64;        memory[17044] <=  8'h6f;        memory[17045] <=  8'h77;        memory[17046] <=  8'h69;        memory[17047] <=  8'h6f;        memory[17048] <=  8'h75;        memory[17049] <=  8'h69;        memory[17050] <=  8'h68;        memory[17051] <=  8'h62;        memory[17052] <=  8'h6e;        memory[17053] <=  8'h6b;        memory[17054] <=  8'h77;        memory[17055] <=  8'h69;        memory[17056] <=  8'h6f;        memory[17057] <=  8'h75;        memory[17058] <=  8'h71;        memory[17059] <=  8'h69;        memory[17060] <=  8'h79;        memory[17061] <=  8'h67;        memory[17062] <=  8'h6a;        memory[17063] <=  8'h64;        memory[17064] <=  8'h61;        memory[17065] <=  8'h76;        memory[17066] <=  8'h62;        memory[17067] <=  8'h6e;        memory[17068] <=  8'h6b;        memory[17069] <=  8'h6f;        memory[17070] <=  8'h70;        memory[17071] <=  8'h64;        memory[17072] <=  8'h76;        memory[17073] <=  8'h69;        memory[17074] <=  8'h6f;        memory[17075] <=  8'h75;        memory[17076] <=  8'h69;        memory[17077] <=  8'h48;        memory[17078] <=  8'h42;        memory[17079] <=  8'h6b;        memory[17080] <=  8'h64;        memory[17081] <=  8'h6e;        memory[17082] <=  8'h6c;        memory[17083] <=  8'h71;        memory[17084] <=  8'h6b;        memory[17085] <=  8'h6d;        memory[17086] <=  8'h6a;        memory[17087] <=  8'h70;        memory[17088] <=  8'h69;        memory[17089] <=  8'h6f;        memory[17090] <=  8'h68;        memory[17091] <=  8'h65;        memory[17092] <=  8'h66;        memory[17093] <=  8'h75;        memory[17094] <=  8'h67;        memory[17095] <=  8'h69;        memory[17096] <=  8'h73;        memory[17097] <=  8'h61;        memory[17098] <=  8'h62;        memory[17099] <=  8'h64;        memory[17100] <=  8'h6b;        memory[17101] <=  8'h6a;        memory[17102] <=  8'h6b;        memory[17103] <=  8'h6c;        memory[17104] <=  8'h6a;        memory[17105] <=  8'h69;        memory[17106] <=  8'h73;        memory[17107] <=  8'h6f;        memory[17108] <=  8'h71;        memory[17109] <=  8'h68;        memory[17110] <=  8'h77;        memory[17111] <=  8'h67;        memory[17112] <=  8'h69;        memory[17113] <=  8'h79;        memory[17114] <=  8'h6a;        memory[17115] <=  8'h64;        memory[17116] <=  8'h76;        memory[17117] <=  8'h62;        memory[17118] <=  8'h6e;        memory[17119] <=  8'h61;        memory[17120] <=  8'h73;        memory[17121] <=  8'h66;        memory[17122] <=  8'h6c;        memory[17123] <=  8'h6b;        memory[17124] <=  8'h64;        memory[17125] <=  8'h6a;        memory[17126] <=  8'h68;        memory[17127] <=  8'h63;        memory[17128] <=  8'h67;        memory[17129] <=  8'h6a;        memory[17130] <=  8'h76;        memory[17131] <=  8'h73;        memory[17132] <=  8'h64;        memory[17133] <=  8'h62;        memory[17134] <=  8'h62;        memory[17135] <=  8'h61;        memory[17136] <=  8'h72;        memory[17137] <=  8'h62;        memory[17138] <=  8'h62;        memory[17139] <=  8'h73;        memory[17140] <=  8'h62;        memory[17141] <=  8'h67;        memory[17142] <=  8'h73;        memory[17143] <=  8'h66;        memory[17144] <=  8'h67;        memory[17145] <=  8'h61;        memory[17146] <=  8'h68;        memory[17147] <=  8'h66;        memory[17148] <=  8'h73;        memory[17149] <=  8'h68;        memory[17150] <=  8'h61;        memory[17151] <=  8'h66;        memory[17152] <=  8'h73;        memory[17153] <=  8'h66;        memory[17154] <=  8'h68;        memory[17155] <=  8'h61;        memory[17156] <=  8'h69;        memory[17157] <=  8'h64;        memory[17158] <=  8'h75;        memory[17159] <=  8'h67;        memory[17160] <=  8'h64;        memory[17161] <=  8'h77;        memory[17162] <=  8'h62;        memory[17163] <=  8'h61;        memory[17164] <=  8'h62;        memory[17165] <=  8'h72;        memory[17166] <=  8'h62;        memory[17167] <=  8'h61;        memory[17168] <=  8'h62;        memory[17169] <=  8'h62;        memory[17170] <=  8'h74;        memory[17171] <=  8'h62;        memory[17172] <=  8'h62;        memory[17173] <=  8'h62;        memory[17174] <=  8'h62;        memory[17175] <=  8'h62;        memory[17176] <=  8'h62;        memory[17177] <=  8'h62;        memory[17178] <=  8'h62;        memory[17179] <=  8'h61;        memory[17180] <=  8'h62;        memory[17181] <=  8'h62;        memory[17182] <=  8'h72;        memory[17183] <=  8'h74;        memory[17184] <=  8'h62;        memory[17185] <=  8'h62;        memory[17186] <=  8'h61;        memory[17187] <=  8'h62;        memory[17188] <=  8'h72;        memory[17189] <=  8'h62;        memory[17190] <=  8'h74;        memory[17191] <=  8'h62;        memory[17192] <=  8'h62;        memory[17193] <=  8'h62;        memory[17194] <=  8'h63;        memory[17195] <=  8'h61;        memory[17196] <=  8'h72;        memory[17197] <=  8'h74;        memory[17198] <=  8'h73;        memory[17199] <=  8'h62;        memory[17200] <=  8'h61;        memory[17201] <=  8'h72;        memory[17202] <=  8'h74;        memory[17203] <=  8'h74;        memory[17204] <=  8'h62;        memory[17205] <=  8'h61;        memory[17206] <=  8'h72;        memory[17207] <=  8'h74;        memory[17208] <=  8'h78;        memory[17209] <=  8'h61;        memory[17210] <=  8'h74;        memory[17211] <=  8'h6b;        memory[17212] <=  8'h73;        memory[17213] <=  8'h68;        memory[17214] <=  8'h63;        memory[17215] <=  8'h66;        memory[17216] <=  8'h69;        memory[17217] <=  8'h77;        memory[17218] <=  8'h68;        memory[17219] <=  8'h61;        memory[17220] <=  8'h74;        memory[17221] <=  8'h61;        memory[17222] <=  8'h6e;        memory[17223] <=  8'h61;        memory[17224] <=  8'h62;        memory[17225] <=  8'h61;        memory[17226] <=  8'h63;        memory[17227] <=  8'h61;        memory[17228] <=  8'h74;        memory[17229] <=  8'h61;        memory[17230] <=  8'h62;        memory[17231] <=  8'h61;        memory[17232] <=  8'h72;        memory[17233] <=  8'h63;        memory[17234] <=  8'h61;        memory[17235] <=  8'h68;        memory[17236] <=  8'h64;        memory[17237] <=  8'h75;        memory[17238] <=  8'h63;        memory[17239] <=  8'h74;        memory[17240] <=  8'h61;        memory[17241] <=  8'h64;        memory[17242] <=  8'h61;        memory[17243] <=  8'h61;        memory[17244] <=  8'h63;        memory[17245] <=  8'h61;        memory[17246] <=  8'h72;        memory[17247] <=  8'h63;        memory[17248] <=  8'h74;        memory[17249] <=  8'h72;        memory[17250] <=  8'h63;        memory[17251] <=  8'h61;        memory[17252] <=  8'h74;        memory[17253] <=  8'h72;        memory[17254] <=  8'h63;        memory[17255] <=  8'h61;        memory[17256] <=  8'h74;        memory[17257] <=  8'h63;        memory[17258] <=  8'h62;        memory[17259] <=  8'h61;        memory[17260] <=  8'h74;        memory[17261] <=  8'h62;        memory[17262] <=  8'h72;        memory[17263] <=  8'h63;        memory[17264] <=  8'h61;        memory[17265] <=  8'h74;        memory[17266] <=  8'h72;        memory[17267] <=  8'h6e;        memory[17268] <=  8'h62;        memory[17269] <=  8'h61;        memory[17270] <=  8'h63;        memory[17271] <=  8'h61;        memory[17272] <=  8'h74;        memory[17273] <=  8'h79;        memory[17274] <=  8'h73;        memory[17275] <=  8'h6e;        memory[17276] <=  8'h63;        memory[17277] <=  8'h74;        memory[17278] <=  8'h61;        memory[17279] <=  8'h6e;        memory[17280] <=  8'h62;        memory[17281] <=  8'h61;        memory[17282] <=  8'h63;        memory[17283] <=  8'h72;        memory[17284] <=  8'h6e;        memory[17285] <=  8'h74;        memory[17286] <=  8'h61;        memory[17287] <=  8'h62;        memory[17288] <=  8'h74;        memory[17289] <=  8'h6e;        memory[17290] <=  8'h61;        memory[17291] <=  8'h72;        memory[17292] <=  8'h62;        memory[17293] <=  8'h78;        memory[17294] <=  8'h74;        memory[17295] <=  8'h61;        memory[17296] <=  8'h72;        memory[17297] <=  8'h62;        memory[17298] <=  8'h61;        memory[17299] <=  8'h72;        memory[17300] <=  8'h74;        memory[17301] <=  8'h74;        memory[17302] <=  8'h62;        memory[17303] <=  8'h61;        memory[17304] <=  8'h72;        memory[17305] <=  8'h74;        memory[17306] <=  8'h78;        memory[17307] <=  8'h61;        memory[17308] <=  8'h74;        memory[17309] <=  8'h6b;        memory[17310] <=  8'h73;        memory[17311] <=  8'h68;        memory[17312] <=  8'h63;        memory[17313] <=  8'h66;        memory[17314] <=  8'h69;        memory[17315] <=  8'h77;        memory[17316] <=  8'h68;        memory[17317] <=  8'h61;        memory[17318] <=  8'h74;        memory[17319] <=  8'h61;        memory[17320] <=  8'h6e;        memory[17321] <=  8'h61;        memory[17322] <=  8'h62;        memory[17323] <=  8'h61;        memory[17324] <=  8'h63;        memory[17325] <=  8'h61;        memory[17326] <=  8'h74;        memory[17327] <=  8'h61;        memory[17328] <=  8'h62;        memory[17329] <=  8'h61;        memory[17330] <=  8'h72;        memory[17331] <=  8'h63;        memory[17332] <=  8'h61;        memory[17333] <=  8'h68;        memory[17334] <=  8'h64;        memory[17335] <=  8'h75;        memory[17336] <=  8'h63;        memory[17337] <=  8'h74;        memory[17338] <=  8'h61;        memory[17339] <=  8'h64;        memory[17340] <=  8'h61;        memory[17341] <=  8'h61;        memory[17342] <=  8'h63;        memory[17343] <=  8'h61;        memory[17344] <=  8'h72;        memory[17345] <=  8'h63;        memory[17346] <=  8'h74;        memory[17347] <=  8'h72;        memory[17348] <=  8'h63;        memory[17349] <=  8'h61;        memory[17350] <=  8'h74;        memory[17351] <=  8'h72;        memory[17352] <=  8'h63;        memory[17353] <=  8'h61;        memory[17354] <=  8'h74;        memory[17355] <=  8'h63;        memory[17356] <=  8'h62;        memory[17357] <=  8'h61;        memory[17358] <=  8'h74;        memory[17359] <=  8'h62;        memory[17360] <=  8'h72;        memory[17361] <=  8'h63;        memory[17362] <=  8'h61;        memory[17363] <=  8'h74;        memory[17364] <=  8'h72;        memory[17365] <=  8'h6e;        memory[17366] <=  8'h62;        memory[17367] <=  8'h61;        memory[17368] <=  8'h63;        memory[17369] <=  8'h61;        memory[17370] <=  8'h74;        memory[17371] <=  8'h79;        memory[17372] <=  8'h73;        memory[17373] <=  8'h6e;        memory[17374] <=  8'h63;        memory[17375] <=  8'h74;        memory[17376] <=  8'h61;        memory[17377] <=  8'h6e;        memory[17378] <=  8'h62;        memory[17379] <=  8'h61;        memory[17380] <=  8'h63;        memory[17381] <=  8'h72;        memory[17382] <=  8'h6e;        memory[17383] <=  8'h74;        memory[17384] <=  8'h61;        memory[17385] <=  8'h62;        memory[17386] <=  8'h74;        memory[17387] <=  8'h6e;        memory[17388] <=  8'h61;        memory[17389] <=  8'h72;        memory[17390] <=  8'h62;        memory[17391] <=  8'h78;        memory[17392] <=  8'h74;        memory[17393] <=  8'h61;        memory[17394] <=  8'h72;        memory[17395] <=  8'h62;        memory[17396] <=  8'h61;        memory[17397] <=  8'h72;        memory[17398] <=  8'h74;        memory[17399] <=  8'h74;        memory[17400] <=  8'h62;        memory[17401] <=  8'h61;        memory[17402] <=  8'h72;        memory[17403] <=  8'h74;        memory[17404] <=  8'h78;        memory[17405] <=  8'h61;        memory[17406] <=  8'h74;        memory[17407] <=  8'h6b;        memory[17408] <=  8'h73;        memory[17409] <=  8'h68;        memory[17410] <=  8'h63;        memory[17411] <=  8'h66;        memory[17412] <=  8'h69;        memory[17413] <=  8'h77;        memory[17414] <=  8'h68;        memory[17415] <=  8'h61;        memory[17416] <=  8'h74;        memory[17417] <=  8'h61;        memory[17418] <=  8'h6e;        memory[17419] <=  8'h61;        memory[17420] <=  8'h62;        memory[17421] <=  8'h61;        memory[17422] <=  8'h63;        memory[17423] <=  8'h61;        memory[17424] <=  8'h74;        memory[17425] <=  8'h61;        memory[17426] <=  8'h62;        memory[17427] <=  8'h61;        memory[17428] <=  8'h72;        memory[17429] <=  8'h63;        memory[17430] <=  8'h61;        memory[17431] <=  8'h68;        memory[17432] <=  8'h64;        memory[17433] <=  8'h75;        memory[17434] <=  8'h63;        memory[17435] <=  8'h74;        memory[17436] <=  8'h61;        memory[17437] <=  8'h64;        memory[17438] <=  8'h61;        memory[17439] <=  8'h61;        memory[17440] <=  8'h63;        memory[17441] <=  8'h61;        memory[17442] <=  8'h72;        memory[17443] <=  8'h63;        memory[17444] <=  8'h74;        memory[17445] <=  8'h72;        memory[17446] <=  8'h63;        memory[17447] <=  8'h61;        memory[17448] <=  8'h74;        memory[17449] <=  8'h72;        memory[17450] <=  8'h63;        memory[17451] <=  8'h61;        memory[17452] <=  8'h74;        memory[17453] <=  8'h63;        memory[17454] <=  8'h62;        memory[17455] <=  8'h61;        memory[17456] <=  8'h74;        memory[17457] <=  8'h62;        memory[17458] <=  8'h72;        memory[17459] <=  8'h63;        memory[17460] <=  8'h61;        memory[17461] <=  8'h74;        memory[17462] <=  8'h72;        memory[17463] <=  8'h6e;        memory[17464] <=  8'h62;        memory[17465] <=  8'h61;        memory[17466] <=  8'h63;        memory[17467] <=  8'h61;        memory[17468] <=  8'h74;        memory[17469] <=  8'h79;        memory[17470] <=  8'h73;        memory[17471] <=  8'h6e;        memory[17472] <=  8'h63;        memory[17473] <=  8'h74;        memory[17474] <=  8'h61;        memory[17475] <=  8'h6e;        memory[17476] <=  8'h62;        memory[17477] <=  8'h61;        memory[17478] <=  8'h63;        memory[17479] <=  8'h72;        memory[17480] <=  8'h6e;        memory[17481] <=  8'h74;        memory[17482] <=  8'h61;        memory[17483] <=  8'h62;        memory[17484] <=  8'h74;        memory[17485] <=  8'h6e;        memory[17486] <=  8'h61;        memory[17487] <=  8'h72;        memory[17488] <=  8'h62;        memory[17489] <=  8'h78;        memory[17490] <=  8'h74;        memory[17491] <=  8'h61;        memory[17492] <=  8'h72;        memory[17493] <=  8'h5d;        memory[17494] <=  8'h5d;        memory[17495] <=  8'h65;        memory[17496] <=  8'h66;        memory[17497] <=  8'h77;        memory[17498] <=  8'h65;        memory[17499] <=  8'h5d;        memory[17500] <=  8'h65;        memory[17501] <=  8'h67;        memory[17502] <=  8'h73;        memory[17503] <=  8'h67;        memory[17504] <=  8'h66;        memory[17505] <=  8'h62;        memory[17506] <=  8'h61;        memory[17507] <=  8'h72;        memory[17508] <=  8'h74;        memory[17509] <=  8'h74;        memory[17510] <=  8'h62;        memory[17511] <=  8'h61;        memory[17512] <=  8'h72;        memory[17513] <=  8'h74;        memory[17514] <=  8'h78;        memory[17515] <=  8'h61;        memory[17516] <=  8'h74;        memory[17517] <=  8'h6b;        memory[17518] <=  8'h73;        memory[17519] <=  8'h68;        memory[17520] <=  8'h63;        memory[17521] <=  8'h66;        memory[17522] <=  8'h69;        memory[17523] <=  8'h77;        memory[17524] <=  8'h68;        memory[17525] <=  8'h61;        memory[17526] <=  8'h74;        memory[17527] <=  8'h61;        memory[17528] <=  8'h6e;        memory[17529] <=  8'h61;        memory[17530] <=  8'h62;        memory[17531] <=  8'h61;        memory[17532] <=  8'h63;        memory[17533] <=  8'h61;        memory[17534] <=  8'h74;        memory[17535] <=  8'h61;        memory[17536] <=  8'h62;        memory[17537] <=  8'h61;        memory[17538] <=  8'h72;        memory[17539] <=  8'h63;        memory[17540] <=  8'h61;        memory[17541] <=  8'h68;        memory[17542] <=  8'h64;        memory[17543] <=  8'h75;        memory[17544] <=  8'h63;        memory[17545] <=  8'h74;        memory[17546] <=  8'h61;        memory[17547] <=  8'h64;        memory[17548] <=  8'h61;        memory[17549] <=  8'h61;        memory[17550] <=  8'h63;        memory[17551] <=  8'h61;        memory[17552] <=  8'h72;        memory[17553] <=  8'h63;        memory[17554] <=  8'h74;        memory[17555] <=  8'h72;        memory[17556] <=  8'h63;        memory[17557] <=  8'h61;        memory[17558] <=  8'h74;        memory[17559] <=  8'h72;        memory[17560] <=  8'h63;        memory[17561] <=  8'h61;        memory[17562] <=  8'h74;        memory[17563] <=  8'h63;        memory[17564] <=  8'h62;        memory[17565] <=  8'h61;        memory[17566] <=  8'h74;        memory[17567] <=  8'h62;        memory[17568] <=  8'h72;        memory[17569] <=  8'h63;        memory[17570] <=  8'h61;        memory[17571] <=  8'h74;        memory[17572] <=  8'h72;        memory[17573] <=  8'h6e;        memory[17574] <=  8'h62;        memory[17575] <=  8'h61;        memory[17576] <=  8'h63;        memory[17577] <=  8'h61;        memory[17578] <=  8'h74;        memory[17579] <=  8'h79;        memory[17580] <=  8'h73;        memory[17581] <=  8'h6e;        memory[17582] <=  8'h63;        memory[17583] <=  8'h74;        memory[17584] <=  8'h61;        memory[17585] <=  8'h6e;        memory[17586] <=  8'h62;        memory[17587] <=  8'h61;        memory[17588] <=  8'h63;        memory[17589] <=  8'h72;        memory[17590] <=  8'h6e;        memory[17591] <=  8'h74;        memory[17592] <=  8'h61;        memory[17593] <=  8'h62;        memory[17594] <=  8'h74;        memory[17595] <=  8'h6e;        memory[17596] <=  8'h61;        memory[17597] <=  8'h72;        memory[17598] <=  8'h62;        memory[17599] <=  8'h78;        memory[17600] <=  8'h74;        memory[17601] <=  8'h61;        memory[17602] <=  8'h72;        memory[17603] <=  8'h62;        memory[17604] <=  8'h61;        memory[17605] <=  8'h72;        memory[17606] <=  8'h74;        memory[17607] <=  8'h74;        memory[17608] <=  8'h62;        memory[17609] <=  8'h61;        memory[17610] <=  8'h72;        memory[17611] <=  8'h74;        memory[17612] <=  8'h78;        memory[17613] <=  8'h61;        memory[17614] <=  8'h74;        memory[17615] <=  8'h6b;        memory[17616] <=  8'h73;        memory[17617] <=  8'h68;        memory[17618] <=  8'h63;        memory[17619] <=  8'h66;        memory[17620] <=  8'h69;        memory[17621] <=  8'h77;        memory[17622] <=  8'h68;        memory[17623] <=  8'h61;        memory[17624] <=  8'h74;        memory[17625] <=  8'h61;        memory[17626] <=  8'h6e;        memory[17627] <=  8'h61;        memory[17628] <=  8'h62;        memory[17629] <=  8'h61;        memory[17630] <=  8'h63;        memory[17631] <=  8'h61;        memory[17632] <=  8'h74;        memory[17633] <=  8'h61;        memory[17634] <=  8'h62;        memory[17635] <=  8'h61;        memory[17636] <=  8'h72;        memory[17637] <=  8'h63;        memory[17638] <=  8'h61;        memory[17639] <=  8'h68;        memory[17640] <=  8'h64;        memory[17641] <=  8'h75;        memory[17642] <=  8'h63;        memory[17643] <=  8'h74;        memory[17644] <=  8'h61;        memory[17645] <=  8'h64;        memory[17646] <=  8'h61;        memory[17647] <=  8'h61;        memory[17648] <=  8'h63;        memory[17649] <=  8'h61;        memory[17650] <=  8'h72;        memory[17651] <=  8'h63;        memory[17652] <=  8'h74;        memory[17653] <=  8'h72;        memory[17654] <=  8'h63;        memory[17655] <=  8'h61;        memory[17656] <=  8'h74;        memory[17657] <=  8'h72;        memory[17658] <=  8'h63;        memory[17659] <=  8'h61;        memory[17660] <=  8'h74;        memory[17661] <=  8'h63;        memory[17662] <=  8'h62;        memory[17663] <=  8'h61;        memory[17664] <=  8'h74;        memory[17665] <=  8'h62;        memory[17666] <=  8'h72;        memory[17667] <=  8'h63;        memory[17668] <=  8'h61;        memory[17669] <=  8'h74;        memory[17670] <=  8'h72;        memory[17671] <=  8'h6e;        memory[17672] <=  8'h62;        memory[17673] <=  8'h61;        memory[17674] <=  8'h63;        memory[17675] <=  8'h61;        memory[17676] <=  8'h74;        memory[17677] <=  8'h79;        memory[17678] <=  8'h73;        memory[17679] <=  8'h6e;        memory[17680] <=  8'h63;        memory[17681] <=  8'h74;        memory[17682] <=  8'h61;        memory[17683] <=  8'h6e;        memory[17684] <=  8'h62;        memory[17685] <=  8'h61;        memory[17686] <=  8'h63;        memory[17687] <=  8'h72;        memory[17688] <=  8'h6e;        memory[17689] <=  8'h74;        memory[17690] <=  8'h61;        memory[17691] <=  8'h62;        memory[17692] <=  8'h74;        memory[17693] <=  8'h6e;        memory[17694] <=  8'h61;        memory[17695] <=  8'h72;        memory[17696] <=  8'h62;        memory[17697] <=  8'h78;        memory[17698] <=  8'h74;        memory[17699] <=  8'h61;        memory[17700] <=  8'h72;        memory[17701] <=  8'h64;        memory[17702] <=  8'h66;        memory[17703] <=  8'h73;        memory[17704] <=  8'h67;        memory[17705] <=  8'h76;        memory[17706] <=  8'h68;        memory[17707] <=  8'h62;        memory[17708] <=  8'h6b;        memory[17709] <=  8'h6a;        memory[17710] <=  8'h6e;        memory[17711] <=  8'h6d;        memory[17712] <=  8'h62;        memory[17713] <=  8'h76;        memory[17714] <=  8'h78;        memory[17715] <=  8'h63;        memory[17716] <=  8'h73;        memory[17717] <=  8'h66;        memory[17718] <=  8'h72;        memory[17719] <=  8'h74;        memory[17720] <=  8'h79;        memory[17721] <=  8'h75;        memory[17722] <=  8'h6a;        memory[17723] <=  8'h6e;        memory[17724] <=  8'h62;        memory[17725] <=  8'h76;        memory[17726] <=  8'h63;        memory[17727] <=  8'h64;        memory[17728] <=  8'h74;        memory[17729] <=  8'h79;        memory[17730] <=  8'h75;        memory[17731] <=  8'h69;        memory[17732] <=  8'h6b;        memory[17733] <=  8'h6d;        memory[17734] <=  8'h6e;        memory[17735] <=  8'h62;        memory[17736] <=  8'h76;        memory[17737] <=  8'h63;        memory[17738] <=  8'h78;        memory[17739] <=  8'h73;        memory[17740] <=  8'h64;        memory[17741] <=  8'h72;        memory[17742] <=  8'h74;        memory[17743] <=  8'h79;        memory[17744] <=  8'h75;        memory[17745] <=  8'h69;        memory[17746] <=  8'h6b;        memory[17747] <=  8'h6d;        memory[17748] <=  8'h6e;        memory[17749] <=  8'h62;        memory[17750] <=  8'h76;        memory[17751] <=  8'h63;        memory[17752] <=  8'h73;        memory[17753] <=  8'h77;        memory[17754] <=  8'h33;        memory[17755] <=  8'h34;        memory[17756] <=  8'h35;        memory[17757] <=  8'h36;        memory[17758] <=  8'h37;        memory[17759] <=  8'h38;        memory[17760] <=  8'h69;        memory[17761] <=  8'h6b;        memory[17762] <=  8'h6d;        memory[17763] <=  8'h6e;        memory[17764] <=  8'h62;        memory[17765] <=  8'h76;        memory[17766] <=  8'h63;        memory[17767] <=  8'h64;        memory[17768] <=  8'h65;        memory[17769] <=  8'h72;        memory[17770] <=  8'h36;        memory[17771] <=  8'h37;        memory[17772] <=  8'h38;        memory[17773] <=  8'h69;        memory[17774] <=  8'h6f;        memory[17775] <=  8'h6b;        memory[17776] <=  8'h6a;        memory[17777] <=  8'h6e;        memory[17778] <=  8'h62;        memory[17779] <=  8'h76;        memory[17780] <=  8'h63;        memory[17781] <=  8'h64;        memory[17782] <=  8'h72;        memory[17783] <=  8'h74;        memory[17784] <=  8'h79;        memory[17785] <=  8'h75;        memory[17786] <=  8'h73;        memory[17787] <=  8'h6a;        memory[17788] <=  8'h63;        memory[17789] <=  8'h6e;        memory[17790] <=  8'h62;        memory[17791] <=  8'h64;        memory[17792] <=  8'h66;        memory[17793] <=  8'h73;        memory[17794] <=  8'h74;        memory[17795] <=  8'h79;        memory[17796] <=  8'h75;        memory[17797] <=  8'h61;        memory[17798] <=  8'h69;        memory[17799] <=  8'h6b;        memory[17800] <=  8'h78;        memory[17801] <=  8'h6d;        memory[17802] <=  8'h6e;        memory[17803] <=  8'h73;        memory[17804] <=  8'h6a;        memory[17805] <=  8'h6f;        memory[17806] <=  8'h64;        memory[17807] <=  8'h6c;        memory[17808] <=  8'h63;        memory[17809] <=  8'h78;        memory[17810] <=  8'h62;        memory[17811] <=  8'h61;        memory[17812] <=  8'h72;        memory[17813] <=  8'h74;        memory[17814] <=  8'h78;        memory[17815] <=  8'h61;        memory[17816] <=  8'h74;        memory[17817] <=  8'h6b;        memory[17818] <=  8'h73;        memory[17819] <=  8'h68;        memory[17820] <=  8'h63;        memory[17821] <=  8'h66;        memory[17822] <=  8'h69;        memory[17823] <=  8'h77;        memory[17824] <=  8'h68;        memory[17825] <=  8'h61;        memory[17826] <=  8'h74;        memory[17827] <=  8'h61;        memory[17828] <=  8'h6e;        memory[17829] <=  8'h61;        memory[17830] <=  8'h62;        memory[17831] <=  8'h61;        memory[17832] <=  8'h63;        memory[17833] <=  8'h61;        memory[17834] <=  8'h74;        memory[17835] <=  8'h61;        memory[17836] <=  8'h62;        memory[17837] <=  8'h61;        memory[17838] <=  8'h72;        memory[17839] <=  8'h63;        memory[17840] <=  8'h61;        memory[17841] <=  8'h68;        memory[17842] <=  8'h64;        memory[17843] <=  8'h75;        memory[17844] <=  8'h63;        memory[17845] <=  8'h74;        memory[17846] <=  8'h61;        memory[17847] <=  8'h64;        memory[17848] <=  8'h61;        memory[17849] <=  8'h61;        memory[17850] <=  8'h63;        memory[17851] <=  8'h61;        memory[17852] <=  8'h72;        memory[17853] <=  8'h62;        memory[17854] <=  8'h61;        memory[17855] <=  8'h72;        memory[17856] <=  8'h74;        memory[17857] <=  8'h78;        memory[17858] <=  8'h61;        memory[17859] <=  8'h74;        memory[17860] <=  8'h6b;        memory[17861] <=  8'h73;        memory[17862] <=  8'h68;        memory[17863] <=  8'h63;        memory[17864] <=  8'h66;        memory[17865] <=  8'h69;        memory[17866] <=  8'h77;        memory[17867] <=  8'h68;        memory[17868] <=  8'h61;        memory[17869] <=  8'h74;        memory[17870] <=  8'h61;        memory[17871] <=  8'h6e;        memory[17872] <=  8'h61;        memory[17873] <=  8'h62;        memory[17874] <=  8'h61;        memory[17875] <=  8'h63;        memory[17876] <=  8'h61;        memory[17877] <=  8'h74;        memory[17878] <=  8'h61;        memory[17879] <=  8'h62;        memory[17880] <=  8'h61;        memory[17881] <=  8'h72;        memory[17882] <=  8'h63;        memory[17883] <=  8'h61;        memory[17884] <=  8'h68;        memory[17885] <=  8'h64;        memory[17886] <=  8'h75;        memory[17887] <=  8'h63;        memory[17888] <=  8'h74;        memory[17889] <=  8'h61;        memory[17890] <=  8'h64;        memory[17891] <=  8'h61;        memory[17892] <=  8'h61;        memory[17893] <=  8'h63;        memory[17894] <=  8'h61;        memory[17895] <=  8'h72;        memory[17896] <=  8'h62;        memory[17897] <=  8'h61;        memory[17898] <=  8'h72;        memory[17899] <=  8'h74;        memory[17900] <=  8'h78;        memory[17901] <=  8'h61;        memory[17902] <=  8'h74;        memory[17903] <=  8'h6b;        memory[17904] <=  8'h73;        memory[17905] <=  8'h68;        memory[17906] <=  8'h63;        memory[17907] <=  8'h66;        memory[17908] <=  8'h69;        memory[17909] <=  8'h77;        memory[17910] <=  8'h68;        memory[17911] <=  8'h61;        memory[17912] <=  8'h74;        memory[17913] <=  8'h61;        memory[17914] <=  8'h6e;        memory[17915] <=  8'h61;        memory[17916] <=  8'h62;        memory[17917] <=  8'h61;        memory[17918] <=  8'h63;        memory[17919] <=  8'h61;        memory[17920] <=  8'h74;        memory[17921] <=  8'h61;        memory[17922] <=  8'h62;        memory[17923] <=  8'h61;        memory[17924] <=  8'h72;        memory[17925] <=  8'h63;        memory[17926] <=  8'h61;        memory[17927] <=  8'h68;        memory[17928] <=  8'h64;        memory[17929] <=  8'h75;        memory[17930] <=  8'h63;        memory[17931] <=  8'h74;        memory[17932] <=  8'h61;        memory[17933] <=  8'h64;        memory[17934] <=  8'h61;        memory[17935] <=  8'h61;        memory[17936] <=  8'h63;        memory[17937] <=  8'h61;        memory[17938] <=  8'h72;        memory[17939] <=  8'h62;        memory[17940] <=  8'h61;        memory[17941] <=  8'h72;        memory[17942] <=  8'h74;        memory[17943] <=  8'h78;        memory[17944] <=  8'h61;        memory[17945] <=  8'h74;        memory[17946] <=  8'h6b;        memory[17947] <=  8'h73;        memory[17948] <=  8'h68;        memory[17949] <=  8'h63;        memory[17950] <=  8'h66;        memory[17951] <=  8'h69;        memory[17952] <=  8'h77;        memory[17953] <=  8'h68;        memory[17954] <=  8'h61;        memory[17955] <=  8'h74;        memory[17956] <=  8'h61;        memory[17957] <=  8'h6e;        memory[17958] <=  8'h61;        memory[17959] <=  8'h62;        memory[17960] <=  8'h61;        memory[17961] <=  8'h63;        memory[17962] <=  8'h61;        memory[17963] <=  8'h74;        memory[17964] <=  8'h61;        memory[17965] <=  8'h62;        memory[17966] <=  8'h61;        memory[17967] <=  8'h72;        memory[17968] <=  8'h63;        memory[17969] <=  8'h61;        memory[17970] <=  8'h68;        memory[17971] <=  8'h64;        memory[17972] <=  8'h75;        memory[17973] <=  8'h63;        memory[17974] <=  8'h74;        memory[17975] <=  8'h61;        memory[17976] <=  8'h64;        memory[17977] <=  8'h61;        memory[17978] <=  8'h61;        memory[17979] <=  8'h63;        memory[17980] <=  8'h61;        memory[17981] <=  8'h72;        memory[17982] <=  8'h62;        memory[17983] <=  8'h61;        memory[17984] <=  8'h72;        memory[17985] <=  8'h74;        memory[17986] <=  8'h78;        memory[17987] <=  8'h61;        memory[17988] <=  8'h74;        memory[17989] <=  8'h6b;        memory[17990] <=  8'h73;        memory[17991] <=  8'h68;        memory[17992] <=  8'h63;        memory[17993] <=  8'h66;        memory[17994] <=  8'h69;        memory[17995] <=  8'h77;        memory[17996] <=  8'h68;        memory[17997] <=  8'h61;        memory[17998] <=  8'h74;        memory[17999] <=  8'h61;        memory[18000] <=  8'h6e;        memory[18001] <=  8'h61;        memory[18002] <=  8'h62;        memory[18003] <=  8'h61;        memory[18004] <=  8'h63;        memory[18005] <=  8'h61;        memory[18006] <=  8'h74;        memory[18007] <=  8'h61;        memory[18008] <=  8'h62;        memory[18009] <=  8'h61;        memory[18010] <=  8'h72;        memory[18011] <=  8'h63;        memory[18012] <=  8'h61;        memory[18013] <=  8'h68;        memory[18014] <=  8'h64;        memory[18015] <=  8'h75;        memory[18016] <=  8'h63;        memory[18017] <=  8'h74;        memory[18018] <=  8'h61;        memory[18019] <=  8'h64;        memory[18020] <=  8'h61;        memory[18021] <=  8'h61;        memory[18022] <=  8'h63;        memory[18023] <=  8'h61;        memory[18024] <=  8'h72;        memory[18025] <=  8'h62;        memory[18026] <=  8'h61;        memory[18027] <=  8'h72;        memory[18028] <=  8'h74;        memory[18029] <=  8'h78;        memory[18030] <=  8'h61;        memory[18031] <=  8'h74;        memory[18032] <=  8'h6b;        memory[18033] <=  8'h73;        memory[18034] <=  8'h68;        memory[18035] <=  8'h63;        memory[18036] <=  8'h66;        memory[18037] <=  8'h69;        memory[18038] <=  8'h77;        memory[18039] <=  8'h68;        memory[18040] <=  8'h61;        memory[18041] <=  8'h74;        memory[18042] <=  8'h61;        memory[18043] <=  8'h6e;        memory[18044] <=  8'h61;        memory[18045] <=  8'h62;        memory[18046] <=  8'h61;        memory[18047] <=  8'h63;        memory[18048] <=  8'h61;        memory[18049] <=  8'h74;        memory[18050] <=  8'h61;        memory[18051] <=  8'h62;        memory[18052] <=  8'h61;        memory[18053] <=  8'h72;        memory[18054] <=  8'h63;        memory[18055] <=  8'h61;        memory[18056] <=  8'h68;        memory[18057] <=  8'h64;        memory[18058] <=  8'h75;        memory[18059] <=  8'h63;        memory[18060] <=  8'h74;        memory[18061] <=  8'h61;        memory[18062] <=  8'h64;        memory[18063] <=  8'h61;        memory[18064] <=  8'h61;        memory[18065] <=  8'h63;        memory[18066] <=  8'h61;        memory[18067] <=  8'h72;        memory[18068] <=  8'h62;        memory[18069] <=  8'h61;        memory[18070] <=  8'h72;        memory[18071] <=  8'h74;        memory[18072] <=  8'h78;        memory[18073] <=  8'h61;        memory[18074] <=  8'h74;        memory[18075] <=  8'h6b;        memory[18076] <=  8'h73;        memory[18077] <=  8'h68;        memory[18078] <=  8'h63;        memory[18079] <=  8'h66;        memory[18080] <=  8'h69;        memory[18081] <=  8'h77;        memory[18082] <=  8'h68;        memory[18083] <=  8'h61;        memory[18084] <=  8'h74;        memory[18085] <=  8'h61;        memory[18086] <=  8'h6e;        memory[18087] <=  8'h61;        memory[18088] <=  8'h62;        memory[18089] <=  8'h61;        memory[18090] <=  8'h63;        memory[18091] <=  8'h61;        memory[18092] <=  8'h74;        memory[18093] <=  8'h61;        memory[18094] <=  8'h62;        memory[18095] <=  8'h61;        memory[18096] <=  8'h72;        memory[18097] <=  8'h63;        memory[18098] <=  8'h61;        memory[18099] <=  8'h68;        memory[18100] <=  8'h64;        memory[18101] <=  8'h75;        memory[18102] <=  8'h63;        memory[18103] <=  8'h74;        memory[18104] <=  8'h61;        memory[18105] <=  8'h64;        memory[18106] <=  8'h61;        memory[18107] <=  8'h61;        memory[18108] <=  8'h63;        memory[18109] <=  8'h61;        memory[18110] <=  8'h72;        memory[18111] <=  8'h62;        memory[18112] <=  8'h61;        memory[18113] <=  8'h72;        memory[18114] <=  8'h74;        memory[18115] <=  8'h78;        memory[18116] <=  8'h61;        memory[18117] <=  8'h74;        memory[18118] <=  8'h6b;        memory[18119] <=  8'h73;        memory[18120] <=  8'h68;        memory[18121] <=  8'h63;        memory[18122] <=  8'h66;        memory[18123] <=  8'h69;        memory[18124] <=  8'h77;        memory[18125] <=  8'h68;        memory[18126] <=  8'h61;        memory[18127] <=  8'h74;        memory[18128] <=  8'h61;        memory[18129] <=  8'h6e;        memory[18130] <=  8'h61;        memory[18131] <=  8'h62;        memory[18132] <=  8'h61;        memory[18133] <=  8'h63;        memory[18134] <=  8'h61;        memory[18135] <=  8'h74;        memory[18136] <=  8'h61;        memory[18137] <=  8'h62;        memory[18138] <=  8'h61;        memory[18139] <=  8'h72;        memory[18140] <=  8'h63;        memory[18141] <=  8'h61;        memory[18142] <=  8'h68;        memory[18143] <=  8'h64;        memory[18144] <=  8'h75;        memory[18145] <=  8'h63;        memory[18146] <=  8'h74;        memory[18147] <=  8'h61;        memory[18148] <=  8'h64;        memory[18149] <=  8'h61;        memory[18150] <=  8'h61;        memory[18151] <=  8'h63;        memory[18152] <=  8'h61;        memory[18153] <=  8'h72;        memory[18154] <=  8'h62;        memory[18155] <=  8'h61;        memory[18156] <=  8'h72;        memory[18157] <=  8'h74;        memory[18158] <=  8'h78;        memory[18159] <=  8'h61;        memory[18160] <=  8'h74;        memory[18161] <=  8'h6b;        memory[18162] <=  8'h73;        memory[18163] <=  8'h68;        memory[18164] <=  8'h63;        memory[18165] <=  8'h66;        memory[18166] <=  8'h69;        memory[18167] <=  8'h77;        memory[18168] <=  8'h68;        memory[18169] <=  8'h61;        memory[18170] <=  8'h74;        memory[18171] <=  8'h61;        memory[18172] <=  8'h6e;        memory[18173] <=  8'h61;        memory[18174] <=  8'h62;        memory[18175] <=  8'h61;        memory[18176] <=  8'h63;        memory[18177] <=  8'h61;        memory[18178] <=  8'h74;        memory[18179] <=  8'h61;        memory[18180] <=  8'h62;        memory[18181] <=  8'h61;        memory[18182] <=  8'h72;        memory[18183] <=  8'h63;        memory[18184] <=  8'h61;        memory[18185] <=  8'h68;        memory[18186] <=  8'h64;        memory[18187] <=  8'h75;        memory[18188] <=  8'h63;        memory[18189] <=  8'h74;        memory[18190] <=  8'h61;        memory[18191] <=  8'h64;        memory[18192] <=  8'h61;        memory[18193] <=  8'h61;        memory[18194] <=  8'h63;        memory[18195] <=  8'h61;        memory[18196] <=  8'h72;        memory[18197] <=  8'h62;        memory[18198] <=  8'h61;        memory[18199] <=  8'h72;        memory[18200] <=  8'h74;        memory[18201] <=  8'h74;        memory[18202] <=  8'h62;        memory[18203] <=  8'h61;        memory[18204] <=  8'h72;        memory[18205] <=  8'h74;        memory[18206] <=  8'h78;        memory[18207] <=  8'h61;        memory[18208] <=  8'h74;        memory[18209] <=  8'h6b;        memory[18210] <=  8'h73;        memory[18211] <=  8'h68;        memory[18212] <=  8'h63;        memory[18213] <=  8'h66;        memory[18214] <=  8'h69;        memory[18215] <=  8'h77;        memory[18216] <=  8'h68;        memory[18217] <=  8'h61;        memory[18218] <=  8'h74;        memory[18219] <=  8'h61;        memory[18220] <=  8'h6e;        memory[18221] <=  8'h61;        memory[18222] <=  8'h62;        memory[18223] <=  8'h61;        memory[18224] <=  8'h63;        memory[18225] <=  8'h61;        memory[18226] <=  8'h74;        memory[18227] <=  8'h61;        memory[18228] <=  8'h62;        memory[18229] <=  8'h61;        memory[18230] <=  8'h72;        memory[18231] <=  8'h63;        memory[18232] <=  8'h61;        memory[18233] <=  8'h68;        memory[18234] <=  8'h64;        memory[18235] <=  8'h75;        memory[18236] <=  8'h63;        memory[18237] <=  8'h74;        memory[18238] <=  8'h61;        memory[18239] <=  8'h64;        memory[18240] <=  8'h61;        memory[18241] <=  8'h61;        memory[18242] <=  8'h63;        memory[18243] <=  8'h61;        memory[18244] <=  8'h72;        memory[18245] <=  8'h63;        memory[18246] <=  8'h74;        memory[18247] <=  8'h72;        memory[18248] <=  8'h63;        memory[18249] <=  8'h61;        memory[18250] <=  8'h74;        memory[18251] <=  8'h72;        memory[18252] <=  8'h63;        memory[18253] <=  8'h61;        memory[18254] <=  8'h74;        memory[18255] <=  8'h63;        memory[18256] <=  8'h62;        memory[18257] <=  8'h61;        memory[18258] <=  8'h74;        memory[18259] <=  8'h62;        memory[18260] <=  8'h72;        memory[18261] <=  8'h63;        memory[18262] <=  8'h61;        memory[18263] <=  8'h72;        memory[18264] <=  8'h62;        memory[18265] <=  8'h78;        memory[18266] <=  8'h74;        memory[18267] <=  8'h61;        memory[18268] <=  8'h72;        memory[18269] <=  8'h64;        memory[18270] <=  8'h66;        memory[18271] <=  8'h73;        memory[18272] <=  8'h67;        memory[18273] <=  8'h76;        memory[18274] <=  8'h68;        memory[18275] <=  8'h62;        memory[18276] <=  8'h6b;        memory[18277] <=  8'h6a;        memory[18278] <=  8'h6e;        memory[18279] <=  8'h6d;        memory[18280] <=  8'h62;        memory[18281] <=  8'h76;        memory[18282] <=  8'h78;        memory[18283] <=  8'h63;        memory[18284] <=  8'h73;        memory[18285] <=  8'h66;        memory[18286] <=  8'h72;        memory[18287] <=  8'h74;        memory[18288] <=  8'h79;        memory[18289] <=  8'h75;        memory[18290] <=  8'h6a;        memory[18291] <=  8'h6e;        memory[18292] <=  8'h62;        memory[18293] <=  8'h76;        memory[18294] <=  8'h63;        memory[18295] <=  8'h64;        memory[18296] <=  8'h74;        memory[18297] <=  8'h79;        memory[18298] <=  8'h75;        memory[18299] <=  8'h69;        memory[18300] <=  8'h6b;        memory[18301] <=  8'h6d;        memory[18302] <=  8'h6e;        memory[18303] <=  8'h62;        memory[18304] <=  8'h76;        memory[18305] <=  8'h63;        memory[18306] <=  8'h78;        memory[18307] <=  8'h73;        memory[18308] <=  8'h64;        memory[18309] <=  8'h72;        memory[18310] <=  8'h74;        memory[18311] <=  8'h79;        memory[18312] <=  8'h75;        memory[18313] <=  8'h69;        memory[18314] <=  8'h6b;        memory[18315] <=  8'h6d;        memory[18316] <=  8'h6e;        memory[18317] <=  8'h62;        memory[18318] <=  8'h76;        memory[18319] <=  8'h63;        memory[18320] <=  8'h73;        memory[18321] <=  8'h77;        memory[18322] <=  8'h33;        memory[18323] <=  8'h34;        memory[18324] <=  8'h35;        memory[18325] <=  8'h36;        memory[18326] <=  8'h37;        memory[18327] <=  8'h38;        memory[18328] <=  8'h69;        memory[18329] <=  8'h6b;        memory[18330] <=  8'h6d;        memory[18331] <=  8'h6e;        memory[18332] <=  8'h62;        memory[18333] <=  8'h76;        memory[18334] <=  8'h63;        memory[18335] <=  8'h64;        memory[18336] <=  8'h65;        memory[18337] <=  8'h72;        memory[18338] <=  8'h36;        memory[18339] <=  8'h37;        memory[18340] <=  8'h38;        memory[18341] <=  8'h69;        memory[18342] <=  8'h6f;        memory[18343] <=  8'h6b;        memory[18344] <=  8'h6a;        memory[18345] <=  8'h6e;        memory[18346] <=  8'h62;        memory[18347] <=  8'h76;        memory[18348] <=  8'h63;        memory[18349] <=  8'h64;        memory[18350] <=  8'h72;        memory[18351] <=  8'h74;        memory[18352] <=  8'h79;        memory[18353] <=  8'h75;        memory[18354] <=  8'h73;        memory[18355] <=  8'h6a;        memory[18356] <=  8'h63;        memory[18357] <=  8'h6e;        memory[18358] <=  8'h62;        memory[18359] <=  8'h64;        memory[18360] <=  8'h66;        memory[18361] <=  8'h73;        memory[18362] <=  8'h74;        memory[18363] <=  8'h79;        memory[18364] <=  8'h75;        memory[18365] <=  8'h61;        memory[18366] <=  8'h69;        memory[18367] <=  8'h6b;        memory[18368] <=  8'h78;        memory[18369] <=  8'h6d;        memory[18370] <=  8'h6e;        memory[18371] <=  8'h73;        memory[18372] <=  8'h6a;        memory[18373] <=  8'h6f;        memory[18374] <=  8'h64;        memory[18375] <=  8'h6c;        memory[18376] <=  8'h63;        memory[18377] <=  8'h78;        memory[18378] <=  8'h2c;        memory[18379] <=  8'h6d;        memory[18380] <=  8'h73;        memory[18381] <=  8'h6b;        memory[18382] <=  8'h64;        memory[18383] <=  8'h6c;        memory[18384] <=  8'h70;        memory[18385] <=  8'h5b;        memory[18386] <=  8'h3b;        memory[18387] <=  8'h73;        memory[18388] <=  8'h6c;        memory[18389] <=  8'h64;        memory[18390] <=  8'h70;        memory[18391] <=  8'h76;        memory[18392] <=  8'h63;        memory[18393] <=  8'h5b;        memory[18394] <=  8'h78;        memory[18395] <=  8'h76;        memory[18396] <=  8'h63;        memory[18397] <=  8'h5b;        memory[18398] <=  8'h78;        memory[18399] <=  8'h70;        memory[18400] <=  8'h6f;        memory[18401] <=  8'h20;        memory[18402] <=  8'h62;        memory[18403] <=  8'h61;        memory[18404] <=  8'h72;        memory[18405] <=  8'h74;        memory[18406] <=  8'h74;        memory[18407] <=  8'h62;        memory[18408] <=  8'h61;        memory[18409] <=  8'h72;        memory[18410] <=  8'h74;        memory[18411] <=  8'h78;        memory[18412] <=  8'h61;        memory[18413] <=  8'h74;        memory[18414] <=  8'h6b;        memory[18415] <=  8'h73;        memory[18416] <=  8'h68;        memory[18417] <=  8'h63;        memory[18418] <=  8'h66;        memory[18419] <=  8'h69;        memory[18420] <=  8'h77;        memory[18421] <=  8'h68;        memory[18422] <=  8'h61;        memory[18423] <=  8'h69;        memory[18424] <=  8'h6a;        memory[18425] <=  8'h78;        memory[18426] <=  8'h5d;        memory[18427] <=  8'h65;        memory[18428] <=  8'h6b;        memory[18429] <=  8'h6f;        memory[18430] <=  8'h39;        memory[18431] <=  8'h64;        memory[18432] <=  8'h75;        memory[18433] <=  8'h38;        memory[18434] <=  8'h79;        memory[18435] <=  8'h20;        memory[18436] <=  8'h37;        memory[18437] <=  8'h63;        memory[18438] <=  8'h67;        memory[18439] <=  8'h78;        memory[18440] <=  8'h63;        memory[18441] <=  8'h75;        memory[18442] <=  8'h68;        memory[18443] <=  8'h69;        memory[18444] <=  8'h6a;        memory[18445] <=  8'h77;        memory[18446] <=  8'h69;        memory[18447] <=  8'h64;        memory[18448] <=  8'h66;        memory[18449] <=  8'h68;        memory[18450] <=  8'h75;        memory[18451] <=  8'h76;        memory[18452] <=  8'h64;        memory[18453] <=  8'h62;        memory[18454] <=  8'h66;        memory[18455] <=  8'h6a;        memory[18456] <=  8'h6e;        memory[18457] <=  8'h6b;        memory[18458] <=  8'h6a;        memory[18459] <=  8'h65;        memory[18460] <=  8'h38;        memory[18461] <=  8'h66;        memory[18462] <=  8'h37;        memory[18463] <=  8'h67;        memory[18464] <=  8'h79;        memory[18465] <=  8'h76;        memory[18466] <=  8'h63;        memory[18467] <=  8'h68;        memory[18468] <=  8'h69;        memory[18469] <=  8'h6a;        memory[18470] <=  8'h33;        memory[18471] <=  8'h65;        memory[18472] <=  8'h67;        memory[18473] <=  8'h79;        memory[18474] <=  8'h72;        memory[18475] <=  8'h64;        memory[18476] <=  8'h62;        memory[18477] <=  8'h6e;        memory[18478] <=  8'h63;        memory[18479] <=  8'h7a;        memory[18480] <=  8'h6a;        memory[18481] <=  8'h6f;        memory[18482] <=  8'h66;        memory[18483] <=  8'h78;        memory[18484] <=  8'h6a;        memory[18485] <=  8'h69;        memory[18486] <=  8'h63;        memory[18487] <=  8'h68;        memory[18488] <=  8'h62;        memory[18489] <=  8'h6e;        memory[18490] <=  8'h6d;        memory[18491] <=  8'h63;        memory[18492] <=  8'h73;        memory[18493] <=  8'h6c;        memory[18494] <=  8'h6b;        memory[18495] <=  8'h6a;        memory[18496] <=  8'h69;        memory[18497] <=  8'h68;        memory[18498] <=  8'h76;        memory[18499] <=  8'h75;        memory[18500] <=  8'h69;        memory[18501] <=  8'h64;        memory[18502] <=  8'h68;        memory[18503] <=  8'h75;        memory[18504] <=  8'h67;        memory[18505] <=  8'h79;        memory[18506] <=  8'h62;        memory[18507] <=  8'h68;        memory[18508] <=  8'h65;        memory[18509] <=  8'h6a;        memory[18510] <=  8'h72;        memory[18511] <=  8'h6b;        memory[18512] <=  8'h6a;        memory[18513] <=  8'h6f;        memory[18514] <=  8'h64;        memory[18515] <=  8'h67;        memory[18516] <=  8'h69;        memory[18517] <=  8'h75;        memory[18518] <=  8'h69;        memory[18519] <=  8'h67;        memory[18520] <=  8'h76;        memory[18521] <=  8'h79;        memory[18522] <=  8'h75;        memory[18523] <=  8'h67;        memory[18524] <=  8'h78;        memory[18525] <=  8'h68;        memory[18526] <=  8'h63;        memory[18527] <=  8'h20;        memory[18528] <=  8'h20;        memory[18529] <=  8'h20;        memory[18530] <=  8'h78;        memory[18531] <=  8'h76;        memory[18532] <=  8'h20;        memory[18533] <=  8'h63;        memory[18534] <=  8'h78;        memory[18535] <=  8'h67;        memory[18536] <=  8'h79;        memory[18537] <=  8'h63;        memory[18538] <=  8'h75;        memory[18539] <=  8'h68;        memory[18540] <=  8'h6a;        memory[18541] <=  8'h6b;        memory[18542] <=  8'h61;        memory[18543] <=  8'h6c;        memory[18544] <=  8'h78;        memory[18545] <=  8'h76;        memory[18546] <=  8'h70;        memory[18547] <=  8'h6f;        memory[18548] <=  8'h69;        memory[18549] <=  8'h6a;        memory[18550] <=  8'h69;        memory[18551] <=  8'h68;        memory[18552] <=  8'h6a;        memory[18553] <=  8'h62;        memory[18554] <=  8'h77;        memory[18555] <=  8'h65;        memory[18556] <=  8'h6e;        memory[18557] <=  8'h61;        memory[18558] <=  8'h66;        memory[18559] <=  8'h6d;        memory[18560] <=  8'h64;        memory[18561] <=  8'h6b;        memory[18562] <=  8'h6d;        memory[18563] <=  8'h76;        memory[18564] <=  8'h6c;        memory[18565] <=  8'h63;        memory[18566] <=  8'h6f;        memory[18567] <=  8'h64;        memory[18568] <=  8'h69;        memory[18569] <=  8'h75;        memory[18570] <=  8'h68;        memory[18571] <=  8'h73;        memory[18572] <=  8'h66;        memory[18573] <=  8'h65;        memory[18574] <=  8'h62;        memory[18575] <=  8'h6e;        memory[18576] <=  8'h64;        memory[18577] <=  8'h73;        memory[18578] <=  8'h63;        memory[18579] <=  8'h6b;        memory[18580] <=  8'h20;        memory[18581] <=  8'h78;        memory[18582] <=  8'h6a;        memory[18583] <=  8'h78;        memory[18584] <=  8'h63;        memory[18585] <=  8'h73;        memory[18586] <=  8'h64;        memory[18587] <=  8'h66;        memory[18588] <=  8'h6b;        memory[18589] <=  8'h64;        memory[18590] <=  8'h6e;        memory[18591] <=  8'h6d;        memory[18592] <=  8'h64;        memory[18593] <=  8'h73;        memory[18594] <=  8'h63;        memory[18595] <=  8'h6b;        memory[18596] <=  8'h78;        memory[18597] <=  8'h6c;        memory[18598] <=  8'h6f;        memory[18599] <=  8'h66;        memory[18600] <=  8'h6a;        memory[18601] <=  8'h69;        memory[18602] <=  8'h61;        memory[18603] <=  8'h62;        memory[18604] <=  8'h6e;        memory[18605] <=  8'h20;        memory[18606] <=  8'h78;        memory[18607] <=  8'h6b;        memory[18608] <=  8'h6d;        memory[18609] <=  8'h20;        memory[18610] <=  8'h6f;        memory[18611] <=  8'h63;        memory[18612] <=  8'h76;        memory[18613] <=  8'h73;        memory[18614] <=  8'h64;        memory[18615] <=  8'h69;        memory[18616] <=  8'h66;        memory[18617] <=  8'h68;        memory[18618] <=  8'h65;        memory[18619] <=  8'h71;        memory[18620] <=  8'h6a;        memory[18621] <=  8'h77;        memory[18622] <=  8'h62;        memory[18623] <=  8'h65;        memory[18624] <=  8'h6e;        memory[18625] <=  8'h20;        memory[18626] <=  8'h6d;        memory[18627] <=  8'h64;        memory[18628] <=  8'h73;        memory[18629] <=  8'h6c;        memory[18630] <=  8'h76;        memory[18631] <=  8'h6b;        memory[18632] <=  8'h63;        memory[18633] <=  8'h78;        memory[18634] <=  8'h20;        memory[18635] <=  8'h6f;        memory[18636] <=  8'h78;        memory[18637] <=  8'h69;        memory[18638] <=  8'h63;        memory[18639] <=  8'h6a;        memory[18640] <=  8'h76;        memory[18641] <=  8'h64;        memory[18642] <=  8'h66;        memory[18643] <=  8'h65;        memory[18644] <=  8'h71;        memory[18645] <=  8'h6e;        memory[18646] <=  8'h20;        memory[18647] <=  8'h64;        memory[18648] <=  8'h6d;        memory[18649] <=  8'h73;        memory[18650] <=  8'h6c;        memory[18651] <=  8'h63;        memory[18652] <=  8'h78;        memory[18653] <=  8'h6b;        memory[18654] <=  8'h20;        memory[18655] <=  8'h6f;        memory[18656] <=  8'h78;        memory[18657] <=  8'h63;        memory[18658] <=  8'h76;        memory[18659] <=  8'h6a;        memory[18660] <=  8'h64;        memory[18661] <=  8'h62;        memory[18662] <=  8'h71;        memory[18663] <=  8'h77;        memory[18664] <=  8'h65;        memory[18665] <=  8'h6e;        memory[18666] <=  8'h6d;        memory[18667] <=  8'h64;        memory[18668] <=  8'h6c;        memory[18669] <=  8'h73;        memory[18670] <=  8'h2c;        memory[18671] <=  8'h76;        memory[18672] <=  8'h63;        memory[18673] <=  8'h78;        memory[18674] <=  8'h20;        memory[18675] <=  8'h63;        memory[18676] <=  8'h6f;        memory[18677] <=  8'h69;        memory[18678] <=  8'h76;        memory[18679] <=  8'h68;        memory[18680] <=  8'h73;        memory[18681] <=  8'h64;        memory[18682] <=  8'h62;        memory[18683] <=  8'h71;        memory[18684] <=  8'h77;        memory[18685] <=  8'h65;        memory[18686] <=  8'h6e;        memory[18687] <=  8'h64;        memory[18688] <=  8'h6b;        memory[18689] <=  8'h73;        memory[18690] <=  8'h76;        memory[18691] <=  8'h6f;        memory[18692] <=  8'h63;        memory[18693] <=  8'h20;        memory[18694] <=  8'h76;        memory[18695] <=  8'h69;        memory[18696] <=  8'h75;        memory[18697] <=  8'h69;        memory[18698] <=  8'h68;        memory[18699] <=  8'h63;        memory[18700] <=  8'h78;        memory[18701] <=  8'h69;        memory[18702] <=  8'h6f;        memory[18703] <=  8'h76;        memory[18704] <=  8'h73;        memory[18705] <=  8'h64;        memory[18706] <=  8'h61;        memory[18707] <=  8'h64;        memory[18708] <=  8'h6e;        memory[18709] <=  8'h77;        memory[18710] <=  8'h71;        memory[18711] <=  8'h6b;        memory[18712] <=  8'h6c;        memory[18713] <=  8'h73;        memory[18714] <=  8'h76;        memory[18715] <=  8'h6e;        memory[18716] <=  8'h62;        memory[18717] <=  8'h20;        memory[18718] <=  8'h64;        memory[18719] <=  8'h66;        memory[18720] <=  8'h6a;        memory[18721] <=  8'h6b;        memory[18722] <=  8'h71;        memory[18723] <=  8'h64;        memory[18724] <=  8'h77;        memory[18725] <=  8'h65;        memory[18726] <=  8'h6e;        memory[18727] <=  8'h62;        memory[18728] <=  8'h20;        memory[18729] <=  8'h64;        memory[18730] <=  8'h73;        memory[18731] <=  8'h76;        memory[18732] <=  8'h68;        memory[18733] <=  8'h64;        memory[18734] <=  8'h61;        memory[18735] <=  8'h71;        memory[18736] <=  8'h77;        memory[18737] <=  8'h6a;        memory[18738] <=  8'h65;        memory[18739] <=  8'h6e;        memory[18740] <=  8'h64;        memory[18741] <=  8'h20;        memory[18742] <=  8'h61;        memory[18743] <=  8'h63;        memory[18744] <=  8'h62;        memory[18745] <=  8'h68;        memory[18746] <=  8'h64;        memory[18747] <=  8'h61;        memory[18748] <=  8'h77;        memory[18749] <=  8'h71;        memory[18750] <=  8'h6e;        memory[18751] <=  8'h20;        memory[18752] <=  8'h62;        memory[18753] <=  8'h73;        memory[18754] <=  8'h76;        memory[18755] <=  8'h61;        memory[18756] <=  8'h67;        memory[18757] <=  8'h76;        memory[18758] <=  8'h68;        memory[18759] <=  8'h67;        memory[18760] <=  8'h61;        memory[18761] <=  8'h73;        memory[18762] <=  8'h6a;        memory[18763] <=  8'h6b;        memory[18764] <=  8'h63;        memory[18765] <=  8'h78;        memory[18766] <=  8'h76;        memory[18767] <=  8'h6e;        memory[18768] <=  8'h73;        memory[18769] <=  8'h64;        memory[18770] <=  8'h20;        memory[18771] <=  8'h66;        memory[18772] <=  8'h62;        memory[18773] <=  8'h64;        memory[18774] <=  8'h61;        memory[18775] <=  8'h73;        memory[18776] <=  8'h76;        memory[18777] <=  8'h67;        memory[18778] <=  8'h63;        memory[18779] <=  8'h79;        memory[18780] <=  8'h7a;        memory[18781] <=  8'h78;        memory[18782] <=  8'h79;        memory[18783] <=  8'h75;        memory[18784] <=  8'h20;        memory[18785] <=  8'h69;        memory[18786] <=  8'h6a;        memory[18787] <=  8'h64;        memory[18788] <=  8'h66;        memory[18789] <=  8'h6b;        memory[18790] <=  8'h61;        memory[18791] <=  8'h64;        memory[18792] <=  8'h63;        memory[18793] <=  8'h78;        memory[18794] <=  8'h68;        memory[18795] <=  8'h20;        memory[18796] <=  8'h67;        memory[18797] <=  8'h61;        memory[18798] <=  8'h68;        memory[18799] <=  8'h75;        memory[18800] <=  8'h64;        memory[18801] <=  8'h73;        memory[18802] <=  8'h69;        memory[18803] <=  8'h6a;        memory[18804] <=  8'h61;        memory[18805] <=  8'h6b;        memory[18806] <=  8'h63;        memory[18807] <=  8'h62;        memory[18808] <=  8'h61;        memory[18809] <=  8'h72;        memory[18810] <=  8'h73;        memory[18811] <=  8'h68;        memory[18812] <=  8'h64;        memory[18813] <=  8'h66;        memory[18814] <=  8'h67;        memory[18815] <=  8'h73;        memory[18816] <=  8'h68;        memory[18817] <=  8'h64;        memory[18818] <=  8'h66;        memory[18819] <=  8'h68;        memory[18820] <=  8'h64;        memory[18821] <=  8'h6a;        memory[18822] <=  8'h68;        memory[18823] <=  8'h62;        memory[18824] <=  8'h67;        memory[18825] <=  8'h63;        memory[18826] <=  8'h61;        memory[18827] <=  8'h66;        memory[18828] <=  8'h73;        memory[18829] <=  8'h79;        memory[18830] <=  8'h67;        memory[18831] <=  8'h6b;        memory[18832] <=  8'h75;        memory[18833] <=  8'h64;        memory[18834] <=  8'h68;        memory[18835] <=  8'h62;        memory[18836] <=  8'h77;        memory[18837] <=  8'h76;        memory[18838] <=  8'h67;        memory[18839] <=  8'h61;        memory[18840] <=  8'h66;        memory[18841] <=  8'h64;        memory[18842] <=  8'h74;        memory[18843] <=  8'h75;        memory[18844] <=  8'h66;        memory[18845] <=  8'h79;        memory[18846] <=  8'h67;        memory[18847] <=  8'h69;        memory[18848] <=  8'h75;        memory[18849] <=  8'h68;        memory[18850] <=  8'h6c;        memory[18851] <=  8'h6a;        memory[18852] <=  8'h62;        memory[18853] <=  8'h6b;        memory[18854] <=  8'h68;        memory[18855] <=  8'h76;        memory[18856] <=  8'h67;        memory[18857] <=  8'h63;        memory[18858] <=  8'h66;        memory[18859] <=  8'h78;        memory[18860] <=  8'h64;        memory[18861] <=  8'h74;        memory[18862] <=  8'h75;        memory[18863] <=  8'h79;        memory[18864] <=  8'h69;        memory[18865] <=  8'h75;        memory[18866] <=  8'h68;        memory[18867] <=  8'h6c;        memory[18868] <=  8'h6a;        memory[18869] <=  8'h6b;        memory[18870] <=  8'h67;        memory[18871] <=  8'h6a;        memory[18872] <=  8'h63;        memory[18873] <=  8'h66;        memory[18874] <=  8'h68;        memory[18875] <=  8'h64;        memory[18876] <=  8'h67;        memory[18877] <=  8'h72;        memory[18878] <=  8'h79;        memory[18879] <=  8'h74;        memory[18880] <=  8'h66;        memory[18881] <=  8'h75;        memory[18882] <=  8'h79;        memory[18883] <=  8'h69;        memory[18884] <=  8'h68;        memory[18885] <=  8'h6c;        memory[18886] <=  8'h62;        memory[18887] <=  8'h6d;        memory[18888] <=  8'h76;        memory[18889] <=  8'h6e;        memory[18890] <=  8'h63;        memory[18891] <=  8'h66;        memory[18892] <=  8'h68;        memory[18893] <=  8'h64;        memory[18894] <=  8'h74;        memory[18895] <=  8'h75;        memory[18896] <=  8'h67;        memory[18897] <=  8'h79;        memory[18898] <=  8'h69;        memory[18899] <=  8'h68;        memory[18900] <=  8'h75;        memory[18901] <=  8'h6a;        memory[18902] <=  8'h6c;        memory[18903] <=  8'h62;        memory[18904] <=  8'h6d;        memory[18905] <=  8'h76;        memory[18906] <=  8'h6e;        memory[18907] <=  8'h63;        memory[18908] <=  8'h66;        memory[18909] <=  8'h68;        memory[18910] <=  8'h67;        memory[18911] <=  8'h79;        memory[18912] <=  8'h68;        memory[18913] <=  8'h75;        memory[18914] <=  8'h6a;        memory[18915] <=  8'h6e;        memory[18916] <=  8'h2c;        memory[18917] <=  8'h62;        memory[18918] <=  8'h6e;        memory[18919] <=  8'h6d;        memory[18920] <=  8'h76;        memory[18921] <=  8'h6e;        memory[18922] <=  8'h63;        memory[18923] <=  8'h66;        memory[18924] <=  8'h68;        memory[18925] <=  8'h74;        memory[18926] <=  8'h79;        memory[18927] <=  8'h69;        memory[18928] <=  8'h75;        memory[18929] <=  8'h6c;        memory[18930] <=  8'h6a;        memory[18931] <=  8'h62;        memory[18932] <=  8'h6d;        memory[18933] <=  8'h76;        memory[18934] <=  8'h6e;        memory[18935] <=  8'h63;        memory[18936] <=  8'h66;        memory[18937] <=  8'h74;        memory[18938] <=  8'h75;        memory[18939] <=  8'h79;        memory[18940] <=  8'h69;        memory[18941] <=  8'h68;        memory[18942] <=  8'h6b;        memory[18943] <=  8'h62;        memory[18944] <=  8'h76;        memory[18945] <=  8'h63;        memory[18946] <=  8'h66;        memory[18947] <=  8'h67;        memory[18948] <=  8'h74;        memory[18949] <=  8'h75;        memory[18950] <=  8'h79;        memory[18951] <=  8'h69;        memory[18952] <=  8'h75;        memory[18953] <=  8'h68;        memory[18954] <=  8'h6a;        memory[18955] <=  8'h6b;        memory[18956] <=  8'h62;        memory[18957] <=  8'h76;        memory[18958] <=  8'h63;        memory[18959] <=  8'h66;        memory[18960] <=  8'h74;        memory[18961] <=  8'h75;        memory[18962] <=  8'h79;        memory[18963] <=  8'h69;        memory[18964] <=  8'h75;        memory[18965] <=  8'h6a;        memory[18966] <=  8'h6b;        memory[18967] <=  8'h6e;        memory[18968] <=  8'h62;        memory[18969] <=  8'h76;        memory[18970] <=  8'h67;        memory[18971] <=  8'h66;        memory[18972] <=  8'h74;        memory[18973] <=  8'h79;        memory[18974] <=  8'h75;        memory[18975] <=  8'h75;        memory[18976] <=  8'h69;        memory[18977] <=  8'h6a;        memory[18978] <=  8'h6b;        memory[18979] <=  8'h68;        memory[18980] <=  8'h62;        memory[18981] <=  8'h6a;        memory[18982] <=  8'h67;        memory[18983] <=  8'h68;        memory[18984] <=  8'h66;        memory[18985] <=  8'h79;        memory[18986] <=  8'h74;        memory[18987] <=  8'h79;        memory[18988] <=  8'h69;        memory[18989] <=  8'h75;        memory[18990] <=  8'h64;        memory[18991] <=  8'h6a;        memory[18992] <=  8'h6b;        memory[18993] <=  8'h68;        memory[18994] <=  8'h63;        memory[18995] <=  8'h7a;        memory[18996] <=  8'h67;        memory[18997] <=  8'h68;        memory[18998] <=  8'h74;        memory[18999] <=  8'h75;        memory[19000] <=  8'h79;        memory[19001] <=  8'h69;        memory[19002] <=  8'h61;        memory[19003] <=  8'h73;        memory[19004] <=  8'h75;        memory[19005] <=  8'h6a;        memory[19006] <=  8'h6b;        memory[19007] <=  8'h62;        memory[19008] <=  8'h6e;        memory[19009] <=  8'h61;        memory[19010] <=  8'h76;        memory[19011] <=  8'h63;        memory[19012] <=  8'h66;        memory[19013] <=  8'h68;        memory[19014] <=  8'h75;        memory[19015] <=  8'h61;        memory[19016] <=  8'h73;        memory[19017] <=  8'h79;        memory[19018] <=  8'h64;        memory[19019] <=  8'h75;        memory[19020] <=  8'h69;        memory[19021] <=  8'h6a;        memory[19022] <=  8'h61;        memory[19023] <=  8'h6b;        memory[19024] <=  8'h62;        memory[19025] <=  8'h63;        memory[19026] <=  8'h78;        memory[19027] <=  8'h68;        memory[19028] <=  8'h67;        memory[19029] <=  8'h79;        memory[19030] <=  8'h75;        memory[19031] <=  8'h7a;        memory[19032] <=  8'h63;        memory[19033] <=  8'h61;        memory[19034] <=  8'h73;        memory[19035] <=  8'h69;        memory[19036] <=  8'h75;        memory[19037] <=  8'h6f;        memory[19038] <=  8'h69;        memory[19039] <=  8'h6a;        memory[19040] <=  8'h61;        memory[19041] <=  8'h6c;        memory[19042] <=  8'h63;        memory[19043] <=  8'h78;        memory[19044] <=  8'h62;        memory[19045] <=  8'h63;        memory[19046] <=  8'h20;        memory[19047] <=  8'h6e;        memory[19048] <=  8'h76;        memory[19049] <=  8'h63;        memory[19050] <=  8'h61;        memory[19051] <=  8'h64;        memory[19052] <=  8'h73;        memory[19053] <=  8'h67;        memory[19054] <=  8'h79;        memory[19055] <=  8'h68;        memory[19056] <=  8'h75;        memory[19057] <=  8'h61;        memory[19058] <=  8'h6a;        memory[19059] <=  8'h6b;        memory[19060] <=  8'h78;        memory[19061] <=  8'h62;        memory[19062] <=  8'h20;        memory[19063] <=  8'h6e;        memory[19064] <=  8'h76;        memory[19065] <=  8'h63;        memory[19066] <=  8'h61;        memory[19067] <=  8'h73;        memory[19068] <=  8'h67;        memory[19069] <=  8'h68;        memory[19070] <=  8'h75;        memory[19071] <=  8'h6a;        memory[19072] <=  8'h6c;        memory[19073] <=  8'h6b;        memory[19074] <=  8'h63;        memory[19075] <=  8'h78;        memory[19076] <=  8'h20;        memory[19077] <=  8'h6a;        memory[19078] <=  8'h6b;        memory[19079] <=  8'h68;        memory[19080] <=  8'h61;        memory[19081] <=  8'h73;        memory[19082] <=  8'h76;        memory[19083] <=  8'h64;        memory[19084] <=  8'h6e;        memory[19085] <=  8'h20;        memory[19086] <=  8'h62;        memory[19087] <=  8'h6e;        memory[19088] <=  8'h6d;        memory[19089] <=  8'h6b;        memory[19090] <=  8'h77;        memory[19091] <=  8'h64;        memory[19092] <=  8'h6f;        memory[19093] <=  8'h77;        memory[19094] <=  8'h69;        memory[19095] <=  8'h6f;        memory[19096] <=  8'h75;        memory[19097] <=  8'h69;        memory[19098] <=  8'h68;        memory[19099] <=  8'h62;        memory[19100] <=  8'h6e;        memory[19101] <=  8'h6b;        memory[19102] <=  8'h77;        memory[19103] <=  8'h69;        memory[19104] <=  8'h6f;        memory[19105] <=  8'h75;        memory[19106] <=  8'h71;        memory[19107] <=  8'h69;        memory[19108] <=  8'h79;        memory[19109] <=  8'h67;        memory[19110] <=  8'h6a;        memory[19111] <=  8'h64;        memory[19112] <=  8'h61;        memory[19113] <=  8'h76;        memory[19114] <=  8'h62;        memory[19115] <=  8'h6e;        memory[19116] <=  8'h6b;        memory[19117] <=  8'h6f;        memory[19118] <=  8'h70;        memory[19119] <=  8'h64;        memory[19120] <=  8'h76;        memory[19121] <=  8'h69;        memory[19122] <=  8'h6f;        memory[19123] <=  8'h75;        memory[19124] <=  8'h69;        memory[19125] <=  8'h48;        memory[19126] <=  8'h42;        memory[19127] <=  8'h6b;        memory[19128] <=  8'h64;        memory[19129] <=  8'h6e;        memory[19130] <=  8'h6c;        memory[19131] <=  8'h71;        memory[19132] <=  8'h6b;        memory[19133] <=  8'h6d;        memory[19134] <=  8'h6a;        memory[19135] <=  8'h70;        memory[19136] <=  8'h69;        memory[19137] <=  8'h6f;        memory[19138] <=  8'h68;        memory[19139] <=  8'h65;        memory[19140] <=  8'h66;        memory[19141] <=  8'h75;        memory[19142] <=  8'h67;        memory[19143] <=  8'h69;        memory[19144] <=  8'h73;        memory[19145] <=  8'h61;        memory[19146] <=  8'h62;        memory[19147] <=  8'h64;        memory[19148] <=  8'h6b;        memory[19149] <=  8'h6a;        memory[19150] <=  8'h6b;        memory[19151] <=  8'h6c;        memory[19152] <=  8'h6a;        memory[19153] <=  8'h69;        memory[19154] <=  8'h73;        memory[19155] <=  8'h6f;        memory[19156] <=  8'h71;        memory[19157] <=  8'h68;        memory[19158] <=  8'h77;        memory[19159] <=  8'h67;        memory[19160] <=  8'h69;        memory[19161] <=  8'h79;        memory[19162] <=  8'h6a;        memory[19163] <=  8'h64;        memory[19164] <=  8'h76;        memory[19165] <=  8'h62;        memory[19166] <=  8'h6e;        memory[19167] <=  8'h61;        memory[19168] <=  8'h73;        memory[19169] <=  8'h66;        memory[19170] <=  8'h6c;        memory[19171] <=  8'h6b;        memory[19172] <=  8'h64;        memory[19173] <=  8'h6a;        memory[19174] <=  8'h68;        memory[19175] <=  8'h63;        memory[19176] <=  8'h67;        memory[19177] <=  8'h6a;        memory[19178] <=  8'h76;        memory[19179] <=  8'h73;        memory[19180] <=  8'h64;        memory[19181] <=  8'h62;        memory[19182] <=  8'h62;        memory[19183] <=  8'h61;        memory[19184] <=  8'h72;        memory[19185] <=  8'h62;        memory[19186] <=  8'h62;        memory[19187] <=  8'h73;        memory[19188] <=  8'h62;        memory[19189] <=  8'h67;        memory[19190] <=  8'h73;        memory[19191] <=  8'h66;        memory[19192] <=  8'h67;        memory[19193] <=  8'h61;        memory[19194] <=  8'h68;        memory[19195] <=  8'h66;        memory[19196] <=  8'h73;        memory[19197] <=  8'h68;        memory[19198] <=  8'h61;        memory[19199] <=  8'h66;        memory[19200] <=  8'h73;        memory[19201] <=  8'h66;        memory[19202] <=  8'h68;        memory[19203] <=  8'h61;        memory[19204] <=  8'h69;        memory[19205] <=  8'h64;        memory[19206] <=  8'h75;        memory[19207] <=  8'h67;        memory[19208] <=  8'h64;        memory[19209] <=  8'h77;        memory[19210] <=  8'h62;        memory[19211] <=  8'h61;        memory[19212] <=  8'h62;        memory[19213] <=  8'h72;        memory[19214] <=  8'h62;        memory[19215] <=  8'h61;        memory[19216] <=  8'h62;        memory[19217] <=  8'h62;        memory[19218] <=  8'h74;        memory[19219] <=  8'h62;        memory[19220] <=  8'h62;        memory[19221] <=  8'h62;        memory[19222] <=  8'h62;        memory[19223] <=  8'h62;        memory[19224] <=  8'h62;        memory[19225] <=  8'h62;        memory[19226] <=  8'h62;        memory[19227] <=  8'h61;        memory[19228] <=  8'h62;        memory[19229] <=  8'h62;        memory[19230] <=  8'h72;        memory[19231] <=  8'h74;        memory[19232] <=  8'h62;        memory[19233] <=  8'h62;        memory[19234] <=  8'h61;        memory[19235] <=  8'h62;        memory[19236] <=  8'h72;        memory[19237] <=  8'h62;        memory[19238] <=  8'h74;        memory[19239] <=  8'h62;        memory[19240] <=  8'h62;        memory[19241] <=  8'h62;        memory[19242] <=  8'h63;        memory[19243] <=  8'h61;        memory[19244] <=  8'h72;        memory[19245] <=  8'h74;        memory[19246] <=  8'h73;        memory[19247] <=  8'h62;        memory[19248] <=  8'h61;        memory[19249] <=  8'h72;        memory[19250] <=  8'h74;        memory[19251] <=  8'h74;        memory[19252] <=  8'h62;        memory[19253] <=  8'h61;        memory[19254] <=  8'h72;        memory[19255] <=  8'h74;        memory[19256] <=  8'h78;        memory[19257] <=  8'h61;        memory[19258] <=  8'h74;        memory[19259] <=  8'h6b;        memory[19260] <=  8'h73;        memory[19261] <=  8'h68;        memory[19262] <=  8'h63;        memory[19263] <=  8'h66;        memory[19264] <=  8'h69;        memory[19265] <=  8'h77;        memory[19266] <=  8'h68;        memory[19267] <=  8'h61;        memory[19268] <=  8'h74;        memory[19269] <=  8'h61;        memory[19270] <=  8'h6e;        memory[19271] <=  8'h61;        memory[19272] <=  8'h62;        memory[19273] <=  8'h61;        memory[19274] <=  8'h63;        memory[19275] <=  8'h61;        memory[19276] <=  8'h74;        memory[19277] <=  8'h61;        memory[19278] <=  8'h62;        memory[19279] <=  8'h61;        memory[19280] <=  8'h72;        memory[19281] <=  8'h63;        memory[19282] <=  8'h61;        memory[19283] <=  8'h68;        memory[19284] <=  8'h64;        memory[19285] <=  8'h75;        memory[19286] <=  8'h63;        memory[19287] <=  8'h74;        memory[19288] <=  8'h61;        memory[19289] <=  8'h64;        memory[19290] <=  8'h61;        memory[19291] <=  8'h61;        memory[19292] <=  8'h63;        memory[19293] <=  8'h61;        memory[19294] <=  8'h72;        memory[19295] <=  8'h63;        memory[19296] <=  8'h74;        memory[19297] <=  8'h72;        memory[19298] <=  8'h63;        memory[19299] <=  8'h61;        memory[19300] <=  8'h74;        memory[19301] <=  8'h72;        memory[19302] <=  8'h63;        memory[19303] <=  8'h61;        memory[19304] <=  8'h74;        memory[19305] <=  8'h63;        memory[19306] <=  8'h62;        memory[19307] <=  8'h61;        memory[19308] <=  8'h74;        memory[19309] <=  8'h62;        memory[19310] <=  8'h72;        memory[19311] <=  8'h63;        memory[19312] <=  8'h61;        memory[19313] <=  8'h74;        memory[19314] <=  8'h72;        memory[19315] <=  8'h6e;        memory[19316] <=  8'h62;        memory[19317] <=  8'h61;        memory[19318] <=  8'h63;        memory[19319] <=  8'h61;        memory[19320] <=  8'h74;        memory[19321] <=  8'h79;        memory[19322] <=  8'h73;        memory[19323] <=  8'h6e;        memory[19324] <=  8'h63;        memory[19325] <=  8'h74;        memory[19326] <=  8'h61;        memory[19327] <=  8'h6e;        memory[19328] <=  8'h62;        memory[19329] <=  8'h61;        memory[19330] <=  8'h63;        memory[19331] <=  8'h72;        memory[19332] <=  8'h6e;        memory[19333] <=  8'h74;        memory[19334] <=  8'h61;        memory[19335] <=  8'h62;        memory[19336] <=  8'h74;        memory[19337] <=  8'h6e;        memory[19338] <=  8'h61;        memory[19339] <=  8'h72;        memory[19340] <=  8'h62;        memory[19341] <=  8'h78;        memory[19342] <=  8'h74;        memory[19343] <=  8'h61;        memory[19344] <=  8'h72;        memory[19345] <=  8'h62;        memory[19346] <=  8'h61;        memory[19347] <=  8'h72;        memory[19348] <=  8'h74;        memory[19349] <=  8'h74;        memory[19350] <=  8'h62;        memory[19351] <=  8'h61;        memory[19352] <=  8'h72;        memory[19353] <=  8'h74;        memory[19354] <=  8'h78;        memory[19355] <=  8'h61;        memory[19356] <=  8'h74;        memory[19357] <=  8'h6b;        memory[19358] <=  8'h73;        memory[19359] <=  8'h68;        memory[19360] <=  8'h63;        memory[19361] <=  8'h66;        memory[19362] <=  8'h69;        memory[19363] <=  8'h77;        memory[19364] <=  8'h68;        memory[19365] <=  8'h61;        memory[19366] <=  8'h74;        memory[19367] <=  8'h61;        memory[19368] <=  8'h6e;        memory[19369] <=  8'h61;        memory[19370] <=  8'h62;        memory[19371] <=  8'h61;        memory[19372] <=  8'h63;        memory[19373] <=  8'h61;        memory[19374] <=  8'h74;        memory[19375] <=  8'h61;        memory[19376] <=  8'h62;        memory[19377] <=  8'h61;        memory[19378] <=  8'h72;        memory[19379] <=  8'h63;        memory[19380] <=  8'h61;        memory[19381] <=  8'h68;        memory[19382] <=  8'h64;        memory[19383] <=  8'h75;        memory[19384] <=  8'h63;        memory[19385] <=  8'h74;        memory[19386] <=  8'h61;        memory[19387] <=  8'h64;        memory[19388] <=  8'h61;        memory[19389] <=  8'h61;        memory[19390] <=  8'h63;        memory[19391] <=  8'h61;        memory[19392] <=  8'h72;        memory[19393] <=  8'h63;        memory[19394] <=  8'h74;        memory[19395] <=  8'h72;        memory[19396] <=  8'h63;        memory[19397] <=  8'h61;        memory[19398] <=  8'h74;        memory[19399] <=  8'h72;        memory[19400] <=  8'h63;        memory[19401] <=  8'h61;        memory[19402] <=  8'h74;        memory[19403] <=  8'h63;        memory[19404] <=  8'h62;        memory[19405] <=  8'h61;        memory[19406] <=  8'h74;        memory[19407] <=  8'h62;        memory[19408] <=  8'h72;        memory[19409] <=  8'h63;        memory[19410] <=  8'h61;        memory[19411] <=  8'h74;        memory[19412] <=  8'h72;        memory[19413] <=  8'h6e;        memory[19414] <=  8'h62;        memory[19415] <=  8'h61;        memory[19416] <=  8'h63;        memory[19417] <=  8'h61;        memory[19418] <=  8'h74;        memory[19419] <=  8'h79;        memory[19420] <=  8'h73;        memory[19421] <=  8'h6e;        memory[19422] <=  8'h63;        memory[19423] <=  8'h74;        memory[19424] <=  8'h61;        memory[19425] <=  8'h6e;        memory[19426] <=  8'h62;        memory[19427] <=  8'h61;        memory[19428] <=  8'h63;        memory[19429] <=  8'h72;        memory[19430] <=  8'h6e;        memory[19431] <=  8'h74;        memory[19432] <=  8'h61;        memory[19433] <=  8'h62;        memory[19434] <=  8'h74;        memory[19435] <=  8'h6e;        memory[19436] <=  8'h61;        memory[19437] <=  8'h72;        memory[19438] <=  8'h62;        memory[19439] <=  8'h78;        memory[19440] <=  8'h74;        memory[19441] <=  8'h61;        memory[19442] <=  8'h72;        memory[19443] <=  8'h62;        memory[19444] <=  8'h61;        memory[19445] <=  8'h72;        memory[19446] <=  8'h74;        memory[19447] <=  8'h74;        memory[19448] <=  8'h62;        memory[19449] <=  8'h61;        memory[19450] <=  8'h72;        memory[19451] <=  8'h74;        memory[19452] <=  8'h78;        memory[19453] <=  8'h61;        memory[19454] <=  8'h74;        memory[19455] <=  8'h6b;        memory[19456] <=  8'h73;        memory[19457] <=  8'h68;        memory[19458] <=  8'h63;        memory[19459] <=  8'h66;        memory[19460] <=  8'h69;        memory[19461] <=  8'h77;        memory[19462] <=  8'h68;        memory[19463] <=  8'h61;        memory[19464] <=  8'h74;        memory[19465] <=  8'h61;        memory[19466] <=  8'h6e;        memory[19467] <=  8'h61;        memory[19468] <=  8'h62;        memory[19469] <=  8'h61;        memory[19470] <=  8'h63;        memory[19471] <=  8'h61;        memory[19472] <=  8'h74;        memory[19473] <=  8'h61;        memory[19474] <=  8'h62;        memory[19475] <=  8'h61;        memory[19476] <=  8'h72;        memory[19477] <=  8'h63;        memory[19478] <=  8'h61;        memory[19479] <=  8'h68;        memory[19480] <=  8'h64;        memory[19481] <=  8'h75;        memory[19482] <=  8'h63;        memory[19483] <=  8'h74;        memory[19484] <=  8'h61;        memory[19485] <=  8'h64;        memory[19486] <=  8'h61;        memory[19487] <=  8'h61;        memory[19488] <=  8'h63;        memory[19489] <=  8'h61;        memory[19490] <=  8'h72;        memory[19491] <=  8'h63;        memory[19492] <=  8'h74;        memory[19493] <=  8'h72;        memory[19494] <=  8'h63;        memory[19495] <=  8'h61;        memory[19496] <=  8'h74;        memory[19497] <=  8'h72;        memory[19498] <=  8'h63;        memory[19499] <=  8'h61;        memory[19500] <=  8'h74;        memory[19501] <=  8'h63;        memory[19502] <=  8'h62;        memory[19503] <=  8'h61;        memory[19504] <=  8'h74;        memory[19505] <=  8'h62;        memory[19506] <=  8'h72;        memory[19507] <=  8'h63;        memory[19508] <=  8'h61;        memory[19509] <=  8'h74;        memory[19510] <=  8'h72;        memory[19511] <=  8'h6e;        memory[19512] <=  8'h62;        memory[19513] <=  8'h61;        memory[19514] <=  8'h63;        memory[19515] <=  8'h61;        memory[19516] <=  8'h74;        memory[19517] <=  8'h79;        memory[19518] <=  8'h73;        memory[19519] <=  8'h6e;        memory[19520] <=  8'h63;        memory[19521] <=  8'h74;        memory[19522] <=  8'h61;        memory[19523] <=  8'h6e;        memory[19524] <=  8'h62;        memory[19525] <=  8'h61;        memory[19526] <=  8'h63;        memory[19527] <=  8'h72;        memory[19528] <=  8'h6e;        memory[19529] <=  8'h74;        memory[19530] <=  8'h61;        memory[19531] <=  8'h62;        memory[19532] <=  8'h74;        memory[19533] <=  8'h6e;        memory[19534] <=  8'h61;        memory[19535] <=  8'h72;        memory[19536] <=  8'h62;        memory[19537] <=  8'h78;        memory[19538] <=  8'h74;        memory[19539] <=  8'h61;        memory[19540] <=  8'h72;        memory[19541] <=  8'h5d;        memory[19542] <=  8'h5d;        memory[19543] <=  8'h65;        memory[19544] <=  8'h66;        memory[19545] <=  8'h77;        memory[19546] <=  8'h65;        memory[19547] <=  8'h5d;        memory[19548] <=  8'h65;        memory[19549] <=  8'h67;        memory[19550] <=  8'h73;        memory[19551] <=  8'h67;        memory[19552] <=  8'h66;        memory[19553] <=  8'h62;        memory[19554] <=  8'h61;        memory[19555] <=  8'h72;        memory[19556] <=  8'h74;        memory[19557] <=  8'h74;        memory[19558] <=  8'h62;        memory[19559] <=  8'h61;        memory[19560] <=  8'h72;        memory[19561] <=  8'h74;        memory[19562] <=  8'h78;        memory[19563] <=  8'h61;        memory[19564] <=  8'h74;        memory[19565] <=  8'h6b;        memory[19566] <=  8'h73;        memory[19567] <=  8'h68;        memory[19568] <=  8'h63;        memory[19569] <=  8'h66;        memory[19570] <=  8'h69;        memory[19571] <=  8'h77;        memory[19572] <=  8'h68;        memory[19573] <=  8'h61;        memory[19574] <=  8'h74;        memory[19575] <=  8'h61;        memory[19576] <=  8'h6e;        memory[19577] <=  8'h61;        memory[19578] <=  8'h62;        memory[19579] <=  8'h61;        memory[19580] <=  8'h63;        memory[19581] <=  8'h61;        memory[19582] <=  8'h74;        memory[19583] <=  8'h61;        memory[19584] <=  8'h62;        memory[19585] <=  8'h61;        memory[19586] <=  8'h72;        memory[19587] <=  8'h63;        memory[19588] <=  8'h61;        memory[19589] <=  8'h68;        memory[19590] <=  8'h64;        memory[19591] <=  8'h75;        memory[19592] <=  8'h63;        memory[19593] <=  8'h74;        memory[19594] <=  8'h61;        memory[19595] <=  8'h64;        memory[19596] <=  8'h61;        memory[19597] <=  8'h61;        memory[19598] <=  8'h63;        memory[19599] <=  8'h61;        memory[19600] <=  8'h72;        memory[19601] <=  8'h63;        memory[19602] <=  8'h74;        memory[19603] <=  8'h72;        memory[19604] <=  8'h63;        memory[19605] <=  8'h61;        memory[19606] <=  8'h74;        memory[19607] <=  8'h72;        memory[19608] <=  8'h63;        memory[19609] <=  8'h61;        memory[19610] <=  8'h74;        memory[19611] <=  8'h63;        memory[19612] <=  8'h62;        memory[19613] <=  8'h61;        memory[19614] <=  8'h74;        memory[19615] <=  8'h62;        memory[19616] <=  8'h72;        memory[19617] <=  8'h63;        memory[19618] <=  8'h61;        memory[19619] <=  8'h74;        memory[19620] <=  8'h72;        memory[19621] <=  8'h6e;        memory[19622] <=  8'h62;        memory[19623] <=  8'h61;        memory[19624] <=  8'h63;        memory[19625] <=  8'h61;        memory[19626] <=  8'h74;        memory[19627] <=  8'h79;        memory[19628] <=  8'h73;        memory[19629] <=  8'h6e;        memory[19630] <=  8'h63;        memory[19631] <=  8'h74;        memory[19632] <=  8'h61;        memory[19633] <=  8'h6e;        memory[19634] <=  8'h62;        memory[19635] <=  8'h61;        memory[19636] <=  8'h63;        memory[19637] <=  8'h72;        memory[19638] <=  8'h6e;        memory[19639] <=  8'h74;        memory[19640] <=  8'h61;        memory[19641] <=  8'h62;        memory[19642] <=  8'h74;        memory[19643] <=  8'h6e;        memory[19644] <=  8'h61;        memory[19645] <=  8'h72;        memory[19646] <=  8'h62;        memory[19647] <=  8'h78;        memory[19648] <=  8'h74;        memory[19649] <=  8'h61;        memory[19650] <=  8'h72;        memory[19651] <=  8'h62;        memory[19652] <=  8'h61;        memory[19653] <=  8'h72;        memory[19654] <=  8'h74;        memory[19655] <=  8'h74;        memory[19656] <=  8'h62;        memory[19657] <=  8'h61;        memory[19658] <=  8'h72;        memory[19659] <=  8'h74;        memory[19660] <=  8'h78;        memory[19661] <=  8'h61;        memory[19662] <=  8'h74;        memory[19663] <=  8'h6b;        memory[19664] <=  8'h73;        memory[19665] <=  8'h68;        memory[19666] <=  8'h63;        memory[19667] <=  8'h66;        memory[19668] <=  8'h69;        memory[19669] <=  8'h77;        memory[19670] <=  8'h68;        memory[19671] <=  8'h61;        memory[19672] <=  8'h74;        memory[19673] <=  8'h61;        memory[19674] <=  8'h6e;        memory[19675] <=  8'h61;        memory[19676] <=  8'h62;        memory[19677] <=  8'h61;        memory[19678] <=  8'h63;        memory[19679] <=  8'h61;        memory[19680] <=  8'h74;        memory[19681] <=  8'h61;        memory[19682] <=  8'h62;        memory[19683] <=  8'h61;        memory[19684] <=  8'h72;        memory[19685] <=  8'h63;        memory[19686] <=  8'h61;        memory[19687] <=  8'h68;        memory[19688] <=  8'h64;        memory[19689] <=  8'h75;        memory[19690] <=  8'h63;        memory[19691] <=  8'h74;        memory[19692] <=  8'h61;        memory[19693] <=  8'h64;        memory[19694] <=  8'h61;        memory[19695] <=  8'h61;        memory[19696] <=  8'h63;        memory[19697] <=  8'h61;        memory[19698] <=  8'h72;        memory[19699] <=  8'h63;        memory[19700] <=  8'h74;        memory[19701] <=  8'h72;        memory[19702] <=  8'h63;        memory[19703] <=  8'h61;        memory[19704] <=  8'h74;        memory[19705] <=  8'h72;        memory[19706] <=  8'h63;        memory[19707] <=  8'h61;        memory[19708] <=  8'h74;        memory[19709] <=  8'h63;        memory[19710] <=  8'h62;        memory[19711] <=  8'h61;        memory[19712] <=  8'h74;        memory[19713] <=  8'h62;        memory[19714] <=  8'h72;        memory[19715] <=  8'h63;        memory[19716] <=  8'h61;        memory[19717] <=  8'h74;        memory[19718] <=  8'h72;        memory[19719] <=  8'h6e;        memory[19720] <=  8'h62;        memory[19721] <=  8'h61;        memory[19722] <=  8'h63;        memory[19723] <=  8'h61;        memory[19724] <=  8'h74;        memory[19725] <=  8'h79;        memory[19726] <=  8'h73;        memory[19727] <=  8'h6e;        memory[19728] <=  8'h63;        memory[19729] <=  8'h74;        memory[19730] <=  8'h61;        memory[19731] <=  8'h6e;        memory[19732] <=  8'h62;        memory[19733] <=  8'h61;        memory[19734] <=  8'h63;        memory[19735] <=  8'h72;        memory[19736] <=  8'h6e;        memory[19737] <=  8'h74;        memory[19738] <=  8'h61;        memory[19739] <=  8'h62;        memory[19740] <=  8'h74;        memory[19741] <=  8'h6e;        memory[19742] <=  8'h61;        memory[19743] <=  8'h72;        memory[19744] <=  8'h62;        memory[19745] <=  8'h78;        memory[19746] <=  8'h74;        memory[19747] <=  8'h61;        memory[19748] <=  8'h72;        memory[19749] <=  8'h64;        memory[19750] <=  8'h66;        memory[19751] <=  8'h73;        memory[19752] <=  8'h67;        memory[19753] <=  8'h76;        memory[19754] <=  8'h68;        memory[19755] <=  8'h62;        memory[19756] <=  8'h6b;        memory[19757] <=  8'h6a;        memory[19758] <=  8'h6e;        memory[19759] <=  8'h6d;        memory[19760] <=  8'h62;        memory[19761] <=  8'h76;        memory[19762] <=  8'h78;        memory[19763] <=  8'h63;        memory[19764] <=  8'h73;        memory[19765] <=  8'h66;        memory[19766] <=  8'h72;        memory[19767] <=  8'h74;        memory[19768] <=  8'h79;        memory[19769] <=  8'h75;        memory[19770] <=  8'h6a;        memory[19771] <=  8'h6e;        memory[19772] <=  8'h62;        memory[19773] <=  8'h76;        memory[19774] <=  8'h63;        memory[19775] <=  8'h64;        memory[19776] <=  8'h74;        memory[19777] <=  8'h79;        memory[19778] <=  8'h75;        memory[19779] <=  8'h69;        memory[19780] <=  8'h6b;        memory[19781] <=  8'h6d;        memory[19782] <=  8'h6e;        memory[19783] <=  8'h62;        memory[19784] <=  8'h76;        memory[19785] <=  8'h63;        memory[19786] <=  8'h78;        memory[19787] <=  8'h73;        memory[19788] <=  8'h64;        memory[19789] <=  8'h72;        memory[19790] <=  8'h74;        memory[19791] <=  8'h79;        memory[19792] <=  8'h75;        memory[19793] <=  8'h69;        memory[19794] <=  8'h6b;        memory[19795] <=  8'h6d;        memory[19796] <=  8'h6e;        memory[19797] <=  8'h62;        memory[19798] <=  8'h76;        memory[19799] <=  8'h63;        memory[19800] <=  8'h73;        memory[19801] <=  8'h77;        memory[19802] <=  8'h33;        memory[19803] <=  8'h34;        memory[19804] <=  8'h35;        memory[19805] <=  8'h36;        memory[19806] <=  8'h37;        memory[19807] <=  8'h38;        memory[19808] <=  8'h69;        memory[19809] <=  8'h6b;        memory[19810] <=  8'h6d;        memory[19811] <=  8'h6e;        memory[19812] <=  8'h62;        memory[19813] <=  8'h76;        memory[19814] <=  8'h63;        memory[19815] <=  8'h64;        memory[19816] <=  8'h65;        memory[19817] <=  8'h72;        memory[19818] <=  8'h36;        memory[19819] <=  8'h37;        memory[19820] <=  8'h38;        memory[19821] <=  8'h69;        memory[19822] <=  8'h6f;        memory[19823] <=  8'h6b;        memory[19824] <=  8'h6a;        memory[19825] <=  8'h6e;        memory[19826] <=  8'h62;        memory[19827] <=  8'h76;        memory[19828] <=  8'h63;        memory[19829] <=  8'h64;        memory[19830] <=  8'h72;        memory[19831] <=  8'h74;        memory[19832] <=  8'h79;        memory[19833] <=  8'h75;        memory[19834] <=  8'h73;        memory[19835] <=  8'h6a;        memory[19836] <=  8'h63;        memory[19837] <=  8'h6e;        memory[19838] <=  8'h62;        memory[19839] <=  8'h64;        memory[19840] <=  8'h66;        memory[19841] <=  8'h73;        memory[19842] <=  8'h74;        memory[19843] <=  8'h79;        memory[19844] <=  8'h75;        memory[19845] <=  8'h61;        memory[19846] <=  8'h69;        memory[19847] <=  8'h6b;        memory[19848] <=  8'h78;        memory[19849] <=  8'h6d;        memory[19850] <=  8'h6e;        memory[19851] <=  8'h73;        memory[19852] <=  8'h6a;        memory[19853] <=  8'h6f;        memory[19854] <=  8'h64;        memory[19855] <=  8'h6c;        memory[19856] <=  8'h63;        memory[19857] <=  8'h78;        memory[19858] <=  8'h62;        memory[19859] <=  8'h61;        memory[19860] <=  8'h72;        memory[19861] <=  8'h74;        memory[19862] <=  8'h78;        memory[19863] <=  8'h61;        memory[19864] <=  8'h74;        memory[19865] <=  8'h6b;        memory[19866] <=  8'h73;        memory[19867] <=  8'h68;        memory[19868] <=  8'h63;        memory[19869] <=  8'h66;        memory[19870] <=  8'h69;        memory[19871] <=  8'h77;        memory[19872] <=  8'h68;        memory[19873] <=  8'h61;        memory[19874] <=  8'h74;        memory[19875] <=  8'h61;        memory[19876] <=  8'h6e;        memory[19877] <=  8'h61;        memory[19878] <=  8'h62;        memory[19879] <=  8'h61;        memory[19880] <=  8'h63;        memory[19881] <=  8'h61;        memory[19882] <=  8'h74;        memory[19883] <=  8'h61;        memory[19884] <=  8'h62;        memory[19885] <=  8'h61;        memory[19886] <=  8'h72;        memory[19887] <=  8'h63;        memory[19888] <=  8'h61;        memory[19889] <=  8'h68;        memory[19890] <=  8'h64;        memory[19891] <=  8'h75;        memory[19892] <=  8'h63;        memory[19893] <=  8'h74;        memory[19894] <=  8'h61;        memory[19895] <=  8'h64;        memory[19896] <=  8'h61;        memory[19897] <=  8'h61;        memory[19898] <=  8'h63;        memory[19899] <=  8'h61;        memory[19900] <=  8'h72;        memory[19901] <=  8'h62;        memory[19902] <=  8'h61;        memory[19903] <=  8'h72;        memory[19904] <=  8'h74;        memory[19905] <=  8'h78;        memory[19906] <=  8'h61;        memory[19907] <=  8'h74;        memory[19908] <=  8'h6b;        memory[19909] <=  8'h73;        memory[19910] <=  8'h68;        memory[19911] <=  8'h63;        memory[19912] <=  8'h66;        memory[19913] <=  8'h69;        memory[19914] <=  8'h77;        memory[19915] <=  8'h68;        memory[19916] <=  8'h61;        memory[19917] <=  8'h74;        memory[19918] <=  8'h61;        memory[19919] <=  8'h6e;        memory[19920] <=  8'h61;        memory[19921] <=  8'h62;        memory[19922] <=  8'h61;        memory[19923] <=  8'h63;        memory[19924] <=  8'h61;        memory[19925] <=  8'h74;        memory[19926] <=  8'h61;        memory[19927] <=  8'h62;        memory[19928] <=  8'h61;        memory[19929] <=  8'h72;        memory[19930] <=  8'h63;        memory[19931] <=  8'h61;        memory[19932] <=  8'h68;        memory[19933] <=  8'h64;        memory[19934] <=  8'h75;        memory[19935] <=  8'h63;        memory[19936] <=  8'h74;        memory[19937] <=  8'h61;        memory[19938] <=  8'h64;        memory[19939] <=  8'h61;        memory[19940] <=  8'h61;        memory[19941] <=  8'h63;        memory[19942] <=  8'h61;        memory[19943] <=  8'h72;        memory[19944] <=  8'h62;        memory[19945] <=  8'h61;        memory[19946] <=  8'h72;        memory[19947] <=  8'h74;        memory[19948] <=  8'h78;        memory[19949] <=  8'h61;        memory[19950] <=  8'h74;        memory[19951] <=  8'h6b;        memory[19952] <=  8'h73;        memory[19953] <=  8'h68;        memory[19954] <=  8'h63;        memory[19955] <=  8'h66;        memory[19956] <=  8'h69;        memory[19957] <=  8'h77;        memory[19958] <=  8'h68;        memory[19959] <=  8'h61;        memory[19960] <=  8'h74;        memory[19961] <=  8'h61;        memory[19962] <=  8'h6e;        memory[19963] <=  8'h61;        memory[19964] <=  8'h62;        memory[19965] <=  8'h61;        memory[19966] <=  8'h63;        memory[19967] <=  8'h61;        memory[19968] <=  8'h74;        memory[19969] <=  8'h61;        memory[19970] <=  8'h62;        memory[19971] <=  8'h61;        memory[19972] <=  8'h72;        memory[19973] <=  8'h63;        memory[19974] <=  8'h61;        memory[19975] <=  8'h68;        memory[19976] <=  8'h64;        memory[19977] <=  8'h75;        memory[19978] <=  8'h63;        memory[19979] <=  8'h74;        memory[19980] <=  8'h61;        memory[19981] <=  8'h64;        memory[19982] <=  8'h61;        memory[19983] <=  8'h61;        memory[19984] <=  8'h63;        memory[19985] <=  8'h61;        memory[19986] <=  8'h72;        memory[19987] <=  8'h62;        memory[19988] <=  8'h61;        memory[19989] <=  8'h72;        memory[19990] <=  8'h74;        memory[19991] <=  8'h78;        memory[19992] <=  8'h61;        memory[19993] <=  8'h74;        memory[19994] <=  8'h6b;        memory[19995] <=  8'h73;        memory[19996] <=  8'h68;        memory[19997] <=  8'h63;        memory[19998] <=  8'h66;        memory[19999] <=  8'h69;        memory[20000] <=  8'h77;        memory[20001] <=  8'h68;        memory[20002] <=  8'h61;        memory[20003] <=  8'h74;        memory[20004] <=  8'h61;        memory[20005] <=  8'h6e;        memory[20006] <=  8'h61;        memory[20007] <=  8'h62;        memory[20008] <=  8'h61;        memory[20009] <=  8'h63;        memory[20010] <=  8'h61;        memory[20011] <=  8'h74;        memory[20012] <=  8'h61;        memory[20013] <=  8'h62;        memory[20014] <=  8'h61;        memory[20015] <=  8'h72;        memory[20016] <=  8'h63;        memory[20017] <=  8'h61;        memory[20018] <=  8'h68;        memory[20019] <=  8'h64;        memory[20020] <=  8'h75;        memory[20021] <=  8'h63;        memory[20022] <=  8'h74;        memory[20023] <=  8'h61;        memory[20024] <=  8'h64;        memory[20025] <=  8'h61;        memory[20026] <=  8'h61;        memory[20027] <=  8'h63;        memory[20028] <=  8'h61;        memory[20029] <=  8'h72;        memory[20030] <=  8'h62;        memory[20031] <=  8'h61;        memory[20032] <=  8'h72;        memory[20033] <=  8'h74;        memory[20034] <=  8'h78;        memory[20035] <=  8'h61;        memory[20036] <=  8'h74;        memory[20037] <=  8'h6b;        memory[20038] <=  8'h73;        memory[20039] <=  8'h68;        memory[20040] <=  8'h63;        memory[20041] <=  8'h66;        memory[20042] <=  8'h69;        memory[20043] <=  8'h77;        memory[20044] <=  8'h68;        memory[20045] <=  8'h61;        memory[20046] <=  8'h74;        memory[20047] <=  8'h61;        memory[20048] <=  8'h6e;        memory[20049] <=  8'h61;        memory[20050] <=  8'h62;        memory[20051] <=  8'h61;        memory[20052] <=  8'h63;        memory[20053] <=  8'h61;        memory[20054] <=  8'h74;        memory[20055] <=  8'h61;        memory[20056] <=  8'h62;        memory[20057] <=  8'h61;        memory[20058] <=  8'h72;        memory[20059] <=  8'h63;        memory[20060] <=  8'h61;        memory[20061] <=  8'h68;        memory[20062] <=  8'h64;        memory[20063] <=  8'h75;        memory[20064] <=  8'h63;        memory[20065] <=  8'h74;        memory[20066] <=  8'h61;        memory[20067] <=  8'h64;        memory[20068] <=  8'h61;        memory[20069] <=  8'h61;        memory[20070] <=  8'h63;        memory[20071] <=  8'h61;        memory[20072] <=  8'h72;        memory[20073] <=  8'h62;        memory[20074] <=  8'h61;        memory[20075] <=  8'h72;        memory[20076] <=  8'h74;        memory[20077] <=  8'h78;        memory[20078] <=  8'h61;        memory[20079] <=  8'h74;        memory[20080] <=  8'h6b;        memory[20081] <=  8'h73;        memory[20082] <=  8'h68;        memory[20083] <=  8'h63;        memory[20084] <=  8'h66;        memory[20085] <=  8'h69;        memory[20086] <=  8'h77;        memory[20087] <=  8'h68;        memory[20088] <=  8'h61;        memory[20089] <=  8'h74;        memory[20090] <=  8'h61;        memory[20091] <=  8'h6e;        memory[20092] <=  8'h61;        memory[20093] <=  8'h62;        memory[20094] <=  8'h61;        memory[20095] <=  8'h63;        memory[20096] <=  8'h61;        memory[20097] <=  8'h74;        memory[20098] <=  8'h61;        memory[20099] <=  8'h62;        memory[20100] <=  8'h61;        memory[20101] <=  8'h72;        memory[20102] <=  8'h63;        memory[20103] <=  8'h61;        memory[20104] <=  8'h68;        memory[20105] <=  8'h64;        memory[20106] <=  8'h75;        memory[20107] <=  8'h63;        memory[20108] <=  8'h74;        memory[20109] <=  8'h61;        memory[20110] <=  8'h64;        memory[20111] <=  8'h61;        memory[20112] <=  8'h61;        memory[20113] <=  8'h63;        memory[20114] <=  8'h61;        memory[20115] <=  8'h72;        memory[20116] <=  8'h62;        memory[20117] <=  8'h61;        memory[20118] <=  8'h72;        memory[20119] <=  8'h74;        memory[20120] <=  8'h78;        memory[20121] <=  8'h61;        memory[20122] <=  8'h74;        memory[20123] <=  8'h6b;        memory[20124] <=  8'h73;        memory[20125] <=  8'h68;        memory[20126] <=  8'h63;        memory[20127] <=  8'h66;        memory[20128] <=  8'h69;        memory[20129] <=  8'h77;        memory[20130] <=  8'h68;        memory[20131] <=  8'h61;        memory[20132] <=  8'h74;        memory[20133] <=  8'h61;        memory[20134] <=  8'h6e;        memory[20135] <=  8'h61;        memory[20136] <=  8'h62;        memory[20137] <=  8'h61;        memory[20138] <=  8'h63;        memory[20139] <=  8'h61;        memory[20140] <=  8'h74;        memory[20141] <=  8'h61;        memory[20142] <=  8'h62;        memory[20143] <=  8'h61;        memory[20144] <=  8'h72;        memory[20145] <=  8'h63;        memory[20146] <=  8'h61;        memory[20147] <=  8'h68;        memory[20148] <=  8'h64;        memory[20149] <=  8'h75;        memory[20150] <=  8'h63;        memory[20151] <=  8'h74;        memory[20152] <=  8'h61;        memory[20153] <=  8'h64;        memory[20154] <=  8'h61;        memory[20155] <=  8'h61;        memory[20156] <=  8'h63;        memory[20157] <=  8'h61;        memory[20158] <=  8'h72;        memory[20159] <=  8'h62;        memory[20160] <=  8'h61;        memory[20161] <=  8'h72;        memory[20162] <=  8'h74;        memory[20163] <=  8'h78;        memory[20164] <=  8'h61;        memory[20165] <=  8'h74;        memory[20166] <=  8'h6b;        memory[20167] <=  8'h73;        memory[20168] <=  8'h68;        memory[20169] <=  8'h63;        memory[20170] <=  8'h66;        memory[20171] <=  8'h69;        memory[20172] <=  8'h77;        memory[20173] <=  8'h68;        memory[20174] <=  8'h61;        memory[20175] <=  8'h74;        memory[20176] <=  8'h61;        memory[20177] <=  8'h6e;        memory[20178] <=  8'h61;        memory[20179] <=  8'h62;        memory[20180] <=  8'h61;        memory[20181] <=  8'h63;        memory[20182] <=  8'h61;        memory[20183] <=  8'h74;        memory[20184] <=  8'h61;        memory[20185] <=  8'h62;        memory[20186] <=  8'h61;        memory[20187] <=  8'h72;        memory[20188] <=  8'h63;        memory[20189] <=  8'h61;        memory[20190] <=  8'h68;        memory[20191] <=  8'h64;        memory[20192] <=  8'h75;        memory[20193] <=  8'h63;        memory[20194] <=  8'h74;        memory[20195] <=  8'h61;        memory[20196] <=  8'h64;        memory[20197] <=  8'h61;        memory[20198] <=  8'h61;        memory[20199] <=  8'h63;        memory[20200] <=  8'h61;        memory[20201] <=  8'h72;        memory[20202] <=  8'h62;        memory[20203] <=  8'h61;        memory[20204] <=  8'h72;        memory[20205] <=  8'h74;        memory[20206] <=  8'h78;        memory[20207] <=  8'h61;        memory[20208] <=  8'h74;        memory[20209] <=  8'h6b;        memory[20210] <=  8'h73;        memory[20211] <=  8'h68;        memory[20212] <=  8'h63;        memory[20213] <=  8'h66;        memory[20214] <=  8'h69;        memory[20215] <=  8'h77;        memory[20216] <=  8'h68;        memory[20217] <=  8'h61;        memory[20218] <=  8'h74;        memory[20219] <=  8'h61;        memory[20220] <=  8'h6e;        memory[20221] <=  8'h61;        memory[20222] <=  8'h62;        memory[20223] <=  8'h61;        memory[20224] <=  8'h63;        memory[20225] <=  8'h61;        memory[20226] <=  8'h74;        memory[20227] <=  8'h61;        memory[20228] <=  8'h62;        memory[20229] <=  8'h61;        memory[20230] <=  8'h72;        memory[20231] <=  8'h63;        memory[20232] <=  8'h61;        memory[20233] <=  8'h68;        memory[20234] <=  8'h64;        memory[20235] <=  8'h75;        memory[20236] <=  8'h63;        memory[20237] <=  8'h74;        memory[20238] <=  8'h61;        memory[20239] <=  8'h64;        memory[20240] <=  8'h61;        memory[20241] <=  8'h61;        memory[20242] <=  8'h63;        memory[20243] <=  8'h61;        memory[20244] <=  8'h72;        memory[20245] <=  8'h62;        memory[20246] <=  8'h61;        memory[20247] <=  8'h72;        memory[20248] <=  8'h74;        memory[20249] <=  8'h74;        memory[20250] <=  8'h62;        memory[20251] <=  8'h61;        memory[20252] <=  8'h72;        memory[20253] <=  8'h74;        memory[20254] <=  8'h78;        memory[20255] <=  8'h61;        memory[20256] <=  8'h74;        memory[20257] <=  8'h6b;        memory[20258] <=  8'h73;        memory[20259] <=  8'h68;        memory[20260] <=  8'h63;        memory[20261] <=  8'h66;        memory[20262] <=  8'h69;        memory[20263] <=  8'h77;        memory[20264] <=  8'h68;        memory[20265] <=  8'h61;        memory[20266] <=  8'h74;        memory[20267] <=  8'h61;        memory[20268] <=  8'h6e;        memory[20269] <=  8'h61;        memory[20270] <=  8'h62;        memory[20271] <=  8'h61;        memory[20272] <=  8'h63;        memory[20273] <=  8'h61;        memory[20274] <=  8'h74;        memory[20275] <=  8'h61;        memory[20276] <=  8'h62;        memory[20277] <=  8'h61;        memory[20278] <=  8'h72;        memory[20279] <=  8'h63;        memory[20280] <=  8'h61;        memory[20281] <=  8'h68;        memory[20282] <=  8'h64;        memory[20283] <=  8'h75;        memory[20284] <=  8'h63;        memory[20285] <=  8'h74;        memory[20286] <=  8'h61;        memory[20287] <=  8'h64;        memory[20288] <=  8'h61;        memory[20289] <=  8'h61;        memory[20290] <=  8'h63;        memory[20291] <=  8'h61;        memory[20292] <=  8'h72;        memory[20293] <=  8'h63;        memory[20294] <=  8'h74;        memory[20295] <=  8'h72;        memory[20296] <=  8'h63;        memory[20297] <=  8'h61;        memory[20298] <=  8'h74;        memory[20299] <=  8'h72;        memory[20300] <=  8'h63;        memory[20301] <=  8'h61;        memory[20302] <=  8'h74;        memory[20303] <=  8'h63;        memory[20304] <=  8'h62;        memory[20305] <=  8'h61;        memory[20306] <=  8'h74;        memory[20307] <=  8'h62;        memory[20308] <=  8'h72;        memory[20309] <=  8'h63;        memory[20310] <=  8'h61;        memory[20311] <=  8'h72;        memory[20312] <=  8'h62;        memory[20313] <=  8'h78;        memory[20314] <=  8'h74;        memory[20315] <=  8'h61;        memory[20316] <=  8'h72;        memory[20317] <=  8'h64;        memory[20318] <=  8'h66;        memory[20319] <=  8'h73;        memory[20320] <=  8'h67;        memory[20321] <=  8'h76;        memory[20322] <=  8'h68;        memory[20323] <=  8'h62;        memory[20324] <=  8'h6b;        memory[20325] <=  8'h6a;        memory[20326] <=  8'h6e;        memory[20327] <=  8'h6d;        memory[20328] <=  8'h62;        memory[20329] <=  8'h76;        memory[20330] <=  8'h78;        memory[20331] <=  8'h63;        memory[20332] <=  8'h73;        memory[20333] <=  8'h66;        memory[20334] <=  8'h72;        memory[20335] <=  8'h74;        memory[20336] <=  8'h79;        memory[20337] <=  8'h75;        memory[20338] <=  8'h6a;        memory[20339] <=  8'h6e;        memory[20340] <=  8'h62;        memory[20341] <=  8'h76;        memory[20342] <=  8'h63;        memory[20343] <=  8'h64;        memory[20344] <=  8'h74;        memory[20345] <=  8'h79;        memory[20346] <=  8'h75;        memory[20347] <=  8'h69;        memory[20348] <=  8'h6b;        memory[20349] <=  8'h6d;        memory[20350] <=  8'h6e;        memory[20351] <=  8'h62;        memory[20352] <=  8'h76;        memory[20353] <=  8'h63;        memory[20354] <=  8'h78;        memory[20355] <=  8'h73;        memory[20356] <=  8'h64;        memory[20357] <=  8'h72;        memory[20358] <=  8'h74;        memory[20359] <=  8'h79;        memory[20360] <=  8'h75;        memory[20361] <=  8'h69;        memory[20362] <=  8'h6b;        memory[20363] <=  8'h6d;        memory[20364] <=  8'h6e;        memory[20365] <=  8'h62;        memory[20366] <=  8'h76;        memory[20367] <=  8'h63;        memory[20368] <=  8'h73;        memory[20369] <=  8'h77;        memory[20370] <=  8'h33;        memory[20371] <=  8'h34;        memory[20372] <=  8'h35;        memory[20373] <=  8'h36;        memory[20374] <=  8'h37;        memory[20375] <=  8'h38;        memory[20376] <=  8'h69;        memory[20377] <=  8'h6b;        memory[20378] <=  8'h6d;        memory[20379] <=  8'h6e;        memory[20380] <=  8'h62;        memory[20381] <=  8'h76;        memory[20382] <=  8'h63;        memory[20383] <=  8'h64;        memory[20384] <=  8'h65;        memory[20385] <=  8'h72;        memory[20386] <=  8'h36;        memory[20387] <=  8'h37;        memory[20388] <=  8'h38;        memory[20389] <=  8'h69;        memory[20390] <=  8'h6f;        memory[20391] <=  8'h6b;        memory[20392] <=  8'h6a;        memory[20393] <=  8'h6e;        memory[20394] <=  8'h62;        memory[20395] <=  8'h76;        memory[20396] <=  8'h63;        memory[20397] <=  8'h64;        memory[20398] <=  8'h72;        memory[20399] <=  8'h74;        memory[20400] <=  8'h79;        memory[20401] <=  8'h75;        memory[20402] <=  8'h73;        memory[20403] <=  8'h6a;        memory[20404] <=  8'h63;        memory[20405] <=  8'h6e;        memory[20406] <=  8'h62;        memory[20407] <=  8'h64;        memory[20408] <=  8'h66;        memory[20409] <=  8'h73;        memory[20410] <=  8'h74;        memory[20411] <=  8'h79;        memory[20412] <=  8'h75;        memory[20413] <=  8'h61;        memory[20414] <=  8'h69;        memory[20415] <=  8'h6b;        memory[20416] <=  8'h78;        memory[20417] <=  8'h6d;        memory[20418] <=  8'h6e;        memory[20419] <=  8'h73;        memory[20420] <=  8'h6a;        memory[20421] <=  8'h6f;        memory[20422] <=  8'h64;        memory[20423] <=  8'h6c;        memory[20424] <=  8'h63;        memory[20425] <=  8'h78;        memory[20426] <=  8'h2c;        memory[20427] <=  8'h6d;        memory[20428] <=  8'h73;        memory[20429] <=  8'h6b;        memory[20430] <=  8'h64;        memory[20431] <=  8'h6c;        memory[20432] <=  8'h70;        memory[20433] <=  8'h5b;        memory[20434] <=  8'h3b;        memory[20435] <=  8'h73;        memory[20436] <=  8'h6c;        memory[20437] <=  8'h64;        memory[20438] <=  8'h70;        memory[20439] <=  8'h76;        memory[20440] <=  8'h63;        memory[20441] <=  8'h5b;        memory[20442] <=  8'h78;        memory[20443] <=  8'h76;        memory[20444] <=  8'h63;        memory[20445] <=  8'h5b;        memory[20446] <=  8'h78;        memory[20447] <=  8'h70;        memory[20448] <=  8'h6f;        memory[20449] <=  8'h20;        memory[20450] <=  8'h62;        memory[20451] <=  8'h61;        memory[20452] <=  8'h72;        memory[20453] <=  8'h74;        memory[20454] <=  8'h74;        memory[20455] <=  8'h62;        memory[20456] <=  8'h61;        memory[20457] <=  8'h72;        memory[20458] <=  8'h74;        memory[20459] <=  8'h78;        memory[20460] <=  8'h61;        memory[20461] <=  8'h74;        memory[20462] <=  8'h6b;        memory[20463] <=  8'h73;        memory[20464] <=  8'h68;        memory[20465] <=  8'h63;        memory[20466] <=  8'h66;        memory[20467] <=  8'h69;        memory[20468] <=  8'h77;        memory[20469] <=  8'h68;        memory[20470] <=  8'h61;        memory[20471] <=  8'h69;        memory[20472] <=  8'h6a;        memory[20473] <=  8'h78;        memory[20474] <=  8'h5d;        memory[20475] <=  8'h65;        memory[20476] <=  8'h6b;        memory[20477] <=  8'h6f;        memory[20478] <=  8'h39;        memory[20479] <=  8'h64;        memory[20480] <=  8'h75;        memory[20481] <=  8'h38;        memory[20482] <=  8'h79;        memory[20483] <=  8'h20;        memory[20484] <=  8'h37;        memory[20485] <=  8'h63;        memory[20486] <=  8'h67;        memory[20487] <=  8'h78;        memory[20488] <=  8'h63;        memory[20489] <=  8'h75;        memory[20490] <=  8'h68;        memory[20491] <=  8'h69;        memory[20492] <=  8'h6a;        memory[20493] <=  8'h77;        memory[20494] <=  8'h69;        memory[20495] <=  8'h64;        memory[20496] <=  8'h66;        memory[20497] <=  8'h68;        memory[20498] <=  8'h75;        memory[20499] <=  8'h76;        memory[20500] <=  8'h64;        memory[20501] <=  8'h62;        memory[20502] <=  8'h66;        memory[20503] <=  8'h6a;        memory[20504] <=  8'h6e;        memory[20505] <=  8'h6b;        memory[20506] <=  8'h6a;        memory[20507] <=  8'h65;        memory[20508] <=  8'h38;        memory[20509] <=  8'h66;        memory[20510] <=  8'h37;        memory[20511] <=  8'h67;        memory[20512] <=  8'h79;        memory[20513] <=  8'h76;        memory[20514] <=  8'h63;        memory[20515] <=  8'h68;        memory[20516] <=  8'h69;        memory[20517] <=  8'h6a;        memory[20518] <=  8'h33;        memory[20519] <=  8'h65;        memory[20520] <=  8'h67;        memory[20521] <=  8'h79;        memory[20522] <=  8'h72;        memory[20523] <=  8'h64;        memory[20524] <=  8'h62;        memory[20525] <=  8'h6e;        memory[20526] <=  8'h63;        memory[20527] <=  8'h7a;        memory[20528] <=  8'h6a;        memory[20529] <=  8'h6f;        memory[20530] <=  8'h66;        memory[20531] <=  8'h78;        memory[20532] <=  8'h6a;        memory[20533] <=  8'h69;        memory[20534] <=  8'h63;        memory[20535] <=  8'h68;        memory[20536] <=  8'h62;        memory[20537] <=  8'h6e;        memory[20538] <=  8'h6d;        memory[20539] <=  8'h63;        memory[20540] <=  8'h73;        memory[20541] <=  8'h6c;        memory[20542] <=  8'h6b;        memory[20543] <=  8'h6a;        memory[20544] <=  8'h69;        memory[20545] <=  8'h68;        memory[20546] <=  8'h76;        memory[20547] <=  8'h75;        memory[20548] <=  8'h69;        memory[20549] <=  8'h64;        memory[20550] <=  8'h68;        memory[20551] <=  8'h75;        memory[20552] <=  8'h67;        memory[20553] <=  8'h79;        memory[20554] <=  8'h62;        memory[20555] <=  8'h68;        memory[20556] <=  8'h65;        memory[20557] <=  8'h6a;        memory[20558] <=  8'h72;        memory[20559] <=  8'h6b;        memory[20560] <=  8'h6a;        memory[20561] <=  8'h6f;        memory[20562] <=  8'h64;        memory[20563] <=  8'h67;        memory[20564] <=  8'h69;        memory[20565] <=  8'h75;        memory[20566] <=  8'h69;        memory[20567] <=  8'h67;        memory[20568] <=  8'h76;        memory[20569] <=  8'h79;        memory[20570] <=  8'h75;        memory[20571] <=  8'h67;        memory[20572] <=  8'h78;        memory[20573] <=  8'h68;        memory[20574] <=  8'h63;        memory[20575] <=  8'h20;        memory[20576] <=  8'h20;        memory[20577] <=  8'h20;        memory[20578] <=  8'h78;        memory[20579] <=  8'h76;        memory[20580] <=  8'h20;        memory[20581] <=  8'h63;        memory[20582] <=  8'h78;        memory[20583] <=  8'h67;        memory[20584] <=  8'h79;        memory[20585] <=  8'h63;        memory[20586] <=  8'h75;        memory[20587] <=  8'h68;        memory[20588] <=  8'h6a;        memory[20589] <=  8'h6b;        memory[20590] <=  8'h61;        memory[20591] <=  8'h6c;        memory[20592] <=  8'h78;        memory[20593] <=  8'h76;        memory[20594] <=  8'h70;        memory[20595] <=  8'h6f;        memory[20596] <=  8'h69;        memory[20597] <=  8'h6a;        memory[20598] <=  8'h69;        memory[20599] <=  8'h68;        memory[20600] <=  8'h6a;        memory[20601] <=  8'h62;        memory[20602] <=  8'h77;        memory[20603] <=  8'h65;        memory[20604] <=  8'h6e;        memory[20605] <=  8'h61;        memory[20606] <=  8'h66;        memory[20607] <=  8'h6d;        memory[20608] <=  8'h64;        memory[20609] <=  8'h6b;        memory[20610] <=  8'h6d;        memory[20611] <=  8'h76;        memory[20612] <=  8'h6c;        memory[20613] <=  8'h63;        memory[20614] <=  8'h6f;        memory[20615] <=  8'h64;        memory[20616] <=  8'h69;        memory[20617] <=  8'h75;        memory[20618] <=  8'h68;        memory[20619] <=  8'h73;        memory[20620] <=  8'h66;        memory[20621] <=  8'h65;        memory[20622] <=  8'h62;        memory[20623] <=  8'h6e;        memory[20624] <=  8'h64;        memory[20625] <=  8'h73;        memory[20626] <=  8'h63;        memory[20627] <=  8'h6b;        memory[20628] <=  8'h20;        memory[20629] <=  8'h78;        memory[20630] <=  8'h6a;        memory[20631] <=  8'h78;        memory[20632] <=  8'h63;        memory[20633] <=  8'h73;        memory[20634] <=  8'h64;        memory[20635] <=  8'h66;        memory[20636] <=  8'h6b;        memory[20637] <=  8'h64;        memory[20638] <=  8'h6e;        memory[20639] <=  8'h6d;        memory[20640] <=  8'h64;        memory[20641] <=  8'h73;        memory[20642] <=  8'h63;        memory[20643] <=  8'h6b;        memory[20644] <=  8'h78;        memory[20645] <=  8'h6c;        memory[20646] <=  8'h6f;        memory[20647] <=  8'h66;        memory[20648] <=  8'h6a;        memory[20649] <=  8'h69;        memory[20650] <=  8'h61;        memory[20651] <=  8'h62;        memory[20652] <=  8'h6e;        memory[20653] <=  8'h20;        memory[20654] <=  8'h78;        memory[20655] <=  8'h6b;        memory[20656] <=  8'h6d;        memory[20657] <=  8'h20;        memory[20658] <=  8'h6f;        memory[20659] <=  8'h63;        memory[20660] <=  8'h76;        memory[20661] <=  8'h73;        memory[20662] <=  8'h64;        memory[20663] <=  8'h69;        memory[20664] <=  8'h66;        memory[20665] <=  8'h68;        memory[20666] <=  8'h65;        memory[20667] <=  8'h71;        memory[20668] <=  8'h6a;        memory[20669] <=  8'h77;        memory[20670] <=  8'h62;        memory[20671] <=  8'h65;        memory[20672] <=  8'h6e;        memory[20673] <=  8'h20;        memory[20674] <=  8'h6d;        memory[20675] <=  8'h64;        memory[20676] <=  8'h73;        memory[20677] <=  8'h6c;        memory[20678] <=  8'h76;        memory[20679] <=  8'h6b;        memory[20680] <=  8'h63;        memory[20681] <=  8'h78;        memory[20682] <=  8'h20;        memory[20683] <=  8'h6f;        memory[20684] <=  8'h78;        memory[20685] <=  8'h69;        memory[20686] <=  8'h63;        memory[20687] <=  8'h6a;        memory[20688] <=  8'h76;        memory[20689] <=  8'h64;        memory[20690] <=  8'h66;        memory[20691] <=  8'h65;        memory[20692] <=  8'h71;        memory[20693] <=  8'h6e;        memory[20694] <=  8'h20;        memory[20695] <=  8'h64;        memory[20696] <=  8'h6d;        memory[20697] <=  8'h73;        memory[20698] <=  8'h6c;        memory[20699] <=  8'h63;        memory[20700] <=  8'h78;        memory[20701] <=  8'h6b;        memory[20702] <=  8'h20;        memory[20703] <=  8'h6f;        memory[20704] <=  8'h78;        memory[20705] <=  8'h63;        memory[20706] <=  8'h76;        memory[20707] <=  8'h6a;        memory[20708] <=  8'h64;        memory[20709] <=  8'h62;        memory[20710] <=  8'h71;        memory[20711] <=  8'h77;        memory[20712] <=  8'h65;        memory[20713] <=  8'h6e;        memory[20714] <=  8'h6d;        memory[20715] <=  8'h64;        memory[20716] <=  8'h6c;        memory[20717] <=  8'h73;        memory[20718] <=  8'h2c;        memory[20719] <=  8'h76;        memory[20720] <=  8'h63;        memory[20721] <=  8'h78;        memory[20722] <=  8'h20;        memory[20723] <=  8'h63;        memory[20724] <=  8'h6f;        memory[20725] <=  8'h69;        memory[20726] <=  8'h76;        memory[20727] <=  8'h68;        memory[20728] <=  8'h73;        memory[20729] <=  8'h64;        memory[20730] <=  8'h62;        memory[20731] <=  8'h71;        memory[20732] <=  8'h77;        memory[20733] <=  8'h65;        memory[20734] <=  8'h6e;        memory[20735] <=  8'h64;        memory[20736] <=  8'h6b;        memory[20737] <=  8'h73;        memory[20738] <=  8'h76;        memory[20739] <=  8'h6f;        memory[20740] <=  8'h63;        memory[20741] <=  8'h20;        memory[20742] <=  8'h76;        memory[20743] <=  8'h69;        memory[20744] <=  8'h75;        memory[20745] <=  8'h69;        memory[20746] <=  8'h68;        memory[20747] <=  8'h63;        memory[20748] <=  8'h78;        memory[20749] <=  8'h69;        memory[20750] <=  8'h6f;        memory[20751] <=  8'h76;        memory[20752] <=  8'h73;        memory[20753] <=  8'h64;        memory[20754] <=  8'h61;        memory[20755] <=  8'h64;        memory[20756] <=  8'h6e;        memory[20757] <=  8'h77;        memory[20758] <=  8'h71;        memory[20759] <=  8'h6b;        memory[20760] <=  8'h6c;        memory[20761] <=  8'h73;        memory[20762] <=  8'h76;        memory[20763] <=  8'h6e;        memory[20764] <=  8'h62;        memory[20765] <=  8'h20;        memory[20766] <=  8'h64;        memory[20767] <=  8'h66;        memory[20768] <=  8'h6a;        memory[20769] <=  8'h6b;        memory[20770] <=  8'h71;        memory[20771] <=  8'h64;        memory[20772] <=  8'h77;        memory[20773] <=  8'h65;        memory[20774] <=  8'h6e;        memory[20775] <=  8'h62;        memory[20776] <=  8'h20;        memory[20777] <=  8'h64;        memory[20778] <=  8'h73;        memory[20779] <=  8'h76;        memory[20780] <=  8'h68;        memory[20781] <=  8'h64;        memory[20782] <=  8'h61;        memory[20783] <=  8'h71;        memory[20784] <=  8'h77;        memory[20785] <=  8'h6a;        memory[20786] <=  8'h65;        memory[20787] <=  8'h6e;        memory[20788] <=  8'h64;        memory[20789] <=  8'h20;        memory[20790] <=  8'h61;        memory[20791] <=  8'h63;        memory[20792] <=  8'h62;        memory[20793] <=  8'h68;        memory[20794] <=  8'h64;        memory[20795] <=  8'h61;        memory[20796] <=  8'h77;        memory[20797] <=  8'h71;        memory[20798] <=  8'h6e;        memory[20799] <=  8'h20;        memory[20800] <=  8'h62;        memory[20801] <=  8'h73;        memory[20802] <=  8'h76;        memory[20803] <=  8'h61;        memory[20804] <=  8'h67;        memory[20805] <=  8'h76;        memory[20806] <=  8'h68;        memory[20807] <=  8'h67;        memory[20808] <=  8'h61;        memory[20809] <=  8'h73;        memory[20810] <=  8'h6a;        memory[20811] <=  8'h6b;        memory[20812] <=  8'h63;        memory[20813] <=  8'h78;        memory[20814] <=  8'h76;        memory[20815] <=  8'h6e;        memory[20816] <=  8'h73;        memory[20817] <=  8'h64;        memory[20818] <=  8'h20;        memory[20819] <=  8'h66;        memory[20820] <=  8'h62;        memory[20821] <=  8'h64;        memory[20822] <=  8'h61;        memory[20823] <=  8'h73;        memory[20824] <=  8'h76;        memory[20825] <=  8'h67;        memory[20826] <=  8'h63;        memory[20827] <=  8'h79;        memory[20828] <=  8'h7a;        memory[20829] <=  8'h78;        memory[20830] <=  8'h79;        memory[20831] <=  8'h75;        memory[20832] <=  8'h20;        memory[20833] <=  8'h69;        memory[20834] <=  8'h6a;        memory[20835] <=  8'h64;        memory[20836] <=  8'h66;        memory[20837] <=  8'h6b;        memory[20838] <=  8'h61;        memory[20839] <=  8'h64;        memory[20840] <=  8'h63;        memory[20841] <=  8'h78;        memory[20842] <=  8'h68;        memory[20843] <=  8'h20;        memory[20844] <=  8'h67;        memory[20845] <=  8'h61;        memory[20846] <=  8'h68;        memory[20847] <=  8'h75;        memory[20848] <=  8'h64;        memory[20849] <=  8'h73;        memory[20850] <=  8'h69;        memory[20851] <=  8'h6a;        memory[20852] <=  8'h61;        memory[20853] <=  8'h6b;        memory[20854] <=  8'h63;        memory[20855] <=  8'h62;        memory[20856] <=  8'h61;        memory[20857] <=  8'h72;        memory[20858] <=  8'h73;        memory[20859] <=  8'h68;        memory[20860] <=  8'h64;        memory[20861] <=  8'h66;        memory[20862] <=  8'h67;        memory[20863] <=  8'h73;        memory[20864] <=  8'h68;        memory[20865] <=  8'h64;        memory[20866] <=  8'h66;        memory[20867] <=  8'h68;        memory[20868] <=  8'h64;        memory[20869] <=  8'h6a;        memory[20870] <=  8'h68;        memory[20871] <=  8'h62;        memory[20872] <=  8'h67;        memory[20873] <=  8'h63;        memory[20874] <=  8'h61;        memory[20875] <=  8'h66;        memory[20876] <=  8'h73;        memory[20877] <=  8'h79;        memory[20878] <=  8'h67;        memory[20879] <=  8'h6b;        memory[20880] <=  8'h75;        memory[20881] <=  8'h64;        memory[20882] <=  8'h68;        memory[20883] <=  8'h62;        memory[20884] <=  8'h77;        memory[20885] <=  8'h76;        memory[20886] <=  8'h67;        memory[20887] <=  8'h61;        memory[20888] <=  8'h66;        memory[20889] <=  8'h64;        memory[20890] <=  8'h74;        memory[20891] <=  8'h75;        memory[20892] <=  8'h66;        memory[20893] <=  8'h79;        memory[20894] <=  8'h67;        memory[20895] <=  8'h69;        memory[20896] <=  8'h75;        memory[20897] <=  8'h68;        memory[20898] <=  8'h6c;        memory[20899] <=  8'h6a;        memory[20900] <=  8'h62;        memory[20901] <=  8'h6b;        memory[20902] <=  8'h68;        memory[20903] <=  8'h76;        memory[20904] <=  8'h67;        memory[20905] <=  8'h63;        memory[20906] <=  8'h66;        memory[20907] <=  8'h78;        memory[20908] <=  8'h64;        memory[20909] <=  8'h74;        memory[20910] <=  8'h75;        memory[20911] <=  8'h79;        memory[20912] <=  8'h69;        memory[20913] <=  8'h75;        memory[20914] <=  8'h68;        memory[20915] <=  8'h6c;        memory[20916] <=  8'h6a;        memory[20917] <=  8'h6b;        memory[20918] <=  8'h67;        memory[20919] <=  8'h6a;        memory[20920] <=  8'h63;        memory[20921] <=  8'h66;        memory[20922] <=  8'h68;        memory[20923] <=  8'h64;        memory[20924] <=  8'h67;        memory[20925] <=  8'h72;        memory[20926] <=  8'h79;        memory[20927] <=  8'h74;        memory[20928] <=  8'h66;        memory[20929] <=  8'h75;        memory[20930] <=  8'h79;        memory[20931] <=  8'h69;        memory[20932] <=  8'h68;        memory[20933] <=  8'h6c;        memory[20934] <=  8'h62;        memory[20935] <=  8'h6d;        memory[20936] <=  8'h76;        memory[20937] <=  8'h6e;        memory[20938] <=  8'h63;        memory[20939] <=  8'h66;        memory[20940] <=  8'h68;        memory[20941] <=  8'h64;        memory[20942] <=  8'h74;        memory[20943] <=  8'h75;        memory[20944] <=  8'h67;        memory[20945] <=  8'h79;        memory[20946] <=  8'h69;        memory[20947] <=  8'h68;        memory[20948] <=  8'h75;        memory[20949] <=  8'h6a;        memory[20950] <=  8'h6c;        memory[20951] <=  8'h62;        memory[20952] <=  8'h6d;        memory[20953] <=  8'h76;        memory[20954] <=  8'h6e;        memory[20955] <=  8'h63;        memory[20956] <=  8'h66;        memory[20957] <=  8'h68;        memory[20958] <=  8'h67;        memory[20959] <=  8'h79;        memory[20960] <=  8'h68;        memory[20961] <=  8'h75;        memory[20962] <=  8'h6a;        memory[20963] <=  8'h6e;        memory[20964] <=  8'h2c;        memory[20965] <=  8'h62;        memory[20966] <=  8'h6e;        memory[20967] <=  8'h6d;        memory[20968] <=  8'h76;        memory[20969] <=  8'h6e;        memory[20970] <=  8'h63;        memory[20971] <=  8'h66;        memory[20972] <=  8'h68;        memory[20973] <=  8'h74;        memory[20974] <=  8'h79;        memory[20975] <=  8'h69;        memory[20976] <=  8'h75;        memory[20977] <=  8'h6c;        memory[20978] <=  8'h6a;        memory[20979] <=  8'h62;        memory[20980] <=  8'h6d;        memory[20981] <=  8'h76;        memory[20982] <=  8'h6e;        memory[20983] <=  8'h63;        memory[20984] <=  8'h66;        memory[20985] <=  8'h74;        memory[20986] <=  8'h75;        memory[20987] <=  8'h79;        memory[20988] <=  8'h69;        memory[20989] <=  8'h68;        memory[20990] <=  8'h6b;        memory[20991] <=  8'h62;        memory[20992] <=  8'h76;        memory[20993] <=  8'h63;        memory[20994] <=  8'h66;        memory[20995] <=  8'h67;        memory[20996] <=  8'h74;        memory[20997] <=  8'h75;        memory[20998] <=  8'h79;        memory[20999] <=  8'h69;        memory[21000] <=  8'h75;        memory[21001] <=  8'h68;        memory[21002] <=  8'h6a;        memory[21003] <=  8'h6b;        memory[21004] <=  8'h62;        memory[21005] <=  8'h76;        memory[21006] <=  8'h63;        memory[21007] <=  8'h66;        memory[21008] <=  8'h74;        memory[21009] <=  8'h75;        memory[21010] <=  8'h79;        memory[21011] <=  8'h69;        memory[21012] <=  8'h75;        memory[21013] <=  8'h6a;        memory[21014] <=  8'h6b;        memory[21015] <=  8'h6e;        memory[21016] <=  8'h62;        memory[21017] <=  8'h76;        memory[21018] <=  8'h67;        memory[21019] <=  8'h66;        memory[21020] <=  8'h74;        memory[21021] <=  8'h79;        memory[21022] <=  8'h75;        memory[21023] <=  8'h75;        memory[21024] <=  8'h69;        memory[21025] <=  8'h6a;        memory[21026] <=  8'h6b;        memory[21027] <=  8'h68;        memory[21028] <=  8'h62;        memory[21029] <=  8'h6a;        memory[21030] <=  8'h67;        memory[21031] <=  8'h68;        memory[21032] <=  8'h66;        memory[21033] <=  8'h79;        memory[21034] <=  8'h74;        memory[21035] <=  8'h79;        memory[21036] <=  8'h69;        memory[21037] <=  8'h75;        memory[21038] <=  8'h64;        memory[21039] <=  8'h6a;        memory[21040] <=  8'h6b;        memory[21041] <=  8'h68;        memory[21042] <=  8'h63;        memory[21043] <=  8'h7a;        memory[21044] <=  8'h67;        memory[21045] <=  8'h68;        memory[21046] <=  8'h74;        memory[21047] <=  8'h75;        memory[21048] <=  8'h79;        memory[21049] <=  8'h69;        memory[21050] <=  8'h61;        memory[21051] <=  8'h73;        memory[21052] <=  8'h75;        memory[21053] <=  8'h6a;        memory[21054] <=  8'h6b;        memory[21055] <=  8'h62;        memory[21056] <=  8'h6e;        memory[21057] <=  8'h61;        memory[21058] <=  8'h76;        memory[21059] <=  8'h63;        memory[21060] <=  8'h66;        memory[21061] <=  8'h68;        memory[21062] <=  8'h75;        memory[21063] <=  8'h61;        memory[21064] <=  8'h73;        memory[21065] <=  8'h79;        memory[21066] <=  8'h64;        memory[21067] <=  8'h75;        memory[21068] <=  8'h69;        memory[21069] <=  8'h6a;        memory[21070] <=  8'h61;        memory[21071] <=  8'h6b;        memory[21072] <=  8'h62;        memory[21073] <=  8'h63;        memory[21074] <=  8'h78;        memory[21075] <=  8'h68;        memory[21076] <=  8'h67;        memory[21077] <=  8'h79;        memory[21078] <=  8'h75;        memory[21079] <=  8'h7a;        memory[21080] <=  8'h63;        memory[21081] <=  8'h61;        memory[21082] <=  8'h73;        memory[21083] <=  8'h69;        memory[21084] <=  8'h75;        memory[21085] <=  8'h6f;        memory[21086] <=  8'h69;        memory[21087] <=  8'h6a;        memory[21088] <=  8'h61;        memory[21089] <=  8'h6c;        memory[21090] <=  8'h63;        memory[21091] <=  8'h78;        memory[21092] <=  8'h62;        memory[21093] <=  8'h63;        memory[21094] <=  8'h20;        memory[21095] <=  8'h6e;        memory[21096] <=  8'h76;        memory[21097] <=  8'h63;        memory[21098] <=  8'h61;        memory[21099] <=  8'h64;        memory[21100] <=  8'h73;        memory[21101] <=  8'h67;        memory[21102] <=  8'h79;        memory[21103] <=  8'h68;        memory[21104] <=  8'h75;        memory[21105] <=  8'h61;        memory[21106] <=  8'h6a;        memory[21107] <=  8'h6b;        memory[21108] <=  8'h78;        memory[21109] <=  8'h62;        memory[21110] <=  8'h20;        memory[21111] <=  8'h6e;        memory[21112] <=  8'h76;        memory[21113] <=  8'h63;        memory[21114] <=  8'h61;        memory[21115] <=  8'h73;        memory[21116] <=  8'h67;        memory[21117] <=  8'h68;        memory[21118] <=  8'h75;        memory[21119] <=  8'h6a;        memory[21120] <=  8'h6c;        memory[21121] <=  8'h6b;        memory[21122] <=  8'h63;        memory[21123] <=  8'h78;        memory[21124] <=  8'h20;        memory[21125] <=  8'h6a;        memory[21126] <=  8'h6b;        memory[21127] <=  8'h68;        memory[21128] <=  8'h61;        memory[21129] <=  8'h73;        memory[21130] <=  8'h76;        memory[21131] <=  8'h64;        memory[21132] <=  8'h6e;        memory[21133] <=  8'h20;        memory[21134] <=  8'h62;        memory[21135] <=  8'h6e;        memory[21136] <=  8'h6d;        memory[21137] <=  8'h6b;        memory[21138] <=  8'h77;        memory[21139] <=  8'h64;        memory[21140] <=  8'h6f;        memory[21141] <=  8'h77;        memory[21142] <=  8'h69;        memory[21143] <=  8'h6f;        memory[21144] <=  8'h75;        memory[21145] <=  8'h69;        memory[21146] <=  8'h68;        memory[21147] <=  8'h62;        memory[21148] <=  8'h6e;        memory[21149] <=  8'h6b;        memory[21150] <=  8'h77;        memory[21151] <=  8'h69;        memory[21152] <=  8'h6f;        memory[21153] <=  8'h75;        memory[21154] <=  8'h71;        memory[21155] <=  8'h69;        memory[21156] <=  8'h79;        memory[21157] <=  8'h67;        memory[21158] <=  8'h6a;        memory[21159] <=  8'h64;        memory[21160] <=  8'h61;        memory[21161] <=  8'h76;        memory[21162] <=  8'h62;        memory[21163] <=  8'h6e;        memory[21164] <=  8'h6b;        memory[21165] <=  8'h6f;        memory[21166] <=  8'h70;        memory[21167] <=  8'h64;        memory[21168] <=  8'h76;        memory[21169] <=  8'h69;        memory[21170] <=  8'h6f;        memory[21171] <=  8'h75;        memory[21172] <=  8'h69;        memory[21173] <=  8'h48;        memory[21174] <=  8'h42;        memory[21175] <=  8'h6b;        memory[21176] <=  8'h64;        memory[21177] <=  8'h6e;        memory[21178] <=  8'h6c;        memory[21179] <=  8'h71;        memory[21180] <=  8'h6b;        memory[21181] <=  8'h6d;        memory[21182] <=  8'h6a;        memory[21183] <=  8'h70;        memory[21184] <=  8'h69;        memory[21185] <=  8'h6f;        memory[21186] <=  8'h68;        memory[21187] <=  8'h65;        memory[21188] <=  8'h66;        memory[21189] <=  8'h75;        memory[21190] <=  8'h67;        memory[21191] <=  8'h69;        memory[21192] <=  8'h73;        memory[21193] <=  8'h61;        memory[21194] <=  8'h62;        memory[21195] <=  8'h64;        memory[21196] <=  8'h6b;        memory[21197] <=  8'h6a;        memory[21198] <=  8'h6b;        memory[21199] <=  8'h6c;        memory[21200] <=  8'h6a;        memory[21201] <=  8'h69;        memory[21202] <=  8'h73;        memory[21203] <=  8'h6f;        memory[21204] <=  8'h71;        memory[21205] <=  8'h68;        memory[21206] <=  8'h77;        memory[21207] <=  8'h67;        memory[21208] <=  8'h69;        memory[21209] <=  8'h79;        memory[21210] <=  8'h6a;        memory[21211] <=  8'h64;        memory[21212] <=  8'h76;        memory[21213] <=  8'h62;        memory[21214] <=  8'h6e;        memory[21215] <=  8'h61;        memory[21216] <=  8'h73;        memory[21217] <=  8'h66;        memory[21218] <=  8'h6c;        memory[21219] <=  8'h6b;        memory[21220] <=  8'h64;        memory[21221] <=  8'h6a;        memory[21222] <=  8'h68;        memory[21223] <=  8'h63;        memory[21224] <=  8'h67;        memory[21225] <=  8'h6a;        memory[21226] <=  8'h76;        memory[21227] <=  8'h73;        memory[21228] <=  8'h64;        memory[21229] <=  8'h62;        memory[21230] <=  8'h62;        memory[21231] <=  8'h61;        memory[21232] <=  8'h72;        memory[21233] <=  8'h62;        memory[21234] <=  8'h62;        memory[21235] <=  8'h73;        memory[21236] <=  8'h62;        memory[21237] <=  8'h67;        memory[21238] <=  8'h73;        memory[21239] <=  8'h66;        memory[21240] <=  8'h67;        memory[21241] <=  8'h61;        memory[21242] <=  8'h68;        memory[21243] <=  8'h66;        memory[21244] <=  8'h73;        memory[21245] <=  8'h68;        memory[21246] <=  8'h61;        memory[21247] <=  8'h66;        memory[21248] <=  8'h73;        memory[21249] <=  8'h66;        memory[21250] <=  8'h68;        memory[21251] <=  8'h61;        memory[21252] <=  8'h69;        memory[21253] <=  8'h64;        memory[21254] <=  8'h75;        memory[21255] <=  8'h67;        memory[21256] <=  8'h64;        memory[21257] <=  8'h77;        memory[21258] <=  8'h62;        memory[21259] <=  8'h61;        memory[21260] <=  8'h62;        memory[21261] <=  8'h72;        memory[21262] <=  8'h62;        memory[21263] <=  8'h61;        memory[21264] <=  8'h62;        memory[21265] <=  8'h62;        memory[21266] <=  8'h74;        memory[21267] <=  8'h62;        memory[21268] <=  8'h62;        memory[21269] <=  8'h62;        memory[21270] <=  8'h62;        memory[21271] <=  8'h62;        memory[21272] <=  8'h62;        memory[21273] <=  8'h62;        memory[21274] <=  8'h62;        memory[21275] <=  8'h61;        memory[21276] <=  8'h62;        memory[21277] <=  8'h62;        memory[21278] <=  8'h72;        memory[21279] <=  8'h74;        memory[21280] <=  8'h62;        memory[21281] <=  8'h62;        memory[21282] <=  8'h61;        memory[21283] <=  8'h62;        memory[21284] <=  8'h72;        memory[21285] <=  8'h62;        memory[21286] <=  8'h74;        memory[21287] <=  8'h62;        memory[21288] <=  8'h62;        memory[21289] <=  8'h62;        memory[21290] <=  8'h63;        memory[21291] <=  8'h61;        memory[21292] <=  8'h72;        memory[21293] <=  8'h74;        memory[21294] <=  8'h73;        memory[21295] <=  8'h62;        memory[21296] <=  8'h61;        memory[21297] <=  8'h72;        memory[21298] <=  8'h74;        memory[21299] <=  8'h74;        memory[21300] <=  8'h62;        memory[21301] <=  8'h61;        memory[21302] <=  8'h72;        memory[21303] <=  8'h74;        memory[21304] <=  8'h78;        memory[21305] <=  8'h61;        memory[21306] <=  8'h74;        memory[21307] <=  8'h6b;        memory[21308] <=  8'h73;        memory[21309] <=  8'h68;        memory[21310] <=  8'h63;        memory[21311] <=  8'h66;        memory[21312] <=  8'h69;        memory[21313] <=  8'h77;        memory[21314] <=  8'h68;        memory[21315] <=  8'h61;        memory[21316] <=  8'h74;        memory[21317] <=  8'h61;        memory[21318] <=  8'h6e;        memory[21319] <=  8'h61;        memory[21320] <=  8'h62;        memory[21321] <=  8'h61;        memory[21322] <=  8'h63;        memory[21323] <=  8'h61;        memory[21324] <=  8'h74;        memory[21325] <=  8'h61;        memory[21326] <=  8'h62;        memory[21327] <=  8'h61;        memory[21328] <=  8'h72;        memory[21329] <=  8'h63;        memory[21330] <=  8'h61;        memory[21331] <=  8'h68;        memory[21332] <=  8'h64;        memory[21333] <=  8'h75;        memory[21334] <=  8'h63;        memory[21335] <=  8'h74;        memory[21336] <=  8'h61;        memory[21337] <=  8'h64;        memory[21338] <=  8'h61;        memory[21339] <=  8'h61;        memory[21340] <=  8'h63;        memory[21341] <=  8'h61;        memory[21342] <=  8'h72;        memory[21343] <=  8'h63;        memory[21344] <=  8'h74;        memory[21345] <=  8'h72;        memory[21346] <=  8'h63;        memory[21347] <=  8'h61;        memory[21348] <=  8'h74;        memory[21349] <=  8'h72;        memory[21350] <=  8'h63;        memory[21351] <=  8'h61;        memory[21352] <=  8'h74;        memory[21353] <=  8'h63;        memory[21354] <=  8'h62;        memory[21355] <=  8'h61;        memory[21356] <=  8'h74;        memory[21357] <=  8'h62;        memory[21358] <=  8'h72;        memory[21359] <=  8'h63;        memory[21360] <=  8'h61;        memory[21361] <=  8'h74;        memory[21362] <=  8'h72;        memory[21363] <=  8'h6e;        memory[21364] <=  8'h62;        memory[21365] <=  8'h61;        memory[21366] <=  8'h63;        memory[21367] <=  8'h61;        memory[21368] <=  8'h74;        memory[21369] <=  8'h79;        memory[21370] <=  8'h73;        memory[21371] <=  8'h6e;        memory[21372] <=  8'h63;        memory[21373] <=  8'h74;        memory[21374] <=  8'h61;        memory[21375] <=  8'h6e;        memory[21376] <=  8'h62;        memory[21377] <=  8'h61;        memory[21378] <=  8'h63;        memory[21379] <=  8'h72;        memory[21380] <=  8'h6e;        memory[21381] <=  8'h74;        memory[21382] <=  8'h61;        memory[21383] <=  8'h62;        memory[21384] <=  8'h74;        memory[21385] <=  8'h6e;        memory[21386] <=  8'h61;        memory[21387] <=  8'h72;        memory[21388] <=  8'h62;        memory[21389] <=  8'h78;        memory[21390] <=  8'h74;        memory[21391] <=  8'h61;        memory[21392] <=  8'h72;        memory[21393] <=  8'h62;        memory[21394] <=  8'h61;        memory[21395] <=  8'h72;        memory[21396] <=  8'h74;        memory[21397] <=  8'h74;        memory[21398] <=  8'h62;        memory[21399] <=  8'h61;        memory[21400] <=  8'h72;        memory[21401] <=  8'h74;        memory[21402] <=  8'h78;        memory[21403] <=  8'h61;        memory[21404] <=  8'h74;        memory[21405] <=  8'h6b;        memory[21406] <=  8'h73;        memory[21407] <=  8'h68;        memory[21408] <=  8'h63;        memory[21409] <=  8'h66;        memory[21410] <=  8'h69;        memory[21411] <=  8'h77;        memory[21412] <=  8'h68;        memory[21413] <=  8'h61;        memory[21414] <=  8'h74;        memory[21415] <=  8'h61;        memory[21416] <=  8'h6e;        memory[21417] <=  8'h61;        memory[21418] <=  8'h62;        memory[21419] <=  8'h61;        memory[21420] <=  8'h63;        memory[21421] <=  8'h61;        memory[21422] <=  8'h74;        memory[21423] <=  8'h61;        memory[21424] <=  8'h62;        memory[21425] <=  8'h61;        memory[21426] <=  8'h72;        memory[21427] <=  8'h63;        memory[21428] <=  8'h61;        memory[21429] <=  8'h68;        memory[21430] <=  8'h64;        memory[21431] <=  8'h75;        memory[21432] <=  8'h63;        memory[21433] <=  8'h74;        memory[21434] <=  8'h61;        memory[21435] <=  8'h64;        memory[21436] <=  8'h61;        memory[21437] <=  8'h61;        memory[21438] <=  8'h63;        memory[21439] <=  8'h61;        memory[21440] <=  8'h72;        memory[21441] <=  8'h63;        memory[21442] <=  8'h74;        memory[21443] <=  8'h72;        memory[21444] <=  8'h63;        memory[21445] <=  8'h61;        memory[21446] <=  8'h74;        memory[21447] <=  8'h72;        memory[21448] <=  8'h63;        memory[21449] <=  8'h61;        memory[21450] <=  8'h74;        memory[21451] <=  8'h63;        memory[21452] <=  8'h62;        memory[21453] <=  8'h61;        memory[21454] <=  8'h74;        memory[21455] <=  8'h62;        memory[21456] <=  8'h72;        memory[21457] <=  8'h63;        memory[21458] <=  8'h61;        memory[21459] <=  8'h74;        memory[21460] <=  8'h72;        memory[21461] <=  8'h6e;        memory[21462] <=  8'h62;        memory[21463] <=  8'h61;        memory[21464] <=  8'h63;        memory[21465] <=  8'h61;        memory[21466] <=  8'h74;        memory[21467] <=  8'h79;        memory[21468] <=  8'h73;        memory[21469] <=  8'h6e;        memory[21470] <=  8'h63;        memory[21471] <=  8'h74;        memory[21472] <=  8'h61;        memory[21473] <=  8'h6e;        memory[21474] <=  8'h62;        memory[21475] <=  8'h61;        memory[21476] <=  8'h63;        memory[21477] <=  8'h72;        memory[21478] <=  8'h6e;        memory[21479] <=  8'h74;        memory[21480] <=  8'h61;        memory[21481] <=  8'h62;        memory[21482] <=  8'h74;        memory[21483] <=  8'h6e;        memory[21484] <=  8'h61;        memory[21485] <=  8'h72;        memory[21486] <=  8'h62;        memory[21487] <=  8'h78;        memory[21488] <=  8'h74;        memory[21489] <=  8'h61;        memory[21490] <=  8'h72;        memory[21491] <=  8'h62;        memory[21492] <=  8'h61;        memory[21493] <=  8'h72;        memory[21494] <=  8'h74;        memory[21495] <=  8'h74;        memory[21496] <=  8'h62;        memory[21497] <=  8'h61;        memory[21498] <=  8'h72;        memory[21499] <=  8'h74;        memory[21500] <=  8'h78;        memory[21501] <=  8'h61;        memory[21502] <=  8'h74;        memory[21503] <=  8'h6b;        memory[21504] <=  8'h73;        memory[21505] <=  8'h68;        memory[21506] <=  8'h63;        memory[21507] <=  8'h66;        memory[21508] <=  8'h69;        memory[21509] <=  8'h77;        memory[21510] <=  8'h68;        memory[21511] <=  8'h61;        memory[21512] <=  8'h74;        memory[21513] <=  8'h61;        memory[21514] <=  8'h6e;        memory[21515] <=  8'h61;        memory[21516] <=  8'h62;        memory[21517] <=  8'h61;        memory[21518] <=  8'h63;        memory[21519] <=  8'h61;        memory[21520] <=  8'h74;        memory[21521] <=  8'h61;        memory[21522] <=  8'h62;        memory[21523] <=  8'h61;        memory[21524] <=  8'h72;        memory[21525] <=  8'h63;        memory[21526] <=  8'h61;        memory[21527] <=  8'h68;        memory[21528] <=  8'h64;        memory[21529] <=  8'h75;        memory[21530] <=  8'h63;        memory[21531] <=  8'h74;        memory[21532] <=  8'h61;        memory[21533] <=  8'h64;        memory[21534] <=  8'h61;        memory[21535] <=  8'h61;        memory[21536] <=  8'h63;        memory[21537] <=  8'h61;        memory[21538] <=  8'h72;        memory[21539] <=  8'h63;        memory[21540] <=  8'h74;        memory[21541] <=  8'h72;        memory[21542] <=  8'h63;        memory[21543] <=  8'h61;        memory[21544] <=  8'h74;        memory[21545] <=  8'h72;        memory[21546] <=  8'h63;        memory[21547] <=  8'h61;        memory[21548] <=  8'h74;        memory[21549] <=  8'h63;        memory[21550] <=  8'h62;        memory[21551] <=  8'h61;        memory[21552] <=  8'h74;        memory[21553] <=  8'h62;        memory[21554] <=  8'h72;        memory[21555] <=  8'h63;        memory[21556] <=  8'h61;        memory[21557] <=  8'h74;        memory[21558] <=  8'h72;        memory[21559] <=  8'h6e;        memory[21560] <=  8'h62;        memory[21561] <=  8'h61;        memory[21562] <=  8'h63;        memory[21563] <=  8'h61;        memory[21564] <=  8'h74;        memory[21565] <=  8'h79;        memory[21566] <=  8'h73;        memory[21567] <=  8'h6e;        memory[21568] <=  8'h63;        memory[21569] <=  8'h74;        memory[21570] <=  8'h61;        memory[21571] <=  8'h6e;        memory[21572] <=  8'h62;        memory[21573] <=  8'h61;        memory[21574] <=  8'h63;        memory[21575] <=  8'h72;        memory[21576] <=  8'h6e;        memory[21577] <=  8'h74;        memory[21578] <=  8'h61;        memory[21579] <=  8'h62;        memory[21580] <=  8'h74;        memory[21581] <=  8'h6e;        memory[21582] <=  8'h61;        memory[21583] <=  8'h72;        memory[21584] <=  8'h62;        memory[21585] <=  8'h78;        memory[21586] <=  8'h74;        memory[21587] <=  8'h61;        memory[21588] <=  8'h72;        memory[21589] <=  8'h5d;        memory[21590] <=  8'h5d;        memory[21591] <=  8'h65;        memory[21592] <=  8'h66;        memory[21593] <=  8'h77;        memory[21594] <=  8'h65;        memory[21595] <=  8'h5d;        memory[21596] <=  8'h65;        memory[21597] <=  8'h67;        memory[21598] <=  8'h73;        memory[21599] <=  8'h67;        memory[21600] <=  8'h66;        memory[21601] <=  8'h62;        memory[21602] <=  8'h61;        memory[21603] <=  8'h72;        memory[21604] <=  8'h74;        memory[21605] <=  8'h74;        memory[21606] <=  8'h62;        memory[21607] <=  8'h61;        memory[21608] <=  8'h72;        memory[21609] <=  8'h74;        memory[21610] <=  8'h78;        memory[21611] <=  8'h61;        memory[21612] <=  8'h74;        memory[21613] <=  8'h6b;        memory[21614] <=  8'h73;        memory[21615] <=  8'h68;        memory[21616] <=  8'h63;        memory[21617] <=  8'h66;        memory[21618] <=  8'h69;        memory[21619] <=  8'h77;        memory[21620] <=  8'h68;        memory[21621] <=  8'h61;        memory[21622] <=  8'h74;        memory[21623] <=  8'h61;        memory[21624] <=  8'h6e;        memory[21625] <=  8'h61;        memory[21626] <=  8'h62;        memory[21627] <=  8'h61;        memory[21628] <=  8'h63;        memory[21629] <=  8'h61;        memory[21630] <=  8'h74;        memory[21631] <=  8'h61;        memory[21632] <=  8'h62;        memory[21633] <=  8'h61;        memory[21634] <=  8'h72;        memory[21635] <=  8'h63;        memory[21636] <=  8'h61;        memory[21637] <=  8'h68;        memory[21638] <=  8'h64;        memory[21639] <=  8'h75;        memory[21640] <=  8'h63;        memory[21641] <=  8'h74;        memory[21642] <=  8'h61;        memory[21643] <=  8'h64;        memory[21644] <=  8'h61;        memory[21645] <=  8'h61;        memory[21646] <=  8'h63;        memory[21647] <=  8'h61;        memory[21648] <=  8'h72;        memory[21649] <=  8'h63;        memory[21650] <=  8'h74;        memory[21651] <=  8'h72;        memory[21652] <=  8'h63;        memory[21653] <=  8'h61;        memory[21654] <=  8'h74;        memory[21655] <=  8'h72;        memory[21656] <=  8'h63;        memory[21657] <=  8'h61;        memory[21658] <=  8'h74;        memory[21659] <=  8'h63;        memory[21660] <=  8'h62;        memory[21661] <=  8'h61;        memory[21662] <=  8'h74;        memory[21663] <=  8'h62;        memory[21664] <=  8'h72;        memory[21665] <=  8'h63;        memory[21666] <=  8'h61;        memory[21667] <=  8'h74;        memory[21668] <=  8'h72;        memory[21669] <=  8'h6e;        memory[21670] <=  8'h62;        memory[21671] <=  8'h61;        memory[21672] <=  8'h63;        memory[21673] <=  8'h61;        memory[21674] <=  8'h74;        memory[21675] <=  8'h79;        memory[21676] <=  8'h73;        memory[21677] <=  8'h6e;        memory[21678] <=  8'h63;        memory[21679] <=  8'h74;        memory[21680] <=  8'h61;        memory[21681] <=  8'h6e;        memory[21682] <=  8'h62;        memory[21683] <=  8'h61;        memory[21684] <=  8'h63;        memory[21685] <=  8'h72;        memory[21686] <=  8'h6e;        memory[21687] <=  8'h74;        memory[21688] <=  8'h61;        memory[21689] <=  8'h62;        memory[21690] <=  8'h74;        memory[21691] <=  8'h6e;        memory[21692] <=  8'h61;        memory[21693] <=  8'h72;        memory[21694] <=  8'h62;        memory[21695] <=  8'h78;        memory[21696] <=  8'h74;        memory[21697] <=  8'h61;        memory[21698] <=  8'h72;        memory[21699] <=  8'h62;        memory[21700] <=  8'h61;        memory[21701] <=  8'h72;        memory[21702] <=  8'h74;        memory[21703] <=  8'h74;        memory[21704] <=  8'h62;        memory[21705] <=  8'h61;        memory[21706] <=  8'h72;        memory[21707] <=  8'h74;        memory[21708] <=  8'h78;        memory[21709] <=  8'h61;        memory[21710] <=  8'h74;        memory[21711] <=  8'h6b;        memory[21712] <=  8'h73;        memory[21713] <=  8'h68;        memory[21714] <=  8'h63;        memory[21715] <=  8'h66;        memory[21716] <=  8'h69;        memory[21717] <=  8'h77;        memory[21718] <=  8'h68;        memory[21719] <=  8'h61;        memory[21720] <=  8'h74;        memory[21721] <=  8'h61;        memory[21722] <=  8'h6e;        memory[21723] <=  8'h61;        memory[21724] <=  8'h62;        memory[21725] <=  8'h61;        memory[21726] <=  8'h63;        memory[21727] <=  8'h61;        memory[21728] <=  8'h74;        memory[21729] <=  8'h61;        memory[21730] <=  8'h62;        memory[21731] <=  8'h61;        memory[21732] <=  8'h72;        memory[21733] <=  8'h63;        memory[21734] <=  8'h61;        memory[21735] <=  8'h68;        memory[21736] <=  8'h64;        memory[21737] <=  8'h75;        memory[21738] <=  8'h63;        memory[21739] <=  8'h74;        memory[21740] <=  8'h61;        memory[21741] <=  8'h64;        memory[21742] <=  8'h61;        memory[21743] <=  8'h61;        memory[21744] <=  8'h63;        memory[21745] <=  8'h61;        memory[21746] <=  8'h72;        memory[21747] <=  8'h63;        memory[21748] <=  8'h74;        memory[21749] <=  8'h72;        memory[21750] <=  8'h63;        memory[21751] <=  8'h61;        memory[21752] <=  8'h74;        memory[21753] <=  8'h72;        memory[21754] <=  8'h63;        memory[21755] <=  8'h61;        memory[21756] <=  8'h74;        memory[21757] <=  8'h63;        memory[21758] <=  8'h62;        memory[21759] <=  8'h61;        memory[21760] <=  8'h74;        memory[21761] <=  8'h62;        memory[21762] <=  8'h72;        memory[21763] <=  8'h63;        memory[21764] <=  8'h61;        memory[21765] <=  8'h74;        memory[21766] <=  8'h72;        memory[21767] <=  8'h6e;        memory[21768] <=  8'h62;        memory[21769] <=  8'h61;        memory[21770] <=  8'h63;        memory[21771] <=  8'h61;        memory[21772] <=  8'h74;        memory[21773] <=  8'h79;        memory[21774] <=  8'h73;        memory[21775] <=  8'h6e;        memory[21776] <=  8'h63;        memory[21777] <=  8'h74;        memory[21778] <=  8'h61;        memory[21779] <=  8'h6e;        memory[21780] <=  8'h62;        memory[21781] <=  8'h61;        memory[21782] <=  8'h63;        memory[21783] <=  8'h72;        memory[21784] <=  8'h6e;        memory[21785] <=  8'h74;        memory[21786] <=  8'h61;        memory[21787] <=  8'h62;        memory[21788] <=  8'h74;        memory[21789] <=  8'h6e;        memory[21790] <=  8'h61;        memory[21791] <=  8'h72;        memory[21792] <=  8'h62;        memory[21793] <=  8'h78;        memory[21794] <=  8'h74;        memory[21795] <=  8'h61;        memory[21796] <=  8'h72;        memory[21797] <=  8'h64;        memory[21798] <=  8'h66;        memory[21799] <=  8'h73;        memory[21800] <=  8'h67;        memory[21801] <=  8'h76;        memory[21802] <=  8'h68;        memory[21803] <=  8'h62;        memory[21804] <=  8'h6b;        memory[21805] <=  8'h6a;        memory[21806] <=  8'h6e;        memory[21807] <=  8'h6d;        memory[21808] <=  8'h62;        memory[21809] <=  8'h76;        memory[21810] <=  8'h78;        memory[21811] <=  8'h63;        memory[21812] <=  8'h73;        memory[21813] <=  8'h66;        memory[21814] <=  8'h72;        memory[21815] <=  8'h74;        memory[21816] <=  8'h79;        memory[21817] <=  8'h75;        memory[21818] <=  8'h6a;        memory[21819] <=  8'h6e;        memory[21820] <=  8'h62;        memory[21821] <=  8'h76;        memory[21822] <=  8'h63;        memory[21823] <=  8'h64;        memory[21824] <=  8'h74;        memory[21825] <=  8'h79;        memory[21826] <=  8'h75;        memory[21827] <=  8'h69;        memory[21828] <=  8'h6b;        memory[21829] <=  8'h6d;        memory[21830] <=  8'h6e;        memory[21831] <=  8'h62;        memory[21832] <=  8'h76;        memory[21833] <=  8'h63;        memory[21834] <=  8'h78;        memory[21835] <=  8'h73;        memory[21836] <=  8'h64;        memory[21837] <=  8'h72;        memory[21838] <=  8'h74;        memory[21839] <=  8'h79;        memory[21840] <=  8'h75;        memory[21841] <=  8'h69;        memory[21842] <=  8'h6b;        memory[21843] <=  8'h6d;        memory[21844] <=  8'h6e;        memory[21845] <=  8'h62;        memory[21846] <=  8'h76;        memory[21847] <=  8'h63;        memory[21848] <=  8'h73;        memory[21849] <=  8'h77;        memory[21850] <=  8'h33;        memory[21851] <=  8'h34;        memory[21852] <=  8'h35;        memory[21853] <=  8'h36;        memory[21854] <=  8'h37;        memory[21855] <=  8'h38;        memory[21856] <=  8'h69;        memory[21857] <=  8'h6b;        memory[21858] <=  8'h6d;        memory[21859] <=  8'h6e;        memory[21860] <=  8'h62;        memory[21861] <=  8'h76;        memory[21862] <=  8'h63;        memory[21863] <=  8'h64;        memory[21864] <=  8'h65;        memory[21865] <=  8'h72;        memory[21866] <=  8'h36;        memory[21867] <=  8'h37;        memory[21868] <=  8'h38;        memory[21869] <=  8'h69;        memory[21870] <=  8'h6f;        memory[21871] <=  8'h6b;        memory[21872] <=  8'h6a;        memory[21873] <=  8'h6e;        memory[21874] <=  8'h62;        memory[21875] <=  8'h76;        memory[21876] <=  8'h63;        memory[21877] <=  8'h64;        memory[21878] <=  8'h72;        memory[21879] <=  8'h74;        memory[21880] <=  8'h79;        memory[21881] <=  8'h75;        memory[21882] <=  8'h73;        memory[21883] <=  8'h6a;        memory[21884] <=  8'h63;        memory[21885] <=  8'h6e;        memory[21886] <=  8'h62;        memory[21887] <=  8'h64;        memory[21888] <=  8'h66;        memory[21889] <=  8'h73;        memory[21890] <=  8'h74;        memory[21891] <=  8'h79;        memory[21892] <=  8'h75;        memory[21893] <=  8'h61;        memory[21894] <=  8'h69;        memory[21895] <=  8'h6b;        memory[21896] <=  8'h78;        memory[21897] <=  8'h6d;        memory[21898] <=  8'h6e;        memory[21899] <=  8'h73;        memory[21900] <=  8'h6a;        memory[21901] <=  8'h6f;        memory[21902] <=  8'h64;        memory[21903] <=  8'h6c;        memory[21904] <=  8'h63;        memory[21905] <=  8'h78;        memory[21906] <=  8'h62;        memory[21907] <=  8'h61;        memory[21908] <=  8'h72;        memory[21909] <=  8'h74;        memory[21910] <=  8'h78;        memory[21911] <=  8'h61;        memory[21912] <=  8'h74;        memory[21913] <=  8'h6b;        memory[21914] <=  8'h73;        memory[21915] <=  8'h68;        memory[21916] <=  8'h63;        memory[21917] <=  8'h66;        memory[21918] <=  8'h69;        memory[21919] <=  8'h77;        memory[21920] <=  8'h68;        memory[21921] <=  8'h61;        memory[21922] <=  8'h74;        memory[21923] <=  8'h61;        memory[21924] <=  8'h6e;        memory[21925] <=  8'h61;        memory[21926] <=  8'h62;        memory[21927] <=  8'h61;        memory[21928] <=  8'h63;        memory[21929] <=  8'h61;        memory[21930] <=  8'h74;        memory[21931] <=  8'h61;        memory[21932] <=  8'h62;        memory[21933] <=  8'h61;        memory[21934] <=  8'h72;        memory[21935] <=  8'h63;        memory[21936] <=  8'h61;        memory[21937] <=  8'h68;        memory[21938] <=  8'h64;        memory[21939] <=  8'h75;        memory[21940] <=  8'h63;        memory[21941] <=  8'h74;        memory[21942] <=  8'h61;        memory[21943] <=  8'h64;        memory[21944] <=  8'h61;        memory[21945] <=  8'h61;        memory[21946] <=  8'h63;        memory[21947] <=  8'h61;        memory[21948] <=  8'h72;        memory[21949] <=  8'h62;        memory[21950] <=  8'h61;        memory[21951] <=  8'h72;        memory[21952] <=  8'h74;        memory[21953] <=  8'h78;        memory[21954] <=  8'h61;        memory[21955] <=  8'h74;        memory[21956] <=  8'h6b;        memory[21957] <=  8'h73;        memory[21958] <=  8'h68;        memory[21959] <=  8'h63;        memory[21960] <=  8'h66;        memory[21961] <=  8'h69;        memory[21962] <=  8'h77;        memory[21963] <=  8'h68;        memory[21964] <=  8'h61;        memory[21965] <=  8'h74;        memory[21966] <=  8'h61;        memory[21967] <=  8'h6e;        memory[21968] <=  8'h61;        memory[21969] <=  8'h62;        memory[21970] <=  8'h61;        memory[21971] <=  8'h63;        memory[21972] <=  8'h61;        memory[21973] <=  8'h74;        memory[21974] <=  8'h61;        memory[21975] <=  8'h62;        memory[21976] <=  8'h61;        memory[21977] <=  8'h72;        memory[21978] <=  8'h63;        memory[21979] <=  8'h61;        memory[21980] <=  8'h68;        memory[21981] <=  8'h64;        memory[21982] <=  8'h75;        memory[21983] <=  8'h63;        memory[21984] <=  8'h74;        memory[21985] <=  8'h61;        memory[21986] <=  8'h64;        memory[21987] <=  8'h61;        memory[21988] <=  8'h61;        memory[21989] <=  8'h63;        memory[21990] <=  8'h61;        memory[21991] <=  8'h72;        memory[21992] <=  8'h62;        memory[21993] <=  8'h61;        memory[21994] <=  8'h72;        memory[21995] <=  8'h74;        memory[21996] <=  8'h78;        memory[21997] <=  8'h61;        memory[21998] <=  8'h74;        memory[21999] <=  8'h6b;        memory[22000] <=  8'h73;        memory[22001] <=  8'h68;        memory[22002] <=  8'h63;        memory[22003] <=  8'h66;        memory[22004] <=  8'h69;        memory[22005] <=  8'h77;        memory[22006] <=  8'h68;        memory[22007] <=  8'h61;        memory[22008] <=  8'h74;        memory[22009] <=  8'h61;        memory[22010] <=  8'h6e;        memory[22011] <=  8'h61;        memory[22012] <=  8'h62;        memory[22013] <=  8'h61;        memory[22014] <=  8'h63;        memory[22015] <=  8'h61;        memory[22016] <=  8'h74;        memory[22017] <=  8'h61;        memory[22018] <=  8'h62;        memory[22019] <=  8'h61;        memory[22020] <=  8'h72;        memory[22021] <=  8'h63;        memory[22022] <=  8'h61;        memory[22023] <=  8'h68;        memory[22024] <=  8'h64;        memory[22025] <=  8'h75;        memory[22026] <=  8'h63;        memory[22027] <=  8'h74;        memory[22028] <=  8'h61;        memory[22029] <=  8'h64;        memory[22030] <=  8'h61;        memory[22031] <=  8'h61;        memory[22032] <=  8'h63;        memory[22033] <=  8'h61;        memory[22034] <=  8'h72;        memory[22035] <=  8'h62;        memory[22036] <=  8'h61;        memory[22037] <=  8'h72;        memory[22038] <=  8'h74;        memory[22039] <=  8'h78;        memory[22040] <=  8'h61;        memory[22041] <=  8'h74;        memory[22042] <=  8'h6b;        memory[22043] <=  8'h73;        memory[22044] <=  8'h68;        memory[22045] <=  8'h63;        memory[22046] <=  8'h66;        memory[22047] <=  8'h69;        memory[22048] <=  8'h77;        memory[22049] <=  8'h68;        memory[22050] <=  8'h61;        memory[22051] <=  8'h74;        memory[22052] <=  8'h61;        memory[22053] <=  8'h6e;        memory[22054] <=  8'h61;        memory[22055] <=  8'h62;        memory[22056] <=  8'h61;        memory[22057] <=  8'h63;        memory[22058] <=  8'h61;        memory[22059] <=  8'h74;        memory[22060] <=  8'h61;        memory[22061] <=  8'h62;        memory[22062] <=  8'h61;        memory[22063] <=  8'h72;        memory[22064] <=  8'h63;        memory[22065] <=  8'h61;        memory[22066] <=  8'h68;        memory[22067] <=  8'h64;        memory[22068] <=  8'h75;        memory[22069] <=  8'h63;        memory[22070] <=  8'h74;        memory[22071] <=  8'h61;        memory[22072] <=  8'h64;        memory[22073] <=  8'h61;        memory[22074] <=  8'h61;        memory[22075] <=  8'h63;        memory[22076] <=  8'h61;        memory[22077] <=  8'h72;        memory[22078] <=  8'h62;        memory[22079] <=  8'h61;        memory[22080] <=  8'h72;        memory[22081] <=  8'h74;        memory[22082] <=  8'h78;        memory[22083] <=  8'h61;        memory[22084] <=  8'h74;        memory[22085] <=  8'h6b;        memory[22086] <=  8'h73;        memory[22087] <=  8'h68;        memory[22088] <=  8'h63;        memory[22089] <=  8'h66;        memory[22090] <=  8'h69;        memory[22091] <=  8'h77;        memory[22092] <=  8'h68;        memory[22093] <=  8'h61;        memory[22094] <=  8'h74;        memory[22095] <=  8'h61;        memory[22096] <=  8'h6e;        memory[22097] <=  8'h61;        memory[22098] <=  8'h62;        memory[22099] <=  8'h61;        memory[22100] <=  8'h63;        memory[22101] <=  8'h61;        memory[22102] <=  8'h74;        memory[22103] <=  8'h61;        memory[22104] <=  8'h62;        memory[22105] <=  8'h61;        memory[22106] <=  8'h72;        memory[22107] <=  8'h63;        memory[22108] <=  8'h61;        memory[22109] <=  8'h68;        memory[22110] <=  8'h64;        memory[22111] <=  8'h75;        memory[22112] <=  8'h63;        memory[22113] <=  8'h74;        memory[22114] <=  8'h61;        memory[22115] <=  8'h64;        memory[22116] <=  8'h61;        memory[22117] <=  8'h61;        memory[22118] <=  8'h63;        memory[22119] <=  8'h61;        memory[22120] <=  8'h72;        memory[22121] <=  8'h62;        memory[22122] <=  8'h61;        memory[22123] <=  8'h72;        memory[22124] <=  8'h74;        memory[22125] <=  8'h78;        memory[22126] <=  8'h61;        memory[22127] <=  8'h74;        memory[22128] <=  8'h6b;        memory[22129] <=  8'h73;        memory[22130] <=  8'h68;        memory[22131] <=  8'h63;        memory[22132] <=  8'h66;        memory[22133] <=  8'h69;        memory[22134] <=  8'h77;        memory[22135] <=  8'h68;        memory[22136] <=  8'h61;        memory[22137] <=  8'h74;        memory[22138] <=  8'h61;        memory[22139] <=  8'h6e;        memory[22140] <=  8'h61;        memory[22141] <=  8'h62;        memory[22142] <=  8'h61;        memory[22143] <=  8'h63;        memory[22144] <=  8'h61;        memory[22145] <=  8'h74;        memory[22146] <=  8'h61;        memory[22147] <=  8'h62;        memory[22148] <=  8'h61;        memory[22149] <=  8'h72;        memory[22150] <=  8'h63;        memory[22151] <=  8'h61;        memory[22152] <=  8'h68;        memory[22153] <=  8'h64;        memory[22154] <=  8'h75;        memory[22155] <=  8'h63;        memory[22156] <=  8'h74;        memory[22157] <=  8'h61;        memory[22158] <=  8'h64;        memory[22159] <=  8'h61;        memory[22160] <=  8'h61;        memory[22161] <=  8'h63;        memory[22162] <=  8'h61;        memory[22163] <=  8'h72;        memory[22164] <=  8'h62;        memory[22165] <=  8'h61;        memory[22166] <=  8'h72;        memory[22167] <=  8'h74;        memory[22168] <=  8'h78;        memory[22169] <=  8'h61;        memory[22170] <=  8'h74;        memory[22171] <=  8'h6b;        memory[22172] <=  8'h73;        memory[22173] <=  8'h68;        memory[22174] <=  8'h63;        memory[22175] <=  8'h66;        memory[22176] <=  8'h69;        memory[22177] <=  8'h77;        memory[22178] <=  8'h68;        memory[22179] <=  8'h61;        memory[22180] <=  8'h74;        memory[22181] <=  8'h61;        memory[22182] <=  8'h6e;        memory[22183] <=  8'h61;        memory[22184] <=  8'h62;        memory[22185] <=  8'h61;        memory[22186] <=  8'h63;        memory[22187] <=  8'h61;        memory[22188] <=  8'h74;        memory[22189] <=  8'h61;        memory[22190] <=  8'h62;        memory[22191] <=  8'h61;        memory[22192] <=  8'h72;        memory[22193] <=  8'h63;        memory[22194] <=  8'h61;        memory[22195] <=  8'h68;        memory[22196] <=  8'h64;        memory[22197] <=  8'h75;        memory[22198] <=  8'h63;        memory[22199] <=  8'h74;        memory[22200] <=  8'h61;        memory[22201] <=  8'h64;        memory[22202] <=  8'h61;        memory[22203] <=  8'h61;        memory[22204] <=  8'h63;        memory[22205] <=  8'h61;        memory[22206] <=  8'h72;        memory[22207] <=  8'h62;        memory[22208] <=  8'h61;        memory[22209] <=  8'h72;        memory[22210] <=  8'h74;        memory[22211] <=  8'h78;        memory[22212] <=  8'h61;        memory[22213] <=  8'h74;        memory[22214] <=  8'h6b;        memory[22215] <=  8'h73;        memory[22216] <=  8'h68;        memory[22217] <=  8'h63;        memory[22218] <=  8'h66;        memory[22219] <=  8'h69;        memory[22220] <=  8'h77;        memory[22221] <=  8'h68;        memory[22222] <=  8'h61;        memory[22223] <=  8'h74;        memory[22224] <=  8'h61;        memory[22225] <=  8'h6e;        memory[22226] <=  8'h61;        memory[22227] <=  8'h62;        memory[22228] <=  8'h61;        memory[22229] <=  8'h63;        memory[22230] <=  8'h61;        memory[22231] <=  8'h74;        memory[22232] <=  8'h61;        memory[22233] <=  8'h62;        memory[22234] <=  8'h61;        memory[22235] <=  8'h72;        memory[22236] <=  8'h63;        memory[22237] <=  8'h61;        memory[22238] <=  8'h68;        memory[22239] <=  8'h64;        memory[22240] <=  8'h75;        memory[22241] <=  8'h63;        memory[22242] <=  8'h74;        memory[22243] <=  8'h61;        memory[22244] <=  8'h64;        memory[22245] <=  8'h61;        memory[22246] <=  8'h61;        memory[22247] <=  8'h63;        memory[22248] <=  8'h61;        memory[22249] <=  8'h72;        memory[22250] <=  8'h62;        memory[22251] <=  8'h61;        memory[22252] <=  8'h72;        memory[22253] <=  8'h74;        memory[22254] <=  8'h78;        memory[22255] <=  8'h61;        memory[22256] <=  8'h74;        memory[22257] <=  8'h6b;        memory[22258] <=  8'h73;        memory[22259] <=  8'h68;        memory[22260] <=  8'h63;        memory[22261] <=  8'h66;        memory[22262] <=  8'h69;        memory[22263] <=  8'h77;        memory[22264] <=  8'h68;        memory[22265] <=  8'h61;        memory[22266] <=  8'h74;        memory[22267] <=  8'h61;        memory[22268] <=  8'h6e;        memory[22269] <=  8'h61;        memory[22270] <=  8'h62;        memory[22271] <=  8'h61;        memory[22272] <=  8'h63;        memory[22273] <=  8'h61;        memory[22274] <=  8'h74;        memory[22275] <=  8'h61;        memory[22276] <=  8'h62;        memory[22277] <=  8'h61;        memory[22278] <=  8'h72;        memory[22279] <=  8'h63;        memory[22280] <=  8'h61;        memory[22281] <=  8'h68;        memory[22282] <=  8'h64;        memory[22283] <=  8'h75;        memory[22284] <=  8'h63;        memory[22285] <=  8'h74;        memory[22286] <=  8'h61;        memory[22287] <=  8'h64;        memory[22288] <=  8'h61;        memory[22289] <=  8'h61;        memory[22290] <=  8'h63;        memory[22291] <=  8'h61;        memory[22292] <=  8'h72;        memory[22293] <=  8'h62;        memory[22294] <=  8'h61;        memory[22295] <=  8'h72;        memory[22296] <=  8'h74;        memory[22297] <=  8'h74;        memory[22298] <=  8'h62;        memory[22299] <=  8'h61;        memory[22300] <=  8'h72;        memory[22301] <=  8'h74;        memory[22302] <=  8'h78;        memory[22303] <=  8'h61;        memory[22304] <=  8'h74;        memory[22305] <=  8'h6b;        memory[22306] <=  8'h73;        memory[22307] <=  8'h68;        memory[22308] <=  8'h63;        memory[22309] <=  8'h66;        memory[22310] <=  8'h69;        memory[22311] <=  8'h77;        memory[22312] <=  8'h68;        memory[22313] <=  8'h61;        memory[22314] <=  8'h74;        memory[22315] <=  8'h61;        memory[22316] <=  8'h6e;        memory[22317] <=  8'h61;        memory[22318] <=  8'h62;        memory[22319] <=  8'h61;        memory[22320] <=  8'h63;        memory[22321] <=  8'h61;        memory[22322] <=  8'h74;        memory[22323] <=  8'h61;        memory[22324] <=  8'h62;        memory[22325] <=  8'h61;        memory[22326] <=  8'h72;        memory[22327] <=  8'h63;        memory[22328] <=  8'h61;        memory[22329] <=  8'h68;        memory[22330] <=  8'h64;        memory[22331] <=  8'h75;        memory[22332] <=  8'h63;        memory[22333] <=  8'h74;        memory[22334] <=  8'h61;        memory[22335] <=  8'h64;        memory[22336] <=  8'h61;        memory[22337] <=  8'h61;        memory[22338] <=  8'h63;        memory[22339] <=  8'h61;        memory[22340] <=  8'h72;        memory[22341] <=  8'h63;        memory[22342] <=  8'h74;        memory[22343] <=  8'h72;        memory[22344] <=  8'h63;        memory[22345] <=  8'h61;        memory[22346] <=  8'h74;        memory[22347] <=  8'h72;        memory[22348] <=  8'h63;        memory[22349] <=  8'h61;        memory[22350] <=  8'h74;        memory[22351] <=  8'h63;        memory[22352] <=  8'h62;        memory[22353] <=  8'h61;        memory[22354] <=  8'h74;        memory[22355] <=  8'h62;        memory[22356] <=  8'h72;        memory[22357] <=  8'h63;        memory[22358] <=  8'h61;        memory[22359] <=  8'h72;        memory[22360] <=  8'h62;        memory[22361] <=  8'h78;        memory[22362] <=  8'h74;        memory[22363] <=  8'h61;        memory[22364] <=  8'h72;        memory[22365] <=  8'h64;        memory[22366] <=  8'h66;        memory[22367] <=  8'h73;        memory[22368] <=  8'h67;        memory[22369] <=  8'h76;        memory[22370] <=  8'h68;        memory[22371] <=  8'h62;        memory[22372] <=  8'h6b;        memory[22373] <=  8'h6a;        memory[22374] <=  8'h6e;        memory[22375] <=  8'h6d;        memory[22376] <=  8'h62;        memory[22377] <=  8'h76;        memory[22378] <=  8'h78;        memory[22379] <=  8'h63;        memory[22380] <=  8'h73;        memory[22381] <=  8'h66;        memory[22382] <=  8'h72;        memory[22383] <=  8'h74;        memory[22384] <=  8'h79;        memory[22385] <=  8'h75;        memory[22386] <=  8'h6a;        memory[22387] <=  8'h6e;        memory[22388] <=  8'h62;        memory[22389] <=  8'h76;        memory[22390] <=  8'h63;        memory[22391] <=  8'h64;        memory[22392] <=  8'h74;        memory[22393] <=  8'h79;        memory[22394] <=  8'h75;        memory[22395] <=  8'h69;        memory[22396] <=  8'h6b;        memory[22397] <=  8'h6d;        memory[22398] <=  8'h6e;        memory[22399] <=  8'h62;        memory[22400] <=  8'h76;        memory[22401] <=  8'h63;        memory[22402] <=  8'h78;        memory[22403] <=  8'h73;        memory[22404] <=  8'h64;        memory[22405] <=  8'h72;        memory[22406] <=  8'h74;        memory[22407] <=  8'h79;        memory[22408] <=  8'h75;        memory[22409] <=  8'h69;        memory[22410] <=  8'h6b;        memory[22411] <=  8'h6d;        memory[22412] <=  8'h6e;        memory[22413] <=  8'h62;        memory[22414] <=  8'h76;        memory[22415] <=  8'h63;        memory[22416] <=  8'h73;        memory[22417] <=  8'h77;        memory[22418] <=  8'h33;        memory[22419] <=  8'h34;        memory[22420] <=  8'h35;        memory[22421] <=  8'h36;        memory[22422] <=  8'h37;        memory[22423] <=  8'h38;        memory[22424] <=  8'h69;        memory[22425] <=  8'h6b;        memory[22426] <=  8'h6d;        memory[22427] <=  8'h6e;        memory[22428] <=  8'h62;        memory[22429] <=  8'h76;        memory[22430] <=  8'h63;        memory[22431] <=  8'h64;        memory[22432] <=  8'h65;        memory[22433] <=  8'h72;        memory[22434] <=  8'h36;        memory[22435] <=  8'h37;        memory[22436] <=  8'h38;        memory[22437] <=  8'h69;        memory[22438] <=  8'h6f;        memory[22439] <=  8'h6b;        memory[22440] <=  8'h6a;        memory[22441] <=  8'h6e;        memory[22442] <=  8'h62;        memory[22443] <=  8'h76;        memory[22444] <=  8'h63;        memory[22445] <=  8'h64;        memory[22446] <=  8'h72;        memory[22447] <=  8'h74;        memory[22448] <=  8'h79;        memory[22449] <=  8'h75;        memory[22450] <=  8'h73;        memory[22451] <=  8'h6a;        memory[22452] <=  8'h63;        memory[22453] <=  8'h6e;        memory[22454] <=  8'h62;        memory[22455] <=  8'h64;        memory[22456] <=  8'h66;        memory[22457] <=  8'h73;        memory[22458] <=  8'h74;        memory[22459] <=  8'h79;        memory[22460] <=  8'h75;        memory[22461] <=  8'h61;        memory[22462] <=  8'h69;        memory[22463] <=  8'h6b;        memory[22464] <=  8'h78;        memory[22465] <=  8'h6d;        memory[22466] <=  8'h6e;        memory[22467] <=  8'h73;        memory[22468] <=  8'h6a;        memory[22469] <=  8'h6f;        memory[22470] <=  8'h64;        memory[22471] <=  8'h6c;        memory[22472] <=  8'h63;        memory[22473] <=  8'h78;        memory[22474] <=  8'h2c;        memory[22475] <=  8'h6d;        memory[22476] <=  8'h73;        memory[22477] <=  8'h6b;        memory[22478] <=  8'h64;        memory[22479] <=  8'h6c;        memory[22480] <=  8'h70;        memory[22481] <=  8'h5b;        memory[22482] <=  8'h3b;        memory[22483] <=  8'h73;        memory[22484] <=  8'h6c;        memory[22485] <=  8'h64;        memory[22486] <=  8'h70;        memory[22487] <=  8'h76;        memory[22488] <=  8'h63;        memory[22489] <=  8'h5b;        memory[22490] <=  8'h78;        memory[22491] <=  8'h76;        memory[22492] <=  8'h63;        memory[22493] <=  8'h5b;        memory[22494] <=  8'h78;        memory[22495] <=  8'h70;        memory[22496] <=  8'h6f;        memory[22497] <=  8'h20;        memory[22498] <=  8'h62;        memory[22499] <=  8'h61;        memory[22500] <=  8'h72;        memory[22501] <=  8'h74;        memory[22502] <=  8'h74;        memory[22503] <=  8'h62;        memory[22504] <=  8'h61;        memory[22505] <=  8'h72;        memory[22506] <=  8'h74;        memory[22507] <=  8'h78;        memory[22508] <=  8'h61;        memory[22509] <=  8'h74;        memory[22510] <=  8'h6b;        memory[22511] <=  8'h73;        memory[22512] <=  8'h68;        memory[22513] <=  8'h63;        memory[22514] <=  8'h66;        memory[22515] <=  8'h69;        memory[22516] <=  8'h77;        memory[22517] <=  8'h68;        memory[22518] <=  8'h61;        memory[22519] <=  8'h69;        memory[22520] <=  8'h6a;        memory[22521] <=  8'h78;        memory[22522] <=  8'h5d;        memory[22523] <=  8'h65;        memory[22524] <=  8'h6b;        memory[22525] <=  8'h6f;        memory[22526] <=  8'h39;        memory[22527] <=  8'h64;        memory[22528] <=  8'h75;        memory[22529] <=  8'h38;        memory[22530] <=  8'h79;        memory[22531] <=  8'h20;        memory[22532] <=  8'h37;        memory[22533] <=  8'h63;        memory[22534] <=  8'h67;        memory[22535] <=  8'h78;        memory[22536] <=  8'h63;        memory[22537] <=  8'h75;        memory[22538] <=  8'h68;        memory[22539] <=  8'h69;        memory[22540] <=  8'h6a;        memory[22541] <=  8'h77;        memory[22542] <=  8'h69;        memory[22543] <=  8'h64;        memory[22544] <=  8'h66;        memory[22545] <=  8'h68;        memory[22546] <=  8'h75;        memory[22547] <=  8'h76;        memory[22548] <=  8'h64;        memory[22549] <=  8'h62;        memory[22550] <=  8'h66;        memory[22551] <=  8'h6a;        memory[22552] <=  8'h6e;        memory[22553] <=  8'h6b;        memory[22554] <=  8'h6a;        memory[22555] <=  8'h65;        memory[22556] <=  8'h38;        memory[22557] <=  8'h66;        memory[22558] <=  8'h37;        memory[22559] <=  8'h67;        memory[22560] <=  8'h79;        memory[22561] <=  8'h76;        memory[22562] <=  8'h63;        memory[22563] <=  8'h68;        memory[22564] <=  8'h69;        memory[22565] <=  8'h6a;        memory[22566] <=  8'h33;        memory[22567] <=  8'h65;        memory[22568] <=  8'h67;        memory[22569] <=  8'h79;        memory[22570] <=  8'h72;        memory[22571] <=  8'h64;        memory[22572] <=  8'h62;        memory[22573] <=  8'h6e;        memory[22574] <=  8'h63;        memory[22575] <=  8'h7a;        memory[22576] <=  8'h6a;        memory[22577] <=  8'h6f;        memory[22578] <=  8'h66;        memory[22579] <=  8'h78;        memory[22580] <=  8'h6a;        memory[22581] <=  8'h69;        memory[22582] <=  8'h63;        memory[22583] <=  8'h68;        memory[22584] <=  8'h62;        memory[22585] <=  8'h6e;        memory[22586] <=  8'h6d;        memory[22587] <=  8'h63;        memory[22588] <=  8'h73;        memory[22589] <=  8'h6c;        memory[22590] <=  8'h6b;        memory[22591] <=  8'h6a;        memory[22592] <=  8'h69;        memory[22593] <=  8'h68;        memory[22594] <=  8'h76;        memory[22595] <=  8'h75;        memory[22596] <=  8'h69;        memory[22597] <=  8'h64;        memory[22598] <=  8'h68;        memory[22599] <=  8'h75;        memory[22600] <=  8'h67;        memory[22601] <=  8'h79;        memory[22602] <=  8'h62;        memory[22603] <=  8'h68;        memory[22604] <=  8'h65;        memory[22605] <=  8'h6a;        memory[22606] <=  8'h72;        memory[22607] <=  8'h6b;        memory[22608] <=  8'h6a;        memory[22609] <=  8'h6f;        memory[22610] <=  8'h64;        memory[22611] <=  8'h67;        memory[22612] <=  8'h69;        memory[22613] <=  8'h75;        memory[22614] <=  8'h69;        memory[22615] <=  8'h67;        memory[22616] <=  8'h76;        memory[22617] <=  8'h79;        memory[22618] <=  8'h75;        memory[22619] <=  8'h67;        memory[22620] <=  8'h78;        memory[22621] <=  8'h68;        memory[22622] <=  8'h63;        memory[22623] <=  8'h20;        memory[22624] <=  8'h20;        memory[22625] <=  8'h20;        memory[22626] <=  8'h78;        memory[22627] <=  8'h76;        memory[22628] <=  8'h20;        memory[22629] <=  8'h63;        memory[22630] <=  8'h78;        memory[22631] <=  8'h67;        memory[22632] <=  8'h79;        memory[22633] <=  8'h63;        memory[22634] <=  8'h75;        memory[22635] <=  8'h68;        memory[22636] <=  8'h6a;        memory[22637] <=  8'h6b;        memory[22638] <=  8'h61;        memory[22639] <=  8'h6c;        memory[22640] <=  8'h78;        memory[22641] <=  8'h76;        memory[22642] <=  8'h70;        memory[22643] <=  8'h6f;        memory[22644] <=  8'h69;        memory[22645] <=  8'h6a;        memory[22646] <=  8'h69;        memory[22647] <=  8'h68;        memory[22648] <=  8'h6a;        memory[22649] <=  8'h62;        memory[22650] <=  8'h77;        memory[22651] <=  8'h65;        memory[22652] <=  8'h6e;        memory[22653] <=  8'h61;        memory[22654] <=  8'h66;        memory[22655] <=  8'h6d;        memory[22656] <=  8'h64;        memory[22657] <=  8'h6b;        memory[22658] <=  8'h6d;        memory[22659] <=  8'h76;        memory[22660] <=  8'h6c;        memory[22661] <=  8'h63;        memory[22662] <=  8'h6f;        memory[22663] <=  8'h64;        memory[22664] <=  8'h69;        memory[22665] <=  8'h75;        memory[22666] <=  8'h68;        memory[22667] <=  8'h73;        memory[22668] <=  8'h66;        memory[22669] <=  8'h65;        memory[22670] <=  8'h62;        memory[22671] <=  8'h6e;        memory[22672] <=  8'h64;        memory[22673] <=  8'h73;        memory[22674] <=  8'h63;        memory[22675] <=  8'h6b;        memory[22676] <=  8'h20;        memory[22677] <=  8'h78;        memory[22678] <=  8'h6a;        memory[22679] <=  8'h78;        memory[22680] <=  8'h63;        memory[22681] <=  8'h73;        memory[22682] <=  8'h64;        memory[22683] <=  8'h66;        memory[22684] <=  8'h6b;        memory[22685] <=  8'h64;        memory[22686] <=  8'h6e;        memory[22687] <=  8'h6d;        memory[22688] <=  8'h64;        memory[22689] <=  8'h73;        memory[22690] <=  8'h63;        memory[22691] <=  8'h6b;        memory[22692] <=  8'h78;        memory[22693] <=  8'h6c;        memory[22694] <=  8'h6f;        memory[22695] <=  8'h66;        memory[22696] <=  8'h6a;        memory[22697] <=  8'h69;        memory[22698] <=  8'h61;        memory[22699] <=  8'h62;        memory[22700] <=  8'h6e;        memory[22701] <=  8'h20;        memory[22702] <=  8'h78;        memory[22703] <=  8'h6b;        memory[22704] <=  8'h6d;        memory[22705] <=  8'h20;        memory[22706] <=  8'h6f;        memory[22707] <=  8'h63;        memory[22708] <=  8'h76;        memory[22709] <=  8'h73;        memory[22710] <=  8'h64;        memory[22711] <=  8'h69;        memory[22712] <=  8'h66;        memory[22713] <=  8'h68;        memory[22714] <=  8'h65;        memory[22715] <=  8'h71;        memory[22716] <=  8'h6a;        memory[22717] <=  8'h77;        memory[22718] <=  8'h62;        memory[22719] <=  8'h65;        memory[22720] <=  8'h6e;        memory[22721] <=  8'h20;        memory[22722] <=  8'h6d;        memory[22723] <=  8'h64;        memory[22724] <=  8'h73;        memory[22725] <=  8'h6c;        memory[22726] <=  8'h76;        memory[22727] <=  8'h6b;        memory[22728] <=  8'h63;        memory[22729] <=  8'h78;        memory[22730] <=  8'h20;        memory[22731] <=  8'h6f;        memory[22732] <=  8'h78;        memory[22733] <=  8'h69;        memory[22734] <=  8'h63;        memory[22735] <=  8'h6a;        memory[22736] <=  8'h76;        memory[22737] <=  8'h64;        memory[22738] <=  8'h66;        memory[22739] <=  8'h65;        memory[22740] <=  8'h71;        memory[22741] <=  8'h6e;        memory[22742] <=  8'h20;        memory[22743] <=  8'h64;        memory[22744] <=  8'h6d;        memory[22745] <=  8'h73;        memory[22746] <=  8'h6c;        memory[22747] <=  8'h63;        memory[22748] <=  8'h78;        memory[22749] <=  8'h6b;        memory[22750] <=  8'h20;        memory[22751] <=  8'h6f;        memory[22752] <=  8'h78;        memory[22753] <=  8'h63;        memory[22754] <=  8'h76;        memory[22755] <=  8'h6a;        memory[22756] <=  8'h64;        memory[22757] <=  8'h62;        memory[22758] <=  8'h71;        memory[22759] <=  8'h77;        memory[22760] <=  8'h65;        memory[22761] <=  8'h6e;        memory[22762] <=  8'h6d;        memory[22763] <=  8'h64;        memory[22764] <=  8'h6c;        memory[22765] <=  8'h73;        memory[22766] <=  8'h2c;        memory[22767] <=  8'h76;        memory[22768] <=  8'h63;        memory[22769] <=  8'h78;        memory[22770] <=  8'h20;        memory[22771] <=  8'h63;        memory[22772] <=  8'h6f;        memory[22773] <=  8'h69;        memory[22774] <=  8'h76;        memory[22775] <=  8'h68;        memory[22776] <=  8'h73;        memory[22777] <=  8'h64;        memory[22778] <=  8'h62;        memory[22779] <=  8'h71;        memory[22780] <=  8'h77;        memory[22781] <=  8'h65;        memory[22782] <=  8'h6e;        memory[22783] <=  8'h64;        memory[22784] <=  8'h6b;        memory[22785] <=  8'h73;        memory[22786] <=  8'h76;        memory[22787] <=  8'h6f;        memory[22788] <=  8'h63;        memory[22789] <=  8'h20;        memory[22790] <=  8'h76;        memory[22791] <=  8'h69;        memory[22792] <=  8'h75;        memory[22793] <=  8'h69;        memory[22794] <=  8'h68;        memory[22795] <=  8'h63;        memory[22796] <=  8'h78;        memory[22797] <=  8'h69;        memory[22798] <=  8'h6f;        memory[22799] <=  8'h76;        memory[22800] <=  8'h73;        memory[22801] <=  8'h64;        memory[22802] <=  8'h61;        memory[22803] <=  8'h64;        memory[22804] <=  8'h6e;        memory[22805] <=  8'h77;        memory[22806] <=  8'h71;        memory[22807] <=  8'h6b;        memory[22808] <=  8'h6c;        memory[22809] <=  8'h73;        memory[22810] <=  8'h76;        memory[22811] <=  8'h6e;        memory[22812] <=  8'h62;        memory[22813] <=  8'h20;        memory[22814] <=  8'h64;        memory[22815] <=  8'h66;        memory[22816] <=  8'h6a;        memory[22817] <=  8'h6b;        memory[22818] <=  8'h71;        memory[22819] <=  8'h64;        memory[22820] <=  8'h77;        memory[22821] <=  8'h65;        memory[22822] <=  8'h6e;        memory[22823] <=  8'h62;        memory[22824] <=  8'h20;        memory[22825] <=  8'h64;        memory[22826] <=  8'h73;        memory[22827] <=  8'h76;        memory[22828] <=  8'h68;        memory[22829] <=  8'h64;        memory[22830] <=  8'h61;        memory[22831] <=  8'h71;        memory[22832] <=  8'h77;        memory[22833] <=  8'h6a;        memory[22834] <=  8'h65;        memory[22835] <=  8'h6e;        memory[22836] <=  8'h64;        memory[22837] <=  8'h20;        memory[22838] <=  8'h61;        memory[22839] <=  8'h63;        memory[22840] <=  8'h62;        memory[22841] <=  8'h68;        memory[22842] <=  8'h64;        memory[22843] <=  8'h61;        memory[22844] <=  8'h77;        memory[22845] <=  8'h71;        memory[22846] <=  8'h6e;        memory[22847] <=  8'h20;        memory[22848] <=  8'h62;        memory[22849] <=  8'h73;        memory[22850] <=  8'h76;        memory[22851] <=  8'h61;        memory[22852] <=  8'h67;        memory[22853] <=  8'h76;        memory[22854] <=  8'h68;        memory[22855] <=  8'h67;        memory[22856] <=  8'h61;        memory[22857] <=  8'h73;        memory[22858] <=  8'h6a;        memory[22859] <=  8'h6b;        memory[22860] <=  8'h63;        memory[22861] <=  8'h78;        memory[22862] <=  8'h76;        memory[22863] <=  8'h6e;        memory[22864] <=  8'h73;        memory[22865] <=  8'h64;        memory[22866] <=  8'h20;        memory[22867] <=  8'h66;        memory[22868] <=  8'h62;        memory[22869] <=  8'h64;        memory[22870] <=  8'h61;        memory[22871] <=  8'h73;        memory[22872] <=  8'h76;        memory[22873] <=  8'h67;        memory[22874] <=  8'h63;        memory[22875] <=  8'h79;        memory[22876] <=  8'h7a;        memory[22877] <=  8'h78;        memory[22878] <=  8'h79;        memory[22879] <=  8'h75;        memory[22880] <=  8'h20;        memory[22881] <=  8'h69;        memory[22882] <=  8'h6a;        memory[22883] <=  8'h64;        memory[22884] <=  8'h66;        memory[22885] <=  8'h6b;        memory[22886] <=  8'h61;        memory[22887] <=  8'h64;        memory[22888] <=  8'h63;        memory[22889] <=  8'h78;        memory[22890] <=  8'h68;        memory[22891] <=  8'h20;        memory[22892] <=  8'h67;        memory[22893] <=  8'h61;        memory[22894] <=  8'h68;        memory[22895] <=  8'h75;        memory[22896] <=  8'h64;        memory[22897] <=  8'h73;        memory[22898] <=  8'h69;        memory[22899] <=  8'h6a;        memory[22900] <=  8'h61;        memory[22901] <=  8'h6b;        memory[22902] <=  8'h63;        memory[22903] <=  8'h62;        memory[22904] <=  8'h61;        memory[22905] <=  8'h72;        memory[22906] <=  8'h73;        memory[22907] <=  8'h68;        memory[22908] <=  8'h64;        memory[22909] <=  8'h66;        memory[22910] <=  8'h67;        memory[22911] <=  8'h73;        memory[22912] <=  8'h68;        memory[22913] <=  8'h64;        memory[22914] <=  8'h66;        memory[22915] <=  8'h68;        memory[22916] <=  8'h64;        memory[22917] <=  8'h6a;        memory[22918] <=  8'h68;        memory[22919] <=  8'h62;        memory[22920] <=  8'h67;        memory[22921] <=  8'h63;        memory[22922] <=  8'h61;        memory[22923] <=  8'h66;        memory[22924] <=  8'h73;        memory[22925] <=  8'h79;        memory[22926] <=  8'h67;        memory[22927] <=  8'h6b;        memory[22928] <=  8'h75;        memory[22929] <=  8'h64;        memory[22930] <=  8'h68;        memory[22931] <=  8'h62;        memory[22932] <=  8'h77;        memory[22933] <=  8'h76;        memory[22934] <=  8'h67;        memory[22935] <=  8'h61;        memory[22936] <=  8'h66;        memory[22937] <=  8'h64;        memory[22938] <=  8'h74;        memory[22939] <=  8'h75;        memory[22940] <=  8'h66;        memory[22941] <=  8'h79;        memory[22942] <=  8'h67;        memory[22943] <=  8'h69;        memory[22944] <=  8'h75;        memory[22945] <=  8'h68;        memory[22946] <=  8'h6c;        memory[22947] <=  8'h6a;        memory[22948] <=  8'h62;        memory[22949] <=  8'h6b;        memory[22950] <=  8'h68;        memory[22951] <=  8'h76;        memory[22952] <=  8'h67;        memory[22953] <=  8'h63;        memory[22954] <=  8'h66;        memory[22955] <=  8'h78;        memory[22956] <=  8'h64;        memory[22957] <=  8'h74;        memory[22958] <=  8'h75;        memory[22959] <=  8'h79;        memory[22960] <=  8'h69;        memory[22961] <=  8'h75;        memory[22962] <=  8'h68;        memory[22963] <=  8'h6c;        memory[22964] <=  8'h6a;        memory[22965] <=  8'h6b;        memory[22966] <=  8'h67;        memory[22967] <=  8'h6a;        memory[22968] <=  8'h63;        memory[22969] <=  8'h66;        memory[22970] <=  8'h68;        memory[22971] <=  8'h64;        memory[22972] <=  8'h67;        memory[22973] <=  8'h72;        memory[22974] <=  8'h79;        memory[22975] <=  8'h74;        memory[22976] <=  8'h66;        memory[22977] <=  8'h75;        memory[22978] <=  8'h79;        memory[22979] <=  8'h69;        memory[22980] <=  8'h68;        memory[22981] <=  8'h6c;        memory[22982] <=  8'h62;        memory[22983] <=  8'h6d;        memory[22984] <=  8'h76;        memory[22985] <=  8'h6e;        memory[22986] <=  8'h63;        memory[22987] <=  8'h66;        memory[22988] <=  8'h68;        memory[22989] <=  8'h64;        memory[22990] <=  8'h74;        memory[22991] <=  8'h75;        memory[22992] <=  8'h67;        memory[22993] <=  8'h79;        memory[22994] <=  8'h69;        memory[22995] <=  8'h68;        memory[22996] <=  8'h75;        memory[22997] <=  8'h6a;        memory[22998] <=  8'h6c;        memory[22999] <=  8'h62;        memory[23000] <=  8'h6d;        memory[23001] <=  8'h76;        memory[23002] <=  8'h6e;        memory[23003] <=  8'h63;        memory[23004] <=  8'h66;        memory[23005] <=  8'h68;        memory[23006] <=  8'h67;        memory[23007] <=  8'h79;        memory[23008] <=  8'h68;        memory[23009] <=  8'h75;        memory[23010] <=  8'h6a;        memory[23011] <=  8'h6e;        memory[23012] <=  8'h2c;        memory[23013] <=  8'h62;        memory[23014] <=  8'h6e;        memory[23015] <=  8'h6d;        memory[23016] <=  8'h76;        memory[23017] <=  8'h6e;        memory[23018] <=  8'h63;        memory[23019] <=  8'h66;        memory[23020] <=  8'h68;        memory[23021] <=  8'h74;        memory[23022] <=  8'h79;        memory[23023] <=  8'h69;        memory[23024] <=  8'h75;        memory[23025] <=  8'h6c;        memory[23026] <=  8'h6a;        memory[23027] <=  8'h62;        memory[23028] <=  8'h6d;        memory[23029] <=  8'h76;        memory[23030] <=  8'h6e;        memory[23031] <=  8'h63;        memory[23032] <=  8'h66;        memory[23033] <=  8'h74;        memory[23034] <=  8'h75;        memory[23035] <=  8'h79;        memory[23036] <=  8'h69;        memory[23037] <=  8'h68;        memory[23038] <=  8'h6b;        memory[23039] <=  8'h62;        memory[23040] <=  8'h76;        memory[23041] <=  8'h63;        memory[23042] <=  8'h66;        memory[23043] <=  8'h67;        memory[23044] <=  8'h74;        memory[23045] <=  8'h75;        memory[23046] <=  8'h79;        memory[23047] <=  8'h69;        memory[23048] <=  8'h75;        memory[23049] <=  8'h68;        memory[23050] <=  8'h6a;        memory[23051] <=  8'h6b;        memory[23052] <=  8'h62;        memory[23053] <=  8'h76;        memory[23054] <=  8'h63;        memory[23055] <=  8'h66;        memory[23056] <=  8'h74;        memory[23057] <=  8'h75;        memory[23058] <=  8'h79;        memory[23059] <=  8'h69;        memory[23060] <=  8'h75;        memory[23061] <=  8'h6a;        memory[23062] <=  8'h6b;        memory[23063] <=  8'h6e;        memory[23064] <=  8'h62;        memory[23065] <=  8'h76;        memory[23066] <=  8'h67;        memory[23067] <=  8'h66;        memory[23068] <=  8'h74;        memory[23069] <=  8'h79;        memory[23070] <=  8'h75;        memory[23071] <=  8'h75;        memory[23072] <=  8'h69;        memory[23073] <=  8'h6a;        memory[23074] <=  8'h6b;        memory[23075] <=  8'h68;        memory[23076] <=  8'h62;        memory[23077] <=  8'h6a;        memory[23078] <=  8'h67;        memory[23079] <=  8'h68;        memory[23080] <=  8'h66;        memory[23081] <=  8'h79;        memory[23082] <=  8'h74;        memory[23083] <=  8'h79;        memory[23084] <=  8'h69;        memory[23085] <=  8'h75;        memory[23086] <=  8'h64;        memory[23087] <=  8'h6a;        memory[23088] <=  8'h6b;        memory[23089] <=  8'h68;        memory[23090] <=  8'h63;        memory[23091] <=  8'h7a;        memory[23092] <=  8'h67;        memory[23093] <=  8'h68;        memory[23094] <=  8'h74;        memory[23095] <=  8'h75;        memory[23096] <=  8'h79;        memory[23097] <=  8'h69;        memory[23098] <=  8'h61;        memory[23099] <=  8'h73;        memory[23100] <=  8'h75;        memory[23101] <=  8'h6a;        memory[23102] <=  8'h6b;        memory[23103] <=  8'h62;        memory[23104] <=  8'h6e;        memory[23105] <=  8'h61;        memory[23106] <=  8'h76;        memory[23107] <=  8'h63;        memory[23108] <=  8'h66;        memory[23109] <=  8'h68;        memory[23110] <=  8'h75;        memory[23111] <=  8'h61;        memory[23112] <=  8'h73;        memory[23113] <=  8'h79;        memory[23114] <=  8'h64;        memory[23115] <=  8'h75;        memory[23116] <=  8'h69;        memory[23117] <=  8'h6a;        memory[23118] <=  8'h61;        memory[23119] <=  8'h6b;        memory[23120] <=  8'h62;        memory[23121] <=  8'h63;        memory[23122] <=  8'h78;        memory[23123] <=  8'h68;        memory[23124] <=  8'h67;        memory[23125] <=  8'h79;        memory[23126] <=  8'h75;        memory[23127] <=  8'h7a;        memory[23128] <=  8'h63;        memory[23129] <=  8'h61;        memory[23130] <=  8'h73;        memory[23131] <=  8'h69;        memory[23132] <=  8'h75;        memory[23133] <=  8'h6f;        memory[23134] <=  8'h69;        memory[23135] <=  8'h6a;        memory[23136] <=  8'h61;        memory[23137] <=  8'h6c;        memory[23138] <=  8'h63;        memory[23139] <=  8'h78;        memory[23140] <=  8'h62;        memory[23141] <=  8'h63;        memory[23142] <=  8'h20;        memory[23143] <=  8'h6e;        memory[23144] <=  8'h76;        memory[23145] <=  8'h63;        memory[23146] <=  8'h61;        memory[23147] <=  8'h64;        memory[23148] <=  8'h73;        memory[23149] <=  8'h67;        memory[23150] <=  8'h79;        memory[23151] <=  8'h68;        memory[23152] <=  8'h75;        memory[23153] <=  8'h61;        memory[23154] <=  8'h6a;        memory[23155] <=  8'h6b;        memory[23156] <=  8'h78;        memory[23157] <=  8'h62;        memory[23158] <=  8'h20;        memory[23159] <=  8'h6e;        memory[23160] <=  8'h76;        memory[23161] <=  8'h63;        memory[23162] <=  8'h61;        memory[23163] <=  8'h73;        memory[23164] <=  8'h67;        memory[23165] <=  8'h68;        memory[23166] <=  8'h75;        memory[23167] <=  8'h6a;        memory[23168] <=  8'h6c;        memory[23169] <=  8'h6b;        memory[23170] <=  8'h63;        memory[23171] <=  8'h78;        memory[23172] <=  8'h20;        memory[23173] <=  8'h6a;        memory[23174] <=  8'h6b;        memory[23175] <=  8'h68;        memory[23176] <=  8'h61;        memory[23177] <=  8'h73;        memory[23178] <=  8'h76;        memory[23179] <=  8'h64;        memory[23180] <=  8'h6e;        memory[23181] <=  8'h20;        memory[23182] <=  8'h62;        memory[23183] <=  8'h6e;        memory[23184] <=  8'h6d;        memory[23185] <=  8'h6b;        memory[23186] <=  8'h77;        memory[23187] <=  8'h64;        memory[23188] <=  8'h6f;        memory[23189] <=  8'h77;        memory[23190] <=  8'h69;        memory[23191] <=  8'h6f;        memory[23192] <=  8'h75;        memory[23193] <=  8'h69;        memory[23194] <=  8'h68;        memory[23195] <=  8'h62;        memory[23196] <=  8'h6e;        memory[23197] <=  8'h6b;        memory[23198] <=  8'h77;        memory[23199] <=  8'h69;        memory[23200] <=  8'h6f;        memory[23201] <=  8'h75;        memory[23202] <=  8'h71;        memory[23203] <=  8'h69;        memory[23204] <=  8'h79;        memory[23205] <=  8'h67;        memory[23206] <=  8'h6a;        memory[23207] <=  8'h64;        memory[23208] <=  8'h61;        memory[23209] <=  8'h76;        memory[23210] <=  8'h62;        memory[23211] <=  8'h6e;        memory[23212] <=  8'h6b;        memory[23213] <=  8'h6f;        memory[23214] <=  8'h70;        memory[23215] <=  8'h64;        memory[23216] <=  8'h76;        memory[23217] <=  8'h69;        memory[23218] <=  8'h6f;        memory[23219] <=  8'h75;        memory[23220] <=  8'h69;        memory[23221] <=  8'h48;        memory[23222] <=  8'h42;        memory[23223] <=  8'h6b;        memory[23224] <=  8'h64;        memory[23225] <=  8'h6e;        memory[23226] <=  8'h6c;        memory[23227] <=  8'h71;        memory[23228] <=  8'h6b;        memory[23229] <=  8'h6d;        memory[23230] <=  8'h6a;        memory[23231] <=  8'h70;        memory[23232] <=  8'h69;        memory[23233] <=  8'h6f;        memory[23234] <=  8'h68;        memory[23235] <=  8'h65;        memory[23236] <=  8'h66;        memory[23237] <=  8'h75;        memory[23238] <=  8'h67;        memory[23239] <=  8'h69;        memory[23240] <=  8'h73;        memory[23241] <=  8'h61;        memory[23242] <=  8'h62;        memory[23243] <=  8'h64;        memory[23244] <=  8'h6b;        memory[23245] <=  8'h6a;        memory[23246] <=  8'h6b;        memory[23247] <=  8'h6c;        memory[23248] <=  8'h6a;        memory[23249] <=  8'h69;        memory[23250] <=  8'h73;        memory[23251] <=  8'h6f;        memory[23252] <=  8'h71;        memory[23253] <=  8'h68;        memory[23254] <=  8'h77;        memory[23255] <=  8'h67;        memory[23256] <=  8'h69;        memory[23257] <=  8'h79;        memory[23258] <=  8'h6a;        memory[23259] <=  8'h64;        memory[23260] <=  8'h76;        memory[23261] <=  8'h62;        memory[23262] <=  8'h6e;        memory[23263] <=  8'h61;        memory[23264] <=  8'h73;        memory[23265] <=  8'h66;        memory[23266] <=  8'h6c;        memory[23267] <=  8'h6b;        memory[23268] <=  8'h64;        memory[23269] <=  8'h6a;        memory[23270] <=  8'h68;        memory[23271] <=  8'h63;        memory[23272] <=  8'h67;        memory[23273] <=  8'h6a;        memory[23274] <=  8'h76;        memory[23275] <=  8'h73;        memory[23276] <=  8'h64;        memory[23277] <=  8'h62;        memory[23278] <=  8'h62;        memory[23279] <=  8'h61;        memory[23280] <=  8'h72;        memory[23281] <=  8'h62;        memory[23282] <=  8'h62;        memory[23283] <=  8'h73;        memory[23284] <=  8'h62;        memory[23285] <=  8'h67;        memory[23286] <=  8'h73;        memory[23287] <=  8'h66;        memory[23288] <=  8'h67;        memory[23289] <=  8'h61;        memory[23290] <=  8'h68;        memory[23291] <=  8'h66;        memory[23292] <=  8'h73;        memory[23293] <=  8'h68;        memory[23294] <=  8'h61;        memory[23295] <=  8'h66;        memory[23296] <=  8'h73;        memory[23297] <=  8'h66;        memory[23298] <=  8'h68;        memory[23299] <=  8'h61;        memory[23300] <=  8'h69;        memory[23301] <=  8'h64;        memory[23302] <=  8'h75;        memory[23303] <=  8'h67;        memory[23304] <=  8'h64;        memory[23305] <=  8'h77;        memory[23306] <=  8'h62;        memory[23307] <=  8'h61;        memory[23308] <=  8'h62;        memory[23309] <=  8'h72;        memory[23310] <=  8'h62;        memory[23311] <=  8'h61;        memory[23312] <=  8'h62;        memory[23313] <=  8'h62;        memory[23314] <=  8'h74;        memory[23315] <=  8'h62;        memory[23316] <=  8'h62;        memory[23317] <=  8'h62;        memory[23318] <=  8'h62;        memory[23319] <=  8'h62;        memory[23320] <=  8'h62;        memory[23321] <=  8'h62;        memory[23322] <=  8'h62;        memory[23323] <=  8'h61;        memory[23324] <=  8'h62;        memory[23325] <=  8'h62;        memory[23326] <=  8'h72;        memory[23327] <=  8'h74;        memory[23328] <=  8'h62;        memory[23329] <=  8'h62;        memory[23330] <=  8'h61;        memory[23331] <=  8'h62;        memory[23332] <=  8'h72;        memory[23333] <=  8'h62;        memory[23334] <=  8'h74;        memory[23335] <=  8'h62;        memory[23336] <=  8'h62;        memory[23337] <=  8'h62;        memory[23338] <=  8'h63;        memory[23339] <=  8'h61;        memory[23340] <=  8'h72;        memory[23341] <=  8'h74;        memory[23342] <=  8'h73;        memory[23343] <=  8'h62;        memory[23344] <=  8'h61;        memory[23345] <=  8'h72;        memory[23346] <=  8'h74;        memory[23347] <=  8'h74;        memory[23348] <=  8'h62;        memory[23349] <=  8'h61;        memory[23350] <=  8'h72;        memory[23351] <=  8'h74;        memory[23352] <=  8'h78;        memory[23353] <=  8'h61;        memory[23354] <=  8'h74;        memory[23355] <=  8'h6b;        memory[23356] <=  8'h73;        memory[23357] <=  8'h68;        memory[23358] <=  8'h63;        memory[23359] <=  8'h66;        memory[23360] <=  8'h69;        memory[23361] <=  8'h77;        memory[23362] <=  8'h68;        memory[23363] <=  8'h61;        memory[23364] <=  8'h74;        memory[23365] <=  8'h61;        memory[23366] <=  8'h6e;        memory[23367] <=  8'h61;        memory[23368] <=  8'h62;        memory[23369] <=  8'h61;        memory[23370] <=  8'h63;        memory[23371] <=  8'h61;        memory[23372] <=  8'h74;        memory[23373] <=  8'h61;        memory[23374] <=  8'h62;        memory[23375] <=  8'h61;        memory[23376] <=  8'h72;        memory[23377] <=  8'h63;        memory[23378] <=  8'h61;        memory[23379] <=  8'h68;        memory[23380] <=  8'h64;        memory[23381] <=  8'h75;        memory[23382] <=  8'h63;        memory[23383] <=  8'h74;        memory[23384] <=  8'h61;        memory[23385] <=  8'h64;        memory[23386] <=  8'h61;        memory[23387] <=  8'h61;        memory[23388] <=  8'h63;        memory[23389] <=  8'h61;        memory[23390] <=  8'h72;        memory[23391] <=  8'h63;        memory[23392] <=  8'h74;        memory[23393] <=  8'h72;        memory[23394] <=  8'h63;        memory[23395] <=  8'h61;        memory[23396] <=  8'h74;        memory[23397] <=  8'h72;        memory[23398] <=  8'h63;        memory[23399] <=  8'h61;        memory[23400] <=  8'h74;        memory[23401] <=  8'h63;        memory[23402] <=  8'h62;        memory[23403] <=  8'h61;        memory[23404] <=  8'h74;        memory[23405] <=  8'h62;        memory[23406] <=  8'h72;        memory[23407] <=  8'h63;        memory[23408] <=  8'h61;        memory[23409] <=  8'h74;        memory[23410] <=  8'h72;        memory[23411] <=  8'h6e;        memory[23412] <=  8'h62;        memory[23413] <=  8'h61;        memory[23414] <=  8'h63;        memory[23415] <=  8'h61;        memory[23416] <=  8'h74;        memory[23417] <=  8'h79;        memory[23418] <=  8'h73;        memory[23419] <=  8'h6e;        memory[23420] <=  8'h63;        memory[23421] <=  8'h74;        memory[23422] <=  8'h61;        memory[23423] <=  8'h6e;        memory[23424] <=  8'h62;        memory[23425] <=  8'h61;        memory[23426] <=  8'h63;        memory[23427] <=  8'h72;        memory[23428] <=  8'h6e;        memory[23429] <=  8'h74;        memory[23430] <=  8'h61;        memory[23431] <=  8'h62;        memory[23432] <=  8'h74;        memory[23433] <=  8'h6e;        memory[23434] <=  8'h61;        memory[23435] <=  8'h72;        memory[23436] <=  8'h62;        memory[23437] <=  8'h78;        memory[23438] <=  8'h74;        memory[23439] <=  8'h61;        memory[23440] <=  8'h72;        memory[23441] <=  8'h62;        memory[23442] <=  8'h61;        memory[23443] <=  8'h72;        memory[23444] <=  8'h74;        memory[23445] <=  8'h74;        memory[23446] <=  8'h62;        memory[23447] <=  8'h61;        memory[23448] <=  8'h72;        memory[23449] <=  8'h74;        memory[23450] <=  8'h78;        memory[23451] <=  8'h61;        memory[23452] <=  8'h74;        memory[23453] <=  8'h6b;        memory[23454] <=  8'h73;        memory[23455] <=  8'h68;        memory[23456] <=  8'h63;        memory[23457] <=  8'h66;        memory[23458] <=  8'h69;        memory[23459] <=  8'h77;        memory[23460] <=  8'h68;        memory[23461] <=  8'h61;        memory[23462] <=  8'h74;        memory[23463] <=  8'h61;        memory[23464] <=  8'h6e;        memory[23465] <=  8'h61;        memory[23466] <=  8'h62;        memory[23467] <=  8'h61;        memory[23468] <=  8'h63;        memory[23469] <=  8'h61;        memory[23470] <=  8'h74;        memory[23471] <=  8'h61;        memory[23472] <=  8'h62;        memory[23473] <=  8'h61;        memory[23474] <=  8'h72;        memory[23475] <=  8'h63;        memory[23476] <=  8'h61;        memory[23477] <=  8'h68;        memory[23478] <=  8'h64;        memory[23479] <=  8'h75;        memory[23480] <=  8'h63;        memory[23481] <=  8'h74;        memory[23482] <=  8'h61;        memory[23483] <=  8'h64;        memory[23484] <=  8'h61;        memory[23485] <=  8'h61;        memory[23486] <=  8'h63;        memory[23487] <=  8'h61;        memory[23488] <=  8'h72;        memory[23489] <=  8'h63;        memory[23490] <=  8'h74;        memory[23491] <=  8'h72;        memory[23492] <=  8'h63;        memory[23493] <=  8'h61;        memory[23494] <=  8'h74;        memory[23495] <=  8'h72;        memory[23496] <=  8'h63;        memory[23497] <=  8'h61;        memory[23498] <=  8'h74;        memory[23499] <=  8'h63;        memory[23500] <=  8'h62;        memory[23501] <=  8'h61;        memory[23502] <=  8'h74;        memory[23503] <=  8'h62;        memory[23504] <=  8'h72;        memory[23505] <=  8'h63;        memory[23506] <=  8'h61;        memory[23507] <=  8'h74;        memory[23508] <=  8'h72;        memory[23509] <=  8'h6e;        memory[23510] <=  8'h62;        memory[23511] <=  8'h61;        memory[23512] <=  8'h63;        memory[23513] <=  8'h61;        memory[23514] <=  8'h74;        memory[23515] <=  8'h79;        memory[23516] <=  8'h73;        memory[23517] <=  8'h6e;        memory[23518] <=  8'h63;        memory[23519] <=  8'h74;        memory[23520] <=  8'h61;        memory[23521] <=  8'h6e;        memory[23522] <=  8'h62;        memory[23523] <=  8'h61;        memory[23524] <=  8'h63;        memory[23525] <=  8'h72;        memory[23526] <=  8'h6e;        memory[23527] <=  8'h74;        memory[23528] <=  8'h61;        memory[23529] <=  8'h62;        memory[23530] <=  8'h74;        memory[23531] <=  8'h6e;        memory[23532] <=  8'h61;        memory[23533] <=  8'h72;        memory[23534] <=  8'h62;        memory[23535] <=  8'h78;        memory[23536] <=  8'h74;        memory[23537] <=  8'h61;        memory[23538] <=  8'h72;        memory[23539] <=  8'h62;        memory[23540] <=  8'h61;        memory[23541] <=  8'h72;        memory[23542] <=  8'h74;        memory[23543] <=  8'h74;        memory[23544] <=  8'h62;        memory[23545] <=  8'h61;        memory[23546] <=  8'h72;        memory[23547] <=  8'h74;        memory[23548] <=  8'h78;        memory[23549] <=  8'h61;        memory[23550] <=  8'h74;        memory[23551] <=  8'h6b;        memory[23552] <=  8'h73;        memory[23553] <=  8'h68;        memory[23554] <=  8'h63;        memory[23555] <=  8'h66;        memory[23556] <=  8'h69;        memory[23557] <=  8'h77;        memory[23558] <=  8'h68;        memory[23559] <=  8'h61;        memory[23560] <=  8'h74;        memory[23561] <=  8'h61;        memory[23562] <=  8'h6e;        memory[23563] <=  8'h61;        memory[23564] <=  8'h62;        memory[23565] <=  8'h61;        memory[23566] <=  8'h63;        memory[23567] <=  8'h61;        memory[23568] <=  8'h74;        memory[23569] <=  8'h61;        memory[23570] <=  8'h62;        memory[23571] <=  8'h61;        memory[23572] <=  8'h72;        memory[23573] <=  8'h63;        memory[23574] <=  8'h61;        memory[23575] <=  8'h68;        memory[23576] <=  8'h64;        memory[23577] <=  8'h75;        memory[23578] <=  8'h63;        memory[23579] <=  8'h74;        memory[23580] <=  8'h61;        memory[23581] <=  8'h64;        memory[23582] <=  8'h61;        memory[23583] <=  8'h61;        memory[23584] <=  8'h63;        memory[23585] <=  8'h61;        memory[23586] <=  8'h72;        memory[23587] <=  8'h63;        memory[23588] <=  8'h74;        memory[23589] <=  8'h72;        memory[23590] <=  8'h63;        memory[23591] <=  8'h61;        memory[23592] <=  8'h74;        memory[23593] <=  8'h72;        memory[23594] <=  8'h63;        memory[23595] <=  8'h61;        memory[23596] <=  8'h74;        memory[23597] <=  8'h63;        memory[23598] <=  8'h62;        memory[23599] <=  8'h61;        memory[23600] <=  8'h74;        memory[23601] <=  8'h62;        memory[23602] <=  8'h72;        memory[23603] <=  8'h63;        memory[23604] <=  8'h61;        memory[23605] <=  8'h74;        memory[23606] <=  8'h72;        memory[23607] <=  8'h6e;        memory[23608] <=  8'h62;        memory[23609] <=  8'h61;        memory[23610] <=  8'h63;        memory[23611] <=  8'h61;        memory[23612] <=  8'h74;        memory[23613] <=  8'h79;        memory[23614] <=  8'h73;        memory[23615] <=  8'h6e;        memory[23616] <=  8'h63;        memory[23617] <=  8'h74;        memory[23618] <=  8'h61;        memory[23619] <=  8'h6e;        memory[23620] <=  8'h62;        memory[23621] <=  8'h61;        memory[23622] <=  8'h63;        memory[23623] <=  8'h72;        memory[23624] <=  8'h6e;        memory[23625] <=  8'h74;        memory[23626] <=  8'h61;        memory[23627] <=  8'h62;        memory[23628] <=  8'h74;        memory[23629] <=  8'h6e;        memory[23630] <=  8'h61;        memory[23631] <=  8'h72;        memory[23632] <=  8'h62;        memory[23633] <=  8'h78;        memory[23634] <=  8'h74;        memory[23635] <=  8'h61;        memory[23636] <=  8'h72;        memory[23637] <=  8'h5d;        memory[23638] <=  8'h5d;        memory[23639] <=  8'h65;        memory[23640] <=  8'h66;        memory[23641] <=  8'h77;        memory[23642] <=  8'h65;        memory[23643] <=  8'h5d;        memory[23644] <=  8'h65;        memory[23645] <=  8'h67;        memory[23646] <=  8'h73;        memory[23647] <=  8'h67;        memory[23648] <=  8'h66;        memory[23649] <=  8'h62;        memory[23650] <=  8'h61;        memory[23651] <=  8'h72;        memory[23652] <=  8'h74;        memory[23653] <=  8'h74;        memory[23654] <=  8'h62;        memory[23655] <=  8'h61;        memory[23656] <=  8'h72;        memory[23657] <=  8'h74;        memory[23658] <=  8'h78;        memory[23659] <=  8'h61;        memory[23660] <=  8'h74;        memory[23661] <=  8'h6b;        memory[23662] <=  8'h73;        memory[23663] <=  8'h68;        memory[23664] <=  8'h63;        memory[23665] <=  8'h66;        memory[23666] <=  8'h69;        memory[23667] <=  8'h77;        memory[23668] <=  8'h68;        memory[23669] <=  8'h61;        memory[23670] <=  8'h74;        memory[23671] <=  8'h61;        memory[23672] <=  8'h6e;        memory[23673] <=  8'h61;        memory[23674] <=  8'h62;        memory[23675] <=  8'h61;        memory[23676] <=  8'h63;        memory[23677] <=  8'h61;        memory[23678] <=  8'h74;        memory[23679] <=  8'h61;        memory[23680] <=  8'h62;        memory[23681] <=  8'h61;        memory[23682] <=  8'h72;        memory[23683] <=  8'h63;        memory[23684] <=  8'h61;        memory[23685] <=  8'h68;        memory[23686] <=  8'h64;        memory[23687] <=  8'h75;        memory[23688] <=  8'h63;        memory[23689] <=  8'h74;        memory[23690] <=  8'h61;        memory[23691] <=  8'h64;        memory[23692] <=  8'h61;        memory[23693] <=  8'h61;        memory[23694] <=  8'h63;        memory[23695] <=  8'h61;        memory[23696] <=  8'h72;        memory[23697] <=  8'h63;        memory[23698] <=  8'h74;        memory[23699] <=  8'h72;        memory[23700] <=  8'h63;        memory[23701] <=  8'h61;        memory[23702] <=  8'h74;        memory[23703] <=  8'h72;        memory[23704] <=  8'h63;        memory[23705] <=  8'h61;        memory[23706] <=  8'h74;        memory[23707] <=  8'h63;        memory[23708] <=  8'h62;        memory[23709] <=  8'h61;        memory[23710] <=  8'h74;        memory[23711] <=  8'h62;        memory[23712] <=  8'h72;        memory[23713] <=  8'h63;        memory[23714] <=  8'h61;        memory[23715] <=  8'h74;        memory[23716] <=  8'h72;        memory[23717] <=  8'h6e;        memory[23718] <=  8'h62;        memory[23719] <=  8'h61;        memory[23720] <=  8'h63;        memory[23721] <=  8'h61;        memory[23722] <=  8'h74;        memory[23723] <=  8'h79;        memory[23724] <=  8'h73;        memory[23725] <=  8'h6e;        memory[23726] <=  8'h63;        memory[23727] <=  8'h74;        memory[23728] <=  8'h61;        memory[23729] <=  8'h6e;        memory[23730] <=  8'h62;        memory[23731] <=  8'h61;        memory[23732] <=  8'h63;        memory[23733] <=  8'h72;        memory[23734] <=  8'h6e;        memory[23735] <=  8'h74;        memory[23736] <=  8'h61;        memory[23737] <=  8'h62;        memory[23738] <=  8'h74;        memory[23739] <=  8'h6e;        memory[23740] <=  8'h61;        memory[23741] <=  8'h72;        memory[23742] <=  8'h62;        memory[23743] <=  8'h78;        memory[23744] <=  8'h74;        memory[23745] <=  8'h61;        memory[23746] <=  8'h72;        memory[23747] <=  8'h62;        memory[23748] <=  8'h61;        memory[23749] <=  8'h72;        memory[23750] <=  8'h74;        memory[23751] <=  8'h74;        memory[23752] <=  8'h62;        memory[23753] <=  8'h61;        memory[23754] <=  8'h72;        memory[23755] <=  8'h74;        memory[23756] <=  8'h78;        memory[23757] <=  8'h61;        memory[23758] <=  8'h74;        memory[23759] <=  8'h6b;        memory[23760] <=  8'h73;        memory[23761] <=  8'h68;        memory[23762] <=  8'h63;        memory[23763] <=  8'h66;        memory[23764] <=  8'h69;        memory[23765] <=  8'h77;        memory[23766] <=  8'h68;        memory[23767] <=  8'h61;        memory[23768] <=  8'h74;        memory[23769] <=  8'h61;        memory[23770] <=  8'h6e;        memory[23771] <=  8'h61;        memory[23772] <=  8'h62;        memory[23773] <=  8'h61;        memory[23774] <=  8'h63;        memory[23775] <=  8'h61;        memory[23776] <=  8'h74;        memory[23777] <=  8'h61;        memory[23778] <=  8'h62;        memory[23779] <=  8'h61;        memory[23780] <=  8'h72;        memory[23781] <=  8'h63;        memory[23782] <=  8'h61;        memory[23783] <=  8'h68;        memory[23784] <=  8'h64;        memory[23785] <=  8'h75;        memory[23786] <=  8'h63;        memory[23787] <=  8'h74;        memory[23788] <=  8'h61;        memory[23789] <=  8'h64;        memory[23790] <=  8'h61;        memory[23791] <=  8'h61;        memory[23792] <=  8'h63;        memory[23793] <=  8'h61;        memory[23794] <=  8'h72;        memory[23795] <=  8'h63;        memory[23796] <=  8'h74;        memory[23797] <=  8'h72;        memory[23798] <=  8'h63;        memory[23799] <=  8'h61;        memory[23800] <=  8'h74;        memory[23801] <=  8'h72;        memory[23802] <=  8'h63;        memory[23803] <=  8'h61;        memory[23804] <=  8'h74;        memory[23805] <=  8'h63;        memory[23806] <=  8'h62;        memory[23807] <=  8'h61;        memory[23808] <=  8'h74;        memory[23809] <=  8'h62;        memory[23810] <=  8'h72;        memory[23811] <=  8'h63;        memory[23812] <=  8'h61;        memory[23813] <=  8'h74;        memory[23814] <=  8'h72;        memory[23815] <=  8'h6e;        memory[23816] <=  8'h62;        memory[23817] <=  8'h61;        memory[23818] <=  8'h63;        memory[23819] <=  8'h61;        memory[23820] <=  8'h74;        memory[23821] <=  8'h79;        memory[23822] <=  8'h73;        memory[23823] <=  8'h6e;        memory[23824] <=  8'h63;        memory[23825] <=  8'h74;        memory[23826] <=  8'h61;        memory[23827] <=  8'h6e;        memory[23828] <=  8'h62;        memory[23829] <=  8'h61;        memory[23830] <=  8'h63;        memory[23831] <=  8'h72;        memory[23832] <=  8'h6e;        memory[23833] <=  8'h74;        memory[23834] <=  8'h61;        memory[23835] <=  8'h62;        memory[23836] <=  8'h74;        memory[23837] <=  8'h6e;        memory[23838] <=  8'h61;        memory[23839] <=  8'h72;        memory[23840] <=  8'h62;        memory[23841] <=  8'h78;        memory[23842] <=  8'h74;        memory[23843] <=  8'h61;        memory[23844] <=  8'h72;        memory[23845] <=  8'h64;        memory[23846] <=  8'h66;        memory[23847] <=  8'h73;        memory[23848] <=  8'h67;        memory[23849] <=  8'h76;        memory[23850] <=  8'h68;        memory[23851] <=  8'h62;        memory[23852] <=  8'h6b;        memory[23853] <=  8'h6a;        memory[23854] <=  8'h6e;        memory[23855] <=  8'h6d;        memory[23856] <=  8'h62;        memory[23857] <=  8'h76;        memory[23858] <=  8'h78;        memory[23859] <=  8'h63;        memory[23860] <=  8'h73;        memory[23861] <=  8'h66;        memory[23862] <=  8'h72;        memory[23863] <=  8'h74;        memory[23864] <=  8'h79;        memory[23865] <=  8'h75;        memory[23866] <=  8'h6a;        memory[23867] <=  8'h6e;        memory[23868] <=  8'h62;        memory[23869] <=  8'h76;        memory[23870] <=  8'h63;        memory[23871] <=  8'h64;        memory[23872] <=  8'h74;        memory[23873] <=  8'h79;        memory[23874] <=  8'h75;        memory[23875] <=  8'h69;        memory[23876] <=  8'h6b;        memory[23877] <=  8'h6d;        memory[23878] <=  8'h6e;        memory[23879] <=  8'h62;        memory[23880] <=  8'h76;        memory[23881] <=  8'h63;        memory[23882] <=  8'h78;        memory[23883] <=  8'h73;        memory[23884] <=  8'h64;        memory[23885] <=  8'h72;        memory[23886] <=  8'h74;        memory[23887] <=  8'h79;        memory[23888] <=  8'h75;        memory[23889] <=  8'h69;        memory[23890] <=  8'h6b;        memory[23891] <=  8'h6d;        memory[23892] <=  8'h6e;        memory[23893] <=  8'h62;        memory[23894] <=  8'h76;        memory[23895] <=  8'h63;        memory[23896] <=  8'h73;        memory[23897] <=  8'h77;        memory[23898] <=  8'h33;        memory[23899] <=  8'h34;        memory[23900] <=  8'h35;        memory[23901] <=  8'h36;        memory[23902] <=  8'h37;        memory[23903] <=  8'h38;        memory[23904] <=  8'h69;        memory[23905] <=  8'h6b;        memory[23906] <=  8'h6d;        memory[23907] <=  8'h6e;        memory[23908] <=  8'h62;        memory[23909] <=  8'h76;        memory[23910] <=  8'h63;        memory[23911] <=  8'h64;        memory[23912] <=  8'h65;        memory[23913] <=  8'h72;        memory[23914] <=  8'h36;        memory[23915] <=  8'h37;        memory[23916] <=  8'h38;        memory[23917] <=  8'h69;        memory[23918] <=  8'h6f;        memory[23919] <=  8'h6b;        memory[23920] <=  8'h6a;        memory[23921] <=  8'h6e;        memory[23922] <=  8'h62;        memory[23923] <=  8'h76;        memory[23924] <=  8'h63;        memory[23925] <=  8'h64;        memory[23926] <=  8'h72;        memory[23927] <=  8'h74;        memory[23928] <=  8'h79;        memory[23929] <=  8'h75;        memory[23930] <=  8'h73;        memory[23931] <=  8'h6a;        memory[23932] <=  8'h63;        memory[23933] <=  8'h6e;        memory[23934] <=  8'h62;        memory[23935] <=  8'h64;        memory[23936] <=  8'h66;        memory[23937] <=  8'h73;        memory[23938] <=  8'h74;        memory[23939] <=  8'h79;        memory[23940] <=  8'h75;        memory[23941] <=  8'h61;        memory[23942] <=  8'h69;        memory[23943] <=  8'h6b;        memory[23944] <=  8'h78;        memory[23945] <=  8'h6d;        memory[23946] <=  8'h6e;        memory[23947] <=  8'h73;        memory[23948] <=  8'h6a;        memory[23949] <=  8'h6f;        memory[23950] <=  8'h64;        memory[23951] <=  8'h6c;        memory[23952] <=  8'h63;        memory[23953] <=  8'h78;        memory[23954] <=  8'h62;        memory[23955] <=  8'h61;        memory[23956] <=  8'h72;        memory[23957] <=  8'h74;        memory[23958] <=  8'h78;        memory[23959] <=  8'h61;        memory[23960] <=  8'h74;        memory[23961] <=  8'h6b;        memory[23962] <=  8'h73;        memory[23963] <=  8'h68;        memory[23964] <=  8'h63;        memory[23965] <=  8'h66;        memory[23966] <=  8'h69;        memory[23967] <=  8'h77;        memory[23968] <=  8'h68;        memory[23969] <=  8'h61;        memory[23970] <=  8'h74;        memory[23971] <=  8'h61;        memory[23972] <=  8'h6e;        memory[23973] <=  8'h61;        memory[23974] <=  8'h62;        memory[23975] <=  8'h61;        memory[23976] <=  8'h63;        memory[23977] <=  8'h61;        memory[23978] <=  8'h74;        memory[23979] <=  8'h61;        memory[23980] <=  8'h62;        memory[23981] <=  8'h61;        memory[23982] <=  8'h72;        memory[23983] <=  8'h63;        memory[23984] <=  8'h61;        memory[23985] <=  8'h68;        memory[23986] <=  8'h64;        memory[23987] <=  8'h75;        memory[23988] <=  8'h63;        memory[23989] <=  8'h74;        memory[23990] <=  8'h61;        memory[23991] <=  8'h64;        memory[23992] <=  8'h61;        memory[23993] <=  8'h61;        memory[23994] <=  8'h63;        memory[23995] <=  8'h61;        memory[23996] <=  8'h72;        memory[23997] <=  8'h62;        memory[23998] <=  8'h61;        memory[23999] <=  8'h72;        memory[24000] <=  8'h74;        memory[24001] <=  8'h78;        memory[24002] <=  8'h61;        memory[24003] <=  8'h74;        memory[24004] <=  8'h6b;        memory[24005] <=  8'h73;        memory[24006] <=  8'h68;        memory[24007] <=  8'h63;        memory[24008] <=  8'h66;        memory[24009] <=  8'h69;        memory[24010] <=  8'h77;        memory[24011] <=  8'h68;        memory[24012] <=  8'h61;        memory[24013] <=  8'h74;        memory[24014] <=  8'h61;        memory[24015] <=  8'h6e;        memory[24016] <=  8'h61;        memory[24017] <=  8'h62;        memory[24018] <=  8'h61;        memory[24019] <=  8'h63;        memory[24020] <=  8'h61;        memory[24021] <=  8'h74;        memory[24022] <=  8'h61;        memory[24023] <=  8'h62;        memory[24024] <=  8'h61;        memory[24025] <=  8'h72;        memory[24026] <=  8'h63;        memory[24027] <=  8'h61;        memory[24028] <=  8'h68;        memory[24029] <=  8'h64;        memory[24030] <=  8'h75;        memory[24031] <=  8'h63;        memory[24032] <=  8'h74;        memory[24033] <=  8'h61;        memory[24034] <=  8'h64;        memory[24035] <=  8'h61;        memory[24036] <=  8'h61;        memory[24037] <=  8'h63;        memory[24038] <=  8'h61;        memory[24039] <=  8'h72;        memory[24040] <=  8'h62;        memory[24041] <=  8'h61;        memory[24042] <=  8'h72;        memory[24043] <=  8'h74;        memory[24044] <=  8'h78;        memory[24045] <=  8'h61;        memory[24046] <=  8'h74;        memory[24047] <=  8'h6b;        memory[24048] <=  8'h73;        memory[24049] <=  8'h68;        memory[24050] <=  8'h63;        memory[24051] <=  8'h66;        memory[24052] <=  8'h69;        memory[24053] <=  8'h77;        memory[24054] <=  8'h68;        memory[24055] <=  8'h61;        memory[24056] <=  8'h74;        memory[24057] <=  8'h61;        memory[24058] <=  8'h6e;        memory[24059] <=  8'h61;        memory[24060] <=  8'h62;        memory[24061] <=  8'h61;        memory[24062] <=  8'h63;        memory[24063] <=  8'h61;        memory[24064] <=  8'h74;        memory[24065] <=  8'h61;        memory[24066] <=  8'h62;        memory[24067] <=  8'h61;        memory[24068] <=  8'h72;        memory[24069] <=  8'h63;        memory[24070] <=  8'h61;        memory[24071] <=  8'h68;        memory[24072] <=  8'h64;        memory[24073] <=  8'h75;        memory[24074] <=  8'h63;        memory[24075] <=  8'h74;        memory[24076] <=  8'h61;        memory[24077] <=  8'h64;        memory[24078] <=  8'h61;        memory[24079] <=  8'h61;        memory[24080] <=  8'h63;        memory[24081] <=  8'h61;        memory[24082] <=  8'h72;        memory[24083] <=  8'h62;        memory[24084] <=  8'h61;        memory[24085] <=  8'h72;        memory[24086] <=  8'h74;        memory[24087] <=  8'h78;        memory[24088] <=  8'h61;        memory[24089] <=  8'h74;        memory[24090] <=  8'h6b;        memory[24091] <=  8'h73;        memory[24092] <=  8'h68;        memory[24093] <=  8'h63;        memory[24094] <=  8'h66;        memory[24095] <=  8'h69;        memory[24096] <=  8'h77;        memory[24097] <=  8'h68;        memory[24098] <=  8'h61;        memory[24099] <=  8'h74;        memory[24100] <=  8'h61;        memory[24101] <=  8'h6e;        memory[24102] <=  8'h61;        memory[24103] <=  8'h62;        memory[24104] <=  8'h61;        memory[24105] <=  8'h63;        memory[24106] <=  8'h61;        memory[24107] <=  8'h74;        memory[24108] <=  8'h61;        memory[24109] <=  8'h62;        memory[24110] <=  8'h61;        memory[24111] <=  8'h72;        memory[24112] <=  8'h63;        memory[24113] <=  8'h61;        memory[24114] <=  8'h68;        memory[24115] <=  8'h64;        memory[24116] <=  8'h75;        memory[24117] <=  8'h63;        memory[24118] <=  8'h74;        memory[24119] <=  8'h61;        memory[24120] <=  8'h64;        memory[24121] <=  8'h61;        memory[24122] <=  8'h61;        memory[24123] <=  8'h63;        memory[24124] <=  8'h61;        memory[24125] <=  8'h72;        memory[24126] <=  8'h62;        memory[24127] <=  8'h61;        memory[24128] <=  8'h72;        memory[24129] <=  8'h74;        memory[24130] <=  8'h78;        memory[24131] <=  8'h61;        memory[24132] <=  8'h74;        memory[24133] <=  8'h6b;        memory[24134] <=  8'h73;        memory[24135] <=  8'h68;        memory[24136] <=  8'h63;        memory[24137] <=  8'h66;        memory[24138] <=  8'h69;        memory[24139] <=  8'h77;        memory[24140] <=  8'h68;        memory[24141] <=  8'h61;        memory[24142] <=  8'h74;        memory[24143] <=  8'h61;        memory[24144] <=  8'h6e;        memory[24145] <=  8'h61;        memory[24146] <=  8'h62;        memory[24147] <=  8'h61;        memory[24148] <=  8'h63;        memory[24149] <=  8'h61;        memory[24150] <=  8'h74;        memory[24151] <=  8'h61;        memory[24152] <=  8'h62;        memory[24153] <=  8'h61;        memory[24154] <=  8'h72;        memory[24155] <=  8'h63;        memory[24156] <=  8'h61;        memory[24157] <=  8'h68;        memory[24158] <=  8'h64;        memory[24159] <=  8'h75;        memory[24160] <=  8'h63;        memory[24161] <=  8'h74;        memory[24162] <=  8'h61;        memory[24163] <=  8'h64;        memory[24164] <=  8'h61;        memory[24165] <=  8'h61;        memory[24166] <=  8'h63;        memory[24167] <=  8'h61;        memory[24168] <=  8'h72;        memory[24169] <=  8'h62;        memory[24170] <=  8'h61;        memory[24171] <=  8'h72;        memory[24172] <=  8'h74;        memory[24173] <=  8'h78;        memory[24174] <=  8'h61;        memory[24175] <=  8'h74;        memory[24176] <=  8'h6b;        memory[24177] <=  8'h73;        memory[24178] <=  8'h68;        memory[24179] <=  8'h63;        memory[24180] <=  8'h66;        memory[24181] <=  8'h69;        memory[24182] <=  8'h77;        memory[24183] <=  8'h68;        memory[24184] <=  8'h61;        memory[24185] <=  8'h74;        memory[24186] <=  8'h61;        memory[24187] <=  8'h6e;        memory[24188] <=  8'h61;        memory[24189] <=  8'h62;        memory[24190] <=  8'h61;        memory[24191] <=  8'h63;        memory[24192] <=  8'h61;        memory[24193] <=  8'h74;        memory[24194] <=  8'h61;        memory[24195] <=  8'h62;        memory[24196] <=  8'h61;        memory[24197] <=  8'h72;        memory[24198] <=  8'h63;        memory[24199] <=  8'h61;        memory[24200] <=  8'h68;        memory[24201] <=  8'h64;        memory[24202] <=  8'h75;        memory[24203] <=  8'h63;        memory[24204] <=  8'h74;        memory[24205] <=  8'h61;        memory[24206] <=  8'h64;        memory[24207] <=  8'h61;        memory[24208] <=  8'h61;        memory[24209] <=  8'h63;        memory[24210] <=  8'h61;        memory[24211] <=  8'h72;        memory[24212] <=  8'h62;        memory[24213] <=  8'h61;        memory[24214] <=  8'h72;        memory[24215] <=  8'h74;        memory[24216] <=  8'h78;        memory[24217] <=  8'h61;        memory[24218] <=  8'h74;        memory[24219] <=  8'h6b;        memory[24220] <=  8'h73;        memory[24221] <=  8'h68;        memory[24222] <=  8'h63;        memory[24223] <=  8'h66;        memory[24224] <=  8'h69;        memory[24225] <=  8'h77;        memory[24226] <=  8'h68;        memory[24227] <=  8'h61;        memory[24228] <=  8'h74;        memory[24229] <=  8'h61;        memory[24230] <=  8'h6e;        memory[24231] <=  8'h61;        memory[24232] <=  8'h62;        memory[24233] <=  8'h61;        memory[24234] <=  8'h63;        memory[24235] <=  8'h61;        memory[24236] <=  8'h74;        memory[24237] <=  8'h61;        memory[24238] <=  8'h62;        memory[24239] <=  8'h61;        memory[24240] <=  8'h72;        memory[24241] <=  8'h63;        memory[24242] <=  8'h61;        memory[24243] <=  8'h68;        memory[24244] <=  8'h64;        memory[24245] <=  8'h75;        memory[24246] <=  8'h63;        memory[24247] <=  8'h74;        memory[24248] <=  8'h61;        memory[24249] <=  8'h64;        memory[24250] <=  8'h61;        memory[24251] <=  8'h61;        memory[24252] <=  8'h63;        memory[24253] <=  8'h61;        memory[24254] <=  8'h72;        memory[24255] <=  8'h62;        memory[24256] <=  8'h61;        memory[24257] <=  8'h72;        memory[24258] <=  8'h74;        memory[24259] <=  8'h78;        memory[24260] <=  8'h61;        memory[24261] <=  8'h74;        memory[24262] <=  8'h6b;        memory[24263] <=  8'h73;        memory[24264] <=  8'h68;        memory[24265] <=  8'h63;        memory[24266] <=  8'h66;        memory[24267] <=  8'h69;        memory[24268] <=  8'h77;        memory[24269] <=  8'h68;        memory[24270] <=  8'h61;        memory[24271] <=  8'h74;        memory[24272] <=  8'h61;        memory[24273] <=  8'h6e;        memory[24274] <=  8'h61;        memory[24275] <=  8'h62;        memory[24276] <=  8'h61;        memory[24277] <=  8'h63;        memory[24278] <=  8'h61;        memory[24279] <=  8'h74;        memory[24280] <=  8'h61;        memory[24281] <=  8'h62;        memory[24282] <=  8'h61;        memory[24283] <=  8'h72;        memory[24284] <=  8'h63;        memory[24285] <=  8'h61;        memory[24286] <=  8'h68;        memory[24287] <=  8'h64;        memory[24288] <=  8'h75;        memory[24289] <=  8'h63;        memory[24290] <=  8'h74;        memory[24291] <=  8'h61;        memory[24292] <=  8'h64;        memory[24293] <=  8'h61;        memory[24294] <=  8'h61;        memory[24295] <=  8'h63;        memory[24296] <=  8'h61;        memory[24297] <=  8'h72;        memory[24298] <=  8'h62;        memory[24299] <=  8'h61;        memory[24300] <=  8'h72;        memory[24301] <=  8'h74;        memory[24302] <=  8'h78;        memory[24303] <=  8'h61;        memory[24304] <=  8'h74;        memory[24305] <=  8'h6b;        memory[24306] <=  8'h73;        memory[24307] <=  8'h68;        memory[24308] <=  8'h63;        memory[24309] <=  8'h66;        memory[24310] <=  8'h69;        memory[24311] <=  8'h77;        memory[24312] <=  8'h68;        memory[24313] <=  8'h61;        memory[24314] <=  8'h74;        memory[24315] <=  8'h61;        memory[24316] <=  8'h6e;        memory[24317] <=  8'h61;        memory[24318] <=  8'h62;        memory[24319] <=  8'h61;        memory[24320] <=  8'h63;        memory[24321] <=  8'h61;        memory[24322] <=  8'h74;        memory[24323] <=  8'h61;        memory[24324] <=  8'h62;        memory[24325] <=  8'h61;        memory[24326] <=  8'h72;        memory[24327] <=  8'h63;        memory[24328] <=  8'h61;        memory[24329] <=  8'h68;        memory[24330] <=  8'h64;        memory[24331] <=  8'h75;        memory[24332] <=  8'h63;        memory[24333] <=  8'h74;        memory[24334] <=  8'h61;        memory[24335] <=  8'h64;        memory[24336] <=  8'h61;        memory[24337] <=  8'h61;        memory[24338] <=  8'h63;        memory[24339] <=  8'h61;        memory[24340] <=  8'h72;        memory[24341] <=  8'h62;        memory[24342] <=  8'h61;        memory[24343] <=  8'h72;        memory[24344] <=  8'h74;        memory[24345] <=  8'h74;        memory[24346] <=  8'h62;        memory[24347] <=  8'h61;        memory[24348] <=  8'h72;        memory[24349] <=  8'h74;        memory[24350] <=  8'h78;        memory[24351] <=  8'h61;        memory[24352] <=  8'h74;        memory[24353] <=  8'h6b;        memory[24354] <=  8'h73;        memory[24355] <=  8'h68;        memory[24356] <=  8'h63;        memory[24357] <=  8'h66;        memory[24358] <=  8'h69;        memory[24359] <=  8'h77;        memory[24360] <=  8'h68;        memory[24361] <=  8'h61;        memory[24362] <=  8'h74;        memory[24363] <=  8'h61;        memory[24364] <=  8'h6e;        memory[24365] <=  8'h61;        memory[24366] <=  8'h62;        memory[24367] <=  8'h61;        memory[24368] <=  8'h63;        memory[24369] <=  8'h61;        memory[24370] <=  8'h74;        memory[24371] <=  8'h61;        memory[24372] <=  8'h62;        memory[24373] <=  8'h61;        memory[24374] <=  8'h72;        memory[24375] <=  8'h63;        memory[24376] <=  8'h61;        memory[24377] <=  8'h68;        memory[24378] <=  8'h64;        memory[24379] <=  8'h75;        memory[24380] <=  8'h63;        memory[24381] <=  8'h74;        memory[24382] <=  8'h61;        memory[24383] <=  8'h64;        memory[24384] <=  8'h61;        memory[24385] <=  8'h61;        memory[24386] <=  8'h63;        memory[24387] <=  8'h61;        memory[24388] <=  8'h72;        memory[24389] <=  8'h63;        memory[24390] <=  8'h74;        memory[24391] <=  8'h72;        memory[24392] <=  8'h63;        memory[24393] <=  8'h61;        memory[24394] <=  8'h74;        memory[24395] <=  8'h72;        memory[24396] <=  8'h63;        memory[24397] <=  8'h61;        memory[24398] <=  8'h74;        memory[24399] <=  8'h63;        memory[24400] <=  8'h62;        memory[24401] <=  8'h61;        memory[24402] <=  8'h74;        memory[24403] <=  8'h62;        memory[24404] <=  8'h72;        memory[24405] <=  8'h63;        memory[24406] <=  8'h61;        memory[24407] <=  8'h72;        memory[24408] <=  8'h62;        memory[24409] <=  8'h78;        memory[24410] <=  8'h74;        memory[24411] <=  8'h61;        memory[24412] <=  8'h72;        memory[24413] <=  8'h64;        memory[24414] <=  8'h66;        memory[24415] <=  8'h73;        memory[24416] <=  8'h67;        memory[24417] <=  8'h76;        memory[24418] <=  8'h68;        memory[24419] <=  8'h62;        memory[24420] <=  8'h6b;        memory[24421] <=  8'h6a;        memory[24422] <=  8'h6e;        memory[24423] <=  8'h6d;        memory[24424] <=  8'h62;        memory[24425] <=  8'h76;        memory[24426] <=  8'h78;        memory[24427] <=  8'h63;        memory[24428] <=  8'h73;        memory[24429] <=  8'h66;        memory[24430] <=  8'h72;        memory[24431] <=  8'h74;        memory[24432] <=  8'h79;        memory[24433] <=  8'h75;        memory[24434] <=  8'h6a;        memory[24435] <=  8'h6e;        memory[24436] <=  8'h62;        memory[24437] <=  8'h76;        memory[24438] <=  8'h63;        memory[24439] <=  8'h64;        memory[24440] <=  8'h74;        memory[24441] <=  8'h79;        memory[24442] <=  8'h75;        memory[24443] <=  8'h69;        memory[24444] <=  8'h6b;        memory[24445] <=  8'h6d;        memory[24446] <=  8'h6e;        memory[24447] <=  8'h62;        memory[24448] <=  8'h76;        memory[24449] <=  8'h63;        memory[24450] <=  8'h78;        memory[24451] <=  8'h73;        memory[24452] <=  8'h64;        memory[24453] <=  8'h72;        memory[24454] <=  8'h74;        memory[24455] <=  8'h79;        memory[24456] <=  8'h75;        memory[24457] <=  8'h69;        memory[24458] <=  8'h6b;        memory[24459] <=  8'h6d;        memory[24460] <=  8'h6e;        memory[24461] <=  8'h62;        memory[24462] <=  8'h76;        memory[24463] <=  8'h63;        memory[24464] <=  8'h73;        memory[24465] <=  8'h77;        memory[24466] <=  8'h33;        memory[24467] <=  8'h34;        memory[24468] <=  8'h35;        memory[24469] <=  8'h36;        memory[24470] <=  8'h37;        memory[24471] <=  8'h38;        memory[24472] <=  8'h69;        memory[24473] <=  8'h6b;        memory[24474] <=  8'h6d;        memory[24475] <=  8'h6e;        memory[24476] <=  8'h62;        memory[24477] <=  8'h76;        memory[24478] <=  8'h63;        memory[24479] <=  8'h64;        memory[24480] <=  8'h65;        memory[24481] <=  8'h72;        memory[24482] <=  8'h36;        memory[24483] <=  8'h37;        memory[24484] <=  8'h38;        memory[24485] <=  8'h69;        memory[24486] <=  8'h6f;        memory[24487] <=  8'h6b;        memory[24488] <=  8'h6a;        memory[24489] <=  8'h6e;        memory[24490] <=  8'h62;        memory[24491] <=  8'h76;        memory[24492] <=  8'h63;        memory[24493] <=  8'h64;        memory[24494] <=  8'h72;        memory[24495] <=  8'h74;        memory[24496] <=  8'h79;        memory[24497] <=  8'h75;        memory[24498] <=  8'h73;        memory[24499] <=  8'h6a;        memory[24500] <=  8'h63;        memory[24501] <=  8'h6e;        memory[24502] <=  8'h62;        memory[24503] <=  8'h64;        memory[24504] <=  8'h66;        memory[24505] <=  8'h73;        memory[24506] <=  8'h74;        memory[24507] <=  8'h79;        memory[24508] <=  8'h75;        memory[24509] <=  8'h61;        memory[24510] <=  8'h69;        memory[24511] <=  8'h6b;        memory[24512] <=  8'h78;        memory[24513] <=  8'h6d;        memory[24514] <=  8'h6e;        memory[24515] <=  8'h73;        memory[24516] <=  8'h6a;        memory[24517] <=  8'h6f;        memory[24518] <=  8'h64;        memory[24519] <=  8'h6c;        memory[24520] <=  8'h63;        memory[24521] <=  8'h78;        memory[24522] <=  8'h2c;        memory[24523] <=  8'h6d;        memory[24524] <=  8'h73;        memory[24525] <=  8'h6b;        memory[24526] <=  8'h64;        memory[24527] <=  8'h6c;        memory[24528] <=  8'h70;        memory[24529] <=  8'h5b;        memory[24530] <=  8'h3b;        memory[24531] <=  8'h73;        memory[24532] <=  8'h6c;        memory[24533] <=  8'h64;        memory[24534] <=  8'h70;        memory[24535] <=  8'h76;        memory[24536] <=  8'h63;        memory[24537] <=  8'h5b;        memory[24538] <=  8'h78;        memory[24539] <=  8'h76;        memory[24540] <=  8'h63;        memory[24541] <=  8'h5b;        memory[24542] <=  8'h78;        memory[24543] <=  8'h70;        memory[24544] <=  8'h6f;        memory[24545] <=  8'h20;        memory[24546] <=  8'h62;        memory[24547] <=  8'h61;        memory[24548] <=  8'h72;        memory[24549] <=  8'h74;        memory[24550] <=  8'h74;        memory[24551] <=  8'h62;        memory[24552] <=  8'h61;        memory[24553] <=  8'h72;        memory[24554] <=  8'h74;        memory[24555] <=  8'h78;        memory[24556] <=  8'h61;        memory[24557] <=  8'h74;        memory[24558] <=  8'h6b;        memory[24559] <=  8'h73;        memory[24560] <=  8'h68;        memory[24561] <=  8'h63;        memory[24562] <=  8'h66;        memory[24563] <=  8'h69;        memory[24564] <=  8'h77;        memory[24565] <=  8'h68;        memory[24566] <=  8'h61;        memory[24567] <=  8'h69;        memory[24568] <=  8'h6a;        memory[24569] <=  8'h78;        memory[24570] <=  8'h5d;        memory[24571] <=  8'h65;        memory[24572] <=  8'h6b;        memory[24573] <=  8'h6f;        memory[24574] <=  8'h39;        memory[24575] <=  8'h64;        memory[24576] <=  8'h75;        memory[24577] <=  8'h38;        memory[24578] <=  8'h79;        memory[24579] <=  8'h20;        memory[24580] <=  8'h37;        memory[24581] <=  8'h63;        memory[24582] <=  8'h67;        memory[24583] <=  8'h78;        memory[24584] <=  8'h63;        memory[24585] <=  8'h75;        memory[24586] <=  8'h68;        memory[24587] <=  8'h69;        memory[24588] <=  8'h6a;        memory[24589] <=  8'h77;        memory[24590] <=  8'h69;        memory[24591] <=  8'h64;        memory[24592] <=  8'h66;        memory[24593] <=  8'h68;        memory[24594] <=  8'h75;        memory[24595] <=  8'h76;        memory[24596] <=  8'h64;        memory[24597] <=  8'h62;        memory[24598] <=  8'h66;        memory[24599] <=  8'h6a;        memory[24600] <=  8'h6e;        memory[24601] <=  8'h6b;        memory[24602] <=  8'h6a;        memory[24603] <=  8'h65;        memory[24604] <=  8'h38;        memory[24605] <=  8'h66;        memory[24606] <=  8'h37;        memory[24607] <=  8'h67;        memory[24608] <=  8'h79;        memory[24609] <=  8'h76;        memory[24610] <=  8'h63;        memory[24611] <=  8'h68;        memory[24612] <=  8'h69;        memory[24613] <=  8'h6a;        memory[24614] <=  8'h33;        memory[24615] <=  8'h65;        memory[24616] <=  8'h67;        memory[24617] <=  8'h79;        memory[24618] <=  8'h72;        memory[24619] <=  8'h64;        memory[24620] <=  8'h62;        memory[24621] <=  8'h6e;        memory[24622] <=  8'h63;        memory[24623] <=  8'h7a;        memory[24624] <=  8'h6a;        memory[24625] <=  8'h6f;        memory[24626] <=  8'h66;        memory[24627] <=  8'h78;        memory[24628] <=  8'h6a;        memory[24629] <=  8'h69;        memory[24630] <=  8'h63;        memory[24631] <=  8'h68;        memory[24632] <=  8'h62;        memory[24633] <=  8'h6e;        memory[24634] <=  8'h6d;        memory[24635] <=  8'h63;        memory[24636] <=  8'h73;        memory[24637] <=  8'h6c;        memory[24638] <=  8'h6b;        memory[24639] <=  8'h6a;        memory[24640] <=  8'h69;        memory[24641] <=  8'h68;        memory[24642] <=  8'h76;        memory[24643] <=  8'h75;        memory[24644] <=  8'h69;        memory[24645] <=  8'h64;        memory[24646] <=  8'h68;        memory[24647] <=  8'h75;        memory[24648] <=  8'h67;        memory[24649] <=  8'h79;        memory[24650] <=  8'h62;        memory[24651] <=  8'h68;        memory[24652] <=  8'h65;        memory[24653] <=  8'h6a;        memory[24654] <=  8'h72;        memory[24655] <=  8'h6b;        memory[24656] <=  8'h6a;        memory[24657] <=  8'h6f;        memory[24658] <=  8'h64;        memory[24659] <=  8'h67;        memory[24660] <=  8'h69;        memory[24661] <=  8'h75;        memory[24662] <=  8'h69;        memory[24663] <=  8'h67;        memory[24664] <=  8'h76;        memory[24665] <=  8'h79;        memory[24666] <=  8'h75;        memory[24667] <=  8'h67;        memory[24668] <=  8'h78;        memory[24669] <=  8'h68;        memory[24670] <=  8'h63;        memory[24671] <=  8'h20;        memory[24672] <=  8'h20;        memory[24673] <=  8'h20;        memory[24674] <=  8'h78;        memory[24675] <=  8'h76;        memory[24676] <=  8'h20;        memory[24677] <=  8'h63;        memory[24678] <=  8'h78;        memory[24679] <=  8'h67;        memory[24680] <=  8'h79;        memory[24681] <=  8'h63;        memory[24682] <=  8'h75;        memory[24683] <=  8'h68;        memory[24684] <=  8'h6a;        memory[24685] <=  8'h6b;        memory[24686] <=  8'h61;        memory[24687] <=  8'h6c;        memory[24688] <=  8'h78;        memory[24689] <=  8'h76;        memory[24690] <=  8'h70;        memory[24691] <=  8'h6f;        memory[24692] <=  8'h69;        memory[24693] <=  8'h6a;        memory[24694] <=  8'h69;        memory[24695] <=  8'h68;        memory[24696] <=  8'h6a;        memory[24697] <=  8'h62;        memory[24698] <=  8'h77;        memory[24699] <=  8'h65;        memory[24700] <=  8'h6e;        memory[24701] <=  8'h61;        memory[24702] <=  8'h66;        memory[24703] <=  8'h6d;        memory[24704] <=  8'h64;        memory[24705] <=  8'h6b;        memory[24706] <=  8'h6d;        memory[24707] <=  8'h76;        memory[24708] <=  8'h6c;        memory[24709] <=  8'h63;        memory[24710] <=  8'h6f;        memory[24711] <=  8'h64;        memory[24712] <=  8'h69;        memory[24713] <=  8'h75;        memory[24714] <=  8'h68;        memory[24715] <=  8'h73;        memory[24716] <=  8'h66;        memory[24717] <=  8'h65;        memory[24718] <=  8'h62;        memory[24719] <=  8'h6e;        memory[24720] <=  8'h64;        memory[24721] <=  8'h73;        memory[24722] <=  8'h63;        memory[24723] <=  8'h6b;        memory[24724] <=  8'h20;        memory[24725] <=  8'h78;        memory[24726] <=  8'h6a;        memory[24727] <=  8'h78;        memory[24728] <=  8'h63;        memory[24729] <=  8'h73;        memory[24730] <=  8'h64;        memory[24731] <=  8'h66;        memory[24732] <=  8'h6b;        memory[24733] <=  8'h64;        memory[24734] <=  8'h6e;        memory[24735] <=  8'h6d;        memory[24736] <=  8'h64;        memory[24737] <=  8'h73;        memory[24738] <=  8'h63;        memory[24739] <=  8'h6b;        memory[24740] <=  8'h78;        memory[24741] <=  8'h6c;        memory[24742] <=  8'h6f;        memory[24743] <=  8'h66;        memory[24744] <=  8'h6a;        memory[24745] <=  8'h69;        memory[24746] <=  8'h61;        memory[24747] <=  8'h62;        memory[24748] <=  8'h6e;        memory[24749] <=  8'h20;        memory[24750] <=  8'h78;        memory[24751] <=  8'h6b;        memory[24752] <=  8'h6d;        memory[24753] <=  8'h20;        memory[24754] <=  8'h6f;        memory[24755] <=  8'h63;        memory[24756] <=  8'h76;        memory[24757] <=  8'h73;        memory[24758] <=  8'h64;        memory[24759] <=  8'h69;        memory[24760] <=  8'h66;        memory[24761] <=  8'h68;        memory[24762] <=  8'h65;        memory[24763] <=  8'h71;        memory[24764] <=  8'h6a;        memory[24765] <=  8'h77;        memory[24766] <=  8'h62;        memory[24767] <=  8'h65;        memory[24768] <=  8'h6e;        memory[24769] <=  8'h20;        memory[24770] <=  8'h6d;        memory[24771] <=  8'h64;        memory[24772] <=  8'h73;        memory[24773] <=  8'h6c;        memory[24774] <=  8'h76;        memory[24775] <=  8'h6b;        memory[24776] <=  8'h63;        memory[24777] <=  8'h78;        memory[24778] <=  8'h20;        memory[24779] <=  8'h6f;        memory[24780] <=  8'h78;        memory[24781] <=  8'h69;        memory[24782] <=  8'h63;        memory[24783] <=  8'h6a;        memory[24784] <=  8'h76;        memory[24785] <=  8'h64;        memory[24786] <=  8'h66;        memory[24787] <=  8'h65;        memory[24788] <=  8'h71;        memory[24789] <=  8'h6e;        memory[24790] <=  8'h20;        memory[24791] <=  8'h64;        memory[24792] <=  8'h6d;        memory[24793] <=  8'h73;        memory[24794] <=  8'h6c;        memory[24795] <=  8'h63;        memory[24796] <=  8'h78;        memory[24797] <=  8'h6b;        memory[24798] <=  8'h20;        memory[24799] <=  8'h6f;        memory[24800] <=  8'h78;        memory[24801] <=  8'h63;        memory[24802] <=  8'h76;        memory[24803] <=  8'h6a;        memory[24804] <=  8'h64;        memory[24805] <=  8'h62;        memory[24806] <=  8'h71;        memory[24807] <=  8'h77;        memory[24808] <=  8'h65;        memory[24809] <=  8'h6e;        memory[24810] <=  8'h6d;        memory[24811] <=  8'h64;        memory[24812] <=  8'h6c;        memory[24813] <=  8'h73;        memory[24814] <=  8'h2c;        memory[24815] <=  8'h76;        memory[24816] <=  8'h63;        memory[24817] <=  8'h78;        memory[24818] <=  8'h20;        memory[24819] <=  8'h63;        memory[24820] <=  8'h6f;        memory[24821] <=  8'h69;        memory[24822] <=  8'h76;        memory[24823] <=  8'h68;        memory[24824] <=  8'h73;        memory[24825] <=  8'h64;        memory[24826] <=  8'h62;        memory[24827] <=  8'h71;        memory[24828] <=  8'h77;        memory[24829] <=  8'h65;        memory[24830] <=  8'h6e;        memory[24831] <=  8'h64;        memory[24832] <=  8'h6b;        memory[24833] <=  8'h73;        memory[24834] <=  8'h76;        memory[24835] <=  8'h6f;        memory[24836] <=  8'h63;        memory[24837] <=  8'h20;        memory[24838] <=  8'h76;        memory[24839] <=  8'h69;        memory[24840] <=  8'h75;        memory[24841] <=  8'h69;        memory[24842] <=  8'h68;        memory[24843] <=  8'h63;        memory[24844] <=  8'h78;        memory[24845] <=  8'h69;        memory[24846] <=  8'h6f;        memory[24847] <=  8'h76;        memory[24848] <=  8'h73;        memory[24849] <=  8'h64;        memory[24850] <=  8'h61;        memory[24851] <=  8'h64;        memory[24852] <=  8'h6e;        memory[24853] <=  8'h77;        memory[24854] <=  8'h71;        memory[24855] <=  8'h6b;        memory[24856] <=  8'h6c;        memory[24857] <=  8'h73;        memory[24858] <=  8'h76;        memory[24859] <=  8'h6e;        memory[24860] <=  8'h62;        memory[24861] <=  8'h20;        memory[24862] <=  8'h64;        memory[24863] <=  8'h66;        memory[24864] <=  8'h6a;        memory[24865] <=  8'h6b;        memory[24866] <=  8'h71;        memory[24867] <=  8'h64;        memory[24868] <=  8'h77;        memory[24869] <=  8'h65;        memory[24870] <=  8'h6e;        memory[24871] <=  8'h62;        memory[24872] <=  8'h20;        memory[24873] <=  8'h64;        memory[24874] <=  8'h73;        memory[24875] <=  8'h76;        memory[24876] <=  8'h68;        memory[24877] <=  8'h64;        memory[24878] <=  8'h61;        memory[24879] <=  8'h71;        memory[24880] <=  8'h77;        memory[24881] <=  8'h6a;        memory[24882] <=  8'h65;        memory[24883] <=  8'h6e;        memory[24884] <=  8'h64;        memory[24885] <=  8'h20;        memory[24886] <=  8'h61;        memory[24887] <=  8'h63;        memory[24888] <=  8'h62;        memory[24889] <=  8'h68;        memory[24890] <=  8'h64;        memory[24891] <=  8'h61;        memory[24892] <=  8'h77;        memory[24893] <=  8'h71;        memory[24894] <=  8'h6e;        memory[24895] <=  8'h20;        memory[24896] <=  8'h62;        memory[24897] <=  8'h73;        memory[24898] <=  8'h76;        memory[24899] <=  8'h61;        memory[24900] <=  8'h67;        memory[24901] <=  8'h76;        memory[24902] <=  8'h68;        memory[24903] <=  8'h67;        memory[24904] <=  8'h61;        memory[24905] <=  8'h73;        memory[24906] <=  8'h6a;        memory[24907] <=  8'h6b;        memory[24908] <=  8'h63;        memory[24909] <=  8'h78;        memory[24910] <=  8'h76;        memory[24911] <=  8'h6e;        memory[24912] <=  8'h73;        memory[24913] <=  8'h64;        memory[24914] <=  8'h20;        memory[24915] <=  8'h66;        memory[24916] <=  8'h62;        memory[24917] <=  8'h64;        memory[24918] <=  8'h61;        memory[24919] <=  8'h73;        memory[24920] <=  8'h76;        memory[24921] <=  8'h67;        memory[24922] <=  8'h63;        memory[24923] <=  8'h79;        memory[24924] <=  8'h7a;        memory[24925] <=  8'h78;        memory[24926] <=  8'h79;        memory[24927] <=  8'h75;        memory[24928] <=  8'h20;        memory[24929] <=  8'h69;        memory[24930] <=  8'h6a;        memory[24931] <=  8'h64;        memory[24932] <=  8'h66;        memory[24933] <=  8'h6b;        memory[24934] <=  8'h61;        memory[24935] <=  8'h64;        memory[24936] <=  8'h63;        memory[24937] <=  8'h78;        memory[24938] <=  8'h68;        memory[24939] <=  8'h20;        memory[24940] <=  8'h67;        memory[24941] <=  8'h61;        memory[24942] <=  8'h68;        memory[24943] <=  8'h75;        memory[24944] <=  8'h64;        memory[24945] <=  8'h73;        memory[24946] <=  8'h69;        memory[24947] <=  8'h6a;        memory[24948] <=  8'h61;        memory[24949] <=  8'h6b;        memory[24950] <=  8'h63;        memory[24951] <=  8'h62;        memory[24952] <=  8'h61;        memory[24953] <=  8'h72;        memory[24954] <=  8'h73;        memory[24955] <=  8'h68;        memory[24956] <=  8'h64;        memory[24957] <=  8'h66;        memory[24958] <=  8'h67;        memory[24959] <=  8'h73;        memory[24960] <=  8'h68;        memory[24961] <=  8'h64;        memory[24962] <=  8'h66;        memory[24963] <=  8'h68;        memory[24964] <=  8'h64;        memory[24965] <=  8'h6a;        memory[24966] <=  8'h68;        memory[24967] <=  8'h62;        memory[24968] <=  8'h67;        memory[24969] <=  8'h63;        memory[24970] <=  8'h61;        memory[24971] <=  8'h66;        memory[24972] <=  8'h73;        memory[24973] <=  8'h79;        memory[24974] <=  8'h67;        memory[24975] <=  8'h6b;        memory[24976] <=  8'h75;        memory[24977] <=  8'h64;        memory[24978] <=  8'h68;        memory[24979] <=  8'h62;        memory[24980] <=  8'h77;        memory[24981] <=  8'h76;        memory[24982] <=  8'h67;        memory[24983] <=  8'h61;        memory[24984] <=  8'h66;        memory[24985] <=  8'h64;        memory[24986] <=  8'h74;        memory[24987] <=  8'h75;        memory[24988] <=  8'h66;        memory[24989] <=  8'h79;        memory[24990] <=  8'h67;        memory[24991] <=  8'h69;        memory[24992] <=  8'h75;        memory[24993] <=  8'h68;        memory[24994] <=  8'h6c;        memory[24995] <=  8'h6a;        memory[24996] <=  8'h62;        memory[24997] <=  8'h6b;        memory[24998] <=  8'h68;        memory[24999] <=  8'h76;        memory[25000] <=  8'h67;        memory[25001] <=  8'h63;        memory[25002] <=  8'h66;        memory[25003] <=  8'h78;        memory[25004] <=  8'h64;        memory[25005] <=  8'h74;        memory[25006] <=  8'h75;        memory[25007] <=  8'h79;        memory[25008] <=  8'h69;        memory[25009] <=  8'h75;        memory[25010] <=  8'h68;        memory[25011] <=  8'h6c;        memory[25012] <=  8'h6a;        memory[25013] <=  8'h6b;        memory[25014] <=  8'h67;        memory[25015] <=  8'h6a;        memory[25016] <=  8'h63;        memory[25017] <=  8'h66;        memory[25018] <=  8'h68;        memory[25019] <=  8'h64;        memory[25020] <=  8'h67;        memory[25021] <=  8'h72;        memory[25022] <=  8'h79;        memory[25023] <=  8'h74;        memory[25024] <=  8'h66;        memory[25025] <=  8'h75;        memory[25026] <=  8'h79;        memory[25027] <=  8'h69;        memory[25028] <=  8'h68;        memory[25029] <=  8'h6c;        memory[25030] <=  8'h62;        memory[25031] <=  8'h6d;        memory[25032] <=  8'h76;        memory[25033] <=  8'h6e;        memory[25034] <=  8'h63;        memory[25035] <=  8'h66;        memory[25036] <=  8'h68;        memory[25037] <=  8'h64;        memory[25038] <=  8'h74;        memory[25039] <=  8'h75;        memory[25040] <=  8'h67;        memory[25041] <=  8'h79;        memory[25042] <=  8'h69;        memory[25043] <=  8'h68;        memory[25044] <=  8'h75;        memory[25045] <=  8'h6a;        memory[25046] <=  8'h6c;        memory[25047] <=  8'h62;        memory[25048] <=  8'h6d;        memory[25049] <=  8'h76;        memory[25050] <=  8'h6e;        memory[25051] <=  8'h63;        memory[25052] <=  8'h66;        memory[25053] <=  8'h68;        memory[25054] <=  8'h67;        memory[25055] <=  8'h79;        memory[25056] <=  8'h68;        memory[25057] <=  8'h75;        memory[25058] <=  8'h6a;        memory[25059] <=  8'h6e;        memory[25060] <=  8'h2c;        memory[25061] <=  8'h62;        memory[25062] <=  8'h6e;        memory[25063] <=  8'h6d;        memory[25064] <=  8'h76;        memory[25065] <=  8'h6e;        memory[25066] <=  8'h63;        memory[25067] <=  8'h66;        memory[25068] <=  8'h68;        memory[25069] <=  8'h74;        memory[25070] <=  8'h79;        memory[25071] <=  8'h69;        memory[25072] <=  8'h75;        memory[25073] <=  8'h6c;        memory[25074] <=  8'h6a;        memory[25075] <=  8'h62;        memory[25076] <=  8'h6d;        memory[25077] <=  8'h76;        memory[25078] <=  8'h6e;        memory[25079] <=  8'h63;        memory[25080] <=  8'h66;        memory[25081] <=  8'h74;        memory[25082] <=  8'h75;        memory[25083] <=  8'h79;        memory[25084] <=  8'h69;        memory[25085] <=  8'h68;        memory[25086] <=  8'h6b;        memory[25087] <=  8'h62;        memory[25088] <=  8'h76;        memory[25089] <=  8'h63;        memory[25090] <=  8'h66;        memory[25091] <=  8'h67;        memory[25092] <=  8'h74;        memory[25093] <=  8'h75;        memory[25094] <=  8'h79;        memory[25095] <=  8'h69;        memory[25096] <=  8'h75;        memory[25097] <=  8'h68;        memory[25098] <=  8'h6a;        memory[25099] <=  8'h6b;        memory[25100] <=  8'h62;        memory[25101] <=  8'h76;        memory[25102] <=  8'h63;        memory[25103] <=  8'h66;        memory[25104] <=  8'h74;        memory[25105] <=  8'h75;        memory[25106] <=  8'h79;        memory[25107] <=  8'h69;        memory[25108] <=  8'h75;        memory[25109] <=  8'h6a;        memory[25110] <=  8'h6b;        memory[25111] <=  8'h6e;        memory[25112] <=  8'h62;        memory[25113] <=  8'h76;        memory[25114] <=  8'h67;        memory[25115] <=  8'h66;        memory[25116] <=  8'h74;        memory[25117] <=  8'h79;        memory[25118] <=  8'h75;        memory[25119] <=  8'h75;        memory[25120] <=  8'h69;        memory[25121] <=  8'h6a;        memory[25122] <=  8'h6b;        memory[25123] <=  8'h68;        memory[25124] <=  8'h62;        memory[25125] <=  8'h6a;        memory[25126] <=  8'h67;        memory[25127] <=  8'h68;        memory[25128] <=  8'h66;        memory[25129] <=  8'h79;        memory[25130] <=  8'h74;        memory[25131] <=  8'h79;        memory[25132] <=  8'h69;        memory[25133] <=  8'h75;        memory[25134] <=  8'h64;        memory[25135] <=  8'h6a;        memory[25136] <=  8'h6b;        memory[25137] <=  8'h68;        memory[25138] <=  8'h63;        memory[25139] <=  8'h7a;        memory[25140] <=  8'h67;        memory[25141] <=  8'h68;        memory[25142] <=  8'h74;        memory[25143] <=  8'h75;        memory[25144] <=  8'h79;        memory[25145] <=  8'h69;        memory[25146] <=  8'h61;        memory[25147] <=  8'h73;        memory[25148] <=  8'h75;        memory[25149] <=  8'h6a;        memory[25150] <=  8'h6b;        memory[25151] <=  8'h62;        memory[25152] <=  8'h6e;        memory[25153] <=  8'h61;        memory[25154] <=  8'h76;        memory[25155] <=  8'h63;        memory[25156] <=  8'h66;        memory[25157] <=  8'h68;        memory[25158] <=  8'h75;        memory[25159] <=  8'h61;        memory[25160] <=  8'h73;        memory[25161] <=  8'h79;        memory[25162] <=  8'h64;        memory[25163] <=  8'h75;        memory[25164] <=  8'h69;        memory[25165] <=  8'h6a;        memory[25166] <=  8'h61;        memory[25167] <=  8'h6b;        memory[25168] <=  8'h62;        memory[25169] <=  8'h63;        memory[25170] <=  8'h78;        memory[25171] <=  8'h68;        memory[25172] <=  8'h67;        memory[25173] <=  8'h79;        memory[25174] <=  8'h75;        memory[25175] <=  8'h7a;        memory[25176] <=  8'h63;        memory[25177] <=  8'h61;        memory[25178] <=  8'h73;        memory[25179] <=  8'h69;        memory[25180] <=  8'h75;        memory[25181] <=  8'h6f;        memory[25182] <=  8'h69;        memory[25183] <=  8'h6a;        memory[25184] <=  8'h61;        memory[25185] <=  8'h6c;        memory[25186] <=  8'h63;        memory[25187] <=  8'h78;        memory[25188] <=  8'h62;        memory[25189] <=  8'h63;        memory[25190] <=  8'h20;        memory[25191] <=  8'h6e;        memory[25192] <=  8'h76;        memory[25193] <=  8'h63;        memory[25194] <=  8'h61;        memory[25195] <=  8'h64;        memory[25196] <=  8'h73;        memory[25197] <=  8'h67;        memory[25198] <=  8'h79;        memory[25199] <=  8'h68;        memory[25200] <=  8'h75;        memory[25201] <=  8'h61;        memory[25202] <=  8'h6a;        memory[25203] <=  8'h6b;        memory[25204] <=  8'h78;        memory[25205] <=  8'h62;        memory[25206] <=  8'h20;        memory[25207] <=  8'h6e;        memory[25208] <=  8'h76;        memory[25209] <=  8'h63;        memory[25210] <=  8'h61;        memory[25211] <=  8'h73;        memory[25212] <=  8'h67;        memory[25213] <=  8'h68;        memory[25214] <=  8'h75;        memory[25215] <=  8'h6a;        memory[25216] <=  8'h6c;        memory[25217] <=  8'h6b;        memory[25218] <=  8'h63;        memory[25219] <=  8'h78;        memory[25220] <=  8'h20;        memory[25221] <=  8'h6a;        memory[25222] <=  8'h6b;        memory[25223] <=  8'h68;        memory[25224] <=  8'h61;        memory[25225] <=  8'h73;        memory[25226] <=  8'h76;        memory[25227] <=  8'h64;        memory[25228] <=  8'h6e;        memory[25229] <=  8'h20;        memory[25230] <=  8'h62;        memory[25231] <=  8'h6e;        memory[25232] <=  8'h6d;        memory[25233] <=  8'h6b;        memory[25234] <=  8'h77;        memory[25235] <=  8'h64;        memory[25236] <=  8'h6f;        memory[25237] <=  8'h77;        memory[25238] <=  8'h69;        memory[25239] <=  8'h6f;        memory[25240] <=  8'h75;        memory[25241] <=  8'h69;        memory[25242] <=  8'h68;        memory[25243] <=  8'h62;        memory[25244] <=  8'h6e;        memory[25245] <=  8'h6b;        memory[25246] <=  8'h77;        memory[25247] <=  8'h69;        memory[25248] <=  8'h6f;        memory[25249] <=  8'h75;        memory[25250] <=  8'h71;        memory[25251] <=  8'h69;        memory[25252] <=  8'h79;        memory[25253] <=  8'h67;        memory[25254] <=  8'h6a;        memory[25255] <=  8'h64;        memory[25256] <=  8'h61;        memory[25257] <=  8'h76;        memory[25258] <=  8'h62;        memory[25259] <=  8'h6e;        memory[25260] <=  8'h6b;        memory[25261] <=  8'h6f;        memory[25262] <=  8'h70;        memory[25263] <=  8'h64;        memory[25264] <=  8'h76;        memory[25265] <=  8'h69;        memory[25266] <=  8'h6f;        memory[25267] <=  8'h75;        memory[25268] <=  8'h69;        memory[25269] <=  8'h48;        memory[25270] <=  8'h42;        memory[25271] <=  8'h6b;        memory[25272] <=  8'h64;        memory[25273] <=  8'h6e;        memory[25274] <=  8'h6c;        memory[25275] <=  8'h71;        memory[25276] <=  8'h6b;        memory[25277] <=  8'h6d;        memory[25278] <=  8'h6a;        memory[25279] <=  8'h70;        memory[25280] <=  8'h69;        memory[25281] <=  8'h6f;        memory[25282] <=  8'h68;        memory[25283] <=  8'h65;        memory[25284] <=  8'h66;        memory[25285] <=  8'h75;        memory[25286] <=  8'h67;        memory[25287] <=  8'h69;        memory[25288] <=  8'h73;        memory[25289] <=  8'h61;        memory[25290] <=  8'h62;        memory[25291] <=  8'h64;        memory[25292] <=  8'h6b;        memory[25293] <=  8'h6a;        memory[25294] <=  8'h6b;        memory[25295] <=  8'h6c;        memory[25296] <=  8'h6a;        memory[25297] <=  8'h69;        memory[25298] <=  8'h73;        memory[25299] <=  8'h6f;        memory[25300] <=  8'h71;        memory[25301] <=  8'h68;        memory[25302] <=  8'h77;        memory[25303] <=  8'h67;        memory[25304] <=  8'h69;        memory[25305] <=  8'h79;        memory[25306] <=  8'h6a;        memory[25307] <=  8'h64;        memory[25308] <=  8'h76;        memory[25309] <=  8'h62;        memory[25310] <=  8'h6e;        memory[25311] <=  8'h61;        memory[25312] <=  8'h73;        memory[25313] <=  8'h66;        memory[25314] <=  8'h6c;        memory[25315] <=  8'h6b;        memory[25316] <=  8'h64;        memory[25317] <=  8'h6a;        memory[25318] <=  8'h68;        memory[25319] <=  8'h63;        memory[25320] <=  8'h67;        memory[25321] <=  8'h6a;        memory[25322] <=  8'h76;        memory[25323] <=  8'h73;        memory[25324] <=  8'h64;        memory[25325] <=  8'h62;        memory[25326] <=  8'h62;        memory[25327] <=  8'h61;        memory[25328] <=  8'h72;        memory[25329] <=  8'h62;        memory[25330] <=  8'h62;        memory[25331] <=  8'h73;        memory[25332] <=  8'h62;        memory[25333] <=  8'h67;        memory[25334] <=  8'h73;        memory[25335] <=  8'h66;        memory[25336] <=  8'h67;        memory[25337] <=  8'h61;        memory[25338] <=  8'h68;        memory[25339] <=  8'h66;        memory[25340] <=  8'h73;        memory[25341] <=  8'h68;        memory[25342] <=  8'h61;        memory[25343] <=  8'h66;        memory[25344] <=  8'h73;        memory[25345] <=  8'h66;        memory[25346] <=  8'h68;        memory[25347] <=  8'h61;        memory[25348] <=  8'h69;        memory[25349] <=  8'h64;        memory[25350] <=  8'h75;        memory[25351] <=  8'h67;        memory[25352] <=  8'h64;        memory[25353] <=  8'h77;        memory[25354] <=  8'h62;        memory[25355] <=  8'h61;        memory[25356] <=  8'h62;        memory[25357] <=  8'h72;        memory[25358] <=  8'h62;        memory[25359] <=  8'h61;        memory[25360] <=  8'h62;        memory[25361] <=  8'h62;        memory[25362] <=  8'h74;        memory[25363] <=  8'h62;        memory[25364] <=  8'h62;        memory[25365] <=  8'h62;        memory[25366] <=  8'h62;        memory[25367] <=  8'h62;        memory[25368] <=  8'h62;        memory[25369] <=  8'h62;        memory[25370] <=  8'h62;        memory[25371] <=  8'h61;        memory[25372] <=  8'h62;        memory[25373] <=  8'h62;        memory[25374] <=  8'h72;        memory[25375] <=  8'h74;        memory[25376] <=  8'h62;        memory[25377] <=  8'h62;        memory[25378] <=  8'h61;        memory[25379] <=  8'h62;        memory[25380] <=  8'h72;        memory[25381] <=  8'h62;        memory[25382] <=  8'h74;        memory[25383] <=  8'h62;        memory[25384] <=  8'h62;        memory[25385] <=  8'h62;        memory[25386] <=  8'h63;        memory[25387] <=  8'h61;        memory[25388] <=  8'h72;        memory[25389] <=  8'h74;        memory[25390] <=  8'h73;        memory[25391] <=  8'h62;        memory[25392] <=  8'h61;        memory[25393] <=  8'h72;        memory[25394] <=  8'h74;        memory[25395] <=  8'h74;        memory[25396] <=  8'h62;        memory[25397] <=  8'h61;        memory[25398] <=  8'h72;        memory[25399] <=  8'h74;        memory[25400] <=  8'h78;        memory[25401] <=  8'h61;        memory[25402] <=  8'h74;        memory[25403] <=  8'h6b;        memory[25404] <=  8'h73;        memory[25405] <=  8'h68;        memory[25406] <=  8'h63;        memory[25407] <=  8'h66;        memory[25408] <=  8'h69;        memory[25409] <=  8'h77;        memory[25410] <=  8'h68;        memory[25411] <=  8'h61;        memory[25412] <=  8'h74;        memory[25413] <=  8'h61;        memory[25414] <=  8'h6e;        memory[25415] <=  8'h61;        memory[25416] <=  8'h62;        memory[25417] <=  8'h61;        memory[25418] <=  8'h63;        memory[25419] <=  8'h61;        memory[25420] <=  8'h74;        memory[25421] <=  8'h61;        memory[25422] <=  8'h62;        memory[25423] <=  8'h61;        memory[25424] <=  8'h72;        memory[25425] <=  8'h63;        memory[25426] <=  8'h61;        memory[25427] <=  8'h68;        memory[25428] <=  8'h64;        memory[25429] <=  8'h75;        memory[25430] <=  8'h63;        memory[25431] <=  8'h74;        memory[25432] <=  8'h61;        memory[25433] <=  8'h64;        memory[25434] <=  8'h61;        memory[25435] <=  8'h61;        memory[25436] <=  8'h63;        memory[25437] <=  8'h61;        memory[25438] <=  8'h72;        memory[25439] <=  8'h63;        memory[25440] <=  8'h74;        memory[25441] <=  8'h72;        memory[25442] <=  8'h63;        memory[25443] <=  8'h61;        memory[25444] <=  8'h74;        memory[25445] <=  8'h72;        memory[25446] <=  8'h63;        memory[25447] <=  8'h61;        memory[25448] <=  8'h74;        memory[25449] <=  8'h63;        memory[25450] <=  8'h62;        memory[25451] <=  8'h61;        memory[25452] <=  8'h74;        memory[25453] <=  8'h62;        memory[25454] <=  8'h72;        memory[25455] <=  8'h63;        memory[25456] <=  8'h61;        memory[25457] <=  8'h74;        memory[25458] <=  8'h72;        memory[25459] <=  8'h6e;        memory[25460] <=  8'h62;        memory[25461] <=  8'h61;        memory[25462] <=  8'h63;        memory[25463] <=  8'h61;        memory[25464] <=  8'h74;        memory[25465] <=  8'h79;        memory[25466] <=  8'h73;        memory[25467] <=  8'h6e;        memory[25468] <=  8'h63;        memory[25469] <=  8'h74;        memory[25470] <=  8'h61;        memory[25471] <=  8'h6e;        memory[25472] <=  8'h62;        memory[25473] <=  8'h61;        memory[25474] <=  8'h63;        memory[25475] <=  8'h72;        memory[25476] <=  8'h6e;        memory[25477] <=  8'h74;        memory[25478] <=  8'h61;        memory[25479] <=  8'h62;        memory[25480] <=  8'h74;        memory[25481] <=  8'h6e;        memory[25482] <=  8'h61;        memory[25483] <=  8'h72;        memory[25484] <=  8'h62;        memory[25485] <=  8'h78;        memory[25486] <=  8'h74;        memory[25487] <=  8'h61;        memory[25488] <=  8'h72;        memory[25489] <=  8'h62;        memory[25490] <=  8'h61;        memory[25491] <=  8'h72;        memory[25492] <=  8'h74;        memory[25493] <=  8'h74;        memory[25494] <=  8'h62;        memory[25495] <=  8'h61;        memory[25496] <=  8'h72;        memory[25497] <=  8'h74;        memory[25498] <=  8'h78;        memory[25499] <=  8'h61;        memory[25500] <=  8'h74;        memory[25501] <=  8'h6b;        memory[25502] <=  8'h73;        memory[25503] <=  8'h68;        memory[25504] <=  8'h63;        memory[25505] <=  8'h66;        memory[25506] <=  8'h69;        memory[25507] <=  8'h77;        memory[25508] <=  8'h68;        memory[25509] <=  8'h61;        memory[25510] <=  8'h74;        memory[25511] <=  8'h61;        memory[25512] <=  8'h6e;        memory[25513] <=  8'h61;        memory[25514] <=  8'h62;        memory[25515] <=  8'h61;        memory[25516] <=  8'h63;        memory[25517] <=  8'h61;        memory[25518] <=  8'h74;        memory[25519] <=  8'h61;        memory[25520] <=  8'h62;        memory[25521] <=  8'h61;        memory[25522] <=  8'h72;        memory[25523] <=  8'h63;        memory[25524] <=  8'h61;        memory[25525] <=  8'h68;        memory[25526] <=  8'h64;        memory[25527] <=  8'h75;        memory[25528] <=  8'h63;        memory[25529] <=  8'h74;        memory[25530] <=  8'h61;        memory[25531] <=  8'h64;        memory[25532] <=  8'h61;        memory[25533] <=  8'h61;        memory[25534] <=  8'h63;        memory[25535] <=  8'h61;        memory[25536] <=  8'h72;        memory[25537] <=  8'h63;        memory[25538] <=  8'h74;        memory[25539] <=  8'h72;        memory[25540] <=  8'h63;        memory[25541] <=  8'h61;        memory[25542] <=  8'h74;        memory[25543] <=  8'h72;        memory[25544] <=  8'h63;        memory[25545] <=  8'h61;        memory[25546] <=  8'h74;        memory[25547] <=  8'h63;        memory[25548] <=  8'h62;        memory[25549] <=  8'h61;        memory[25550] <=  8'h74;        memory[25551] <=  8'h62;        memory[25552] <=  8'h72;        memory[25553] <=  8'h63;        memory[25554] <=  8'h61;        memory[25555] <=  8'h74;        memory[25556] <=  8'h72;        memory[25557] <=  8'h6e;        memory[25558] <=  8'h62;        memory[25559] <=  8'h61;        memory[25560] <=  8'h63;        memory[25561] <=  8'h61;        memory[25562] <=  8'h74;        memory[25563] <=  8'h79;        memory[25564] <=  8'h73;        memory[25565] <=  8'h6e;        memory[25566] <=  8'h63;        memory[25567] <=  8'h74;        memory[25568] <=  8'h61;        memory[25569] <=  8'h6e;        memory[25570] <=  8'h62;        memory[25571] <=  8'h61;        memory[25572] <=  8'h63;        memory[25573] <=  8'h72;        memory[25574] <=  8'h6e;        memory[25575] <=  8'h74;        memory[25576] <=  8'h61;        memory[25577] <=  8'h62;        memory[25578] <=  8'h74;        memory[25579] <=  8'h6e;        memory[25580] <=  8'h61;        memory[25581] <=  8'h72;        memory[25582] <=  8'h62;        memory[25583] <=  8'h78;        memory[25584] <=  8'h74;        memory[25585] <=  8'h61;        memory[25586] <=  8'h72;        memory[25587] <=  8'h62;        memory[25588] <=  8'h61;        memory[25589] <=  8'h72;        memory[25590] <=  8'h74;        memory[25591] <=  8'h74;        memory[25592] <=  8'h62;        memory[25593] <=  8'h61;        memory[25594] <=  8'h72;        memory[25595] <=  8'h74;        memory[25596] <=  8'h78;        memory[25597] <=  8'h61;        memory[25598] <=  8'h74;        memory[25599] <=  8'h6b;        memory[25600] <=  8'h73;        memory[25601] <=  8'h68;        memory[25602] <=  8'h63;        memory[25603] <=  8'h66;        memory[25604] <=  8'h69;        memory[25605] <=  8'h77;        memory[25606] <=  8'h68;        memory[25607] <=  8'h61;        memory[25608] <=  8'h74;        memory[25609] <=  8'h61;        memory[25610] <=  8'h6e;        memory[25611] <=  8'h61;        memory[25612] <=  8'h62;        memory[25613] <=  8'h61;        memory[25614] <=  8'h63;        memory[25615] <=  8'h61;        memory[25616] <=  8'h74;        memory[25617] <=  8'h61;        memory[25618] <=  8'h62;        memory[25619] <=  8'h61;        memory[25620] <=  8'h72;        memory[25621] <=  8'h63;        memory[25622] <=  8'h61;        memory[25623] <=  8'h68;        memory[25624] <=  8'h64;        memory[25625] <=  8'h75;        memory[25626] <=  8'h63;        memory[25627] <=  8'h74;        memory[25628] <=  8'h61;        memory[25629] <=  8'h64;        memory[25630] <=  8'h61;        memory[25631] <=  8'h61;        memory[25632] <=  8'h63;        memory[25633] <=  8'h61;        memory[25634] <=  8'h72;        memory[25635] <=  8'h63;        memory[25636] <=  8'h74;        memory[25637] <=  8'h72;        memory[25638] <=  8'h63;        memory[25639] <=  8'h61;        memory[25640] <=  8'h74;        memory[25641] <=  8'h72;        memory[25642] <=  8'h63;        memory[25643] <=  8'h61;        memory[25644] <=  8'h74;        memory[25645] <=  8'h63;        memory[25646] <=  8'h62;        memory[25647] <=  8'h61;        memory[25648] <=  8'h74;        memory[25649] <=  8'h62;        memory[25650] <=  8'h72;        memory[25651] <=  8'h63;        memory[25652] <=  8'h61;        memory[25653] <=  8'h74;        memory[25654] <=  8'h72;        memory[25655] <=  8'h6e;        memory[25656] <=  8'h62;        memory[25657] <=  8'h61;        memory[25658] <=  8'h63;        memory[25659] <=  8'h61;        memory[25660] <=  8'h74;        memory[25661] <=  8'h79;        memory[25662] <=  8'h73;        memory[25663] <=  8'h6e;        memory[25664] <=  8'h63;        memory[25665] <=  8'h74;        memory[25666] <=  8'h61;        memory[25667] <=  8'h6e;        memory[25668] <=  8'h62;        memory[25669] <=  8'h61;        memory[25670] <=  8'h63;        memory[25671] <=  8'h72;        memory[25672] <=  8'h6e;        memory[25673] <=  8'h74;        memory[25674] <=  8'h61;        memory[25675] <=  8'h62;        memory[25676] <=  8'h74;        memory[25677] <=  8'h6e;        memory[25678] <=  8'h61;        memory[25679] <=  8'h72;        memory[25680] <=  8'h62;        memory[25681] <=  8'h78;        memory[25682] <=  8'h74;        memory[25683] <=  8'h61;        memory[25684] <=  8'h72;        memory[25685] <=  8'h5d;        memory[25686] <=  8'h5d;        memory[25687] <=  8'h65;        memory[25688] <=  8'h66;        memory[25689] <=  8'h77;        memory[25690] <=  8'h65;        memory[25691] <=  8'h5d;        memory[25692] <=  8'h65;        memory[25693] <=  8'h67;        memory[25694] <=  8'h73;        memory[25695] <=  8'h67;        memory[25696] <=  8'h66;        memory[25697] <=  8'h62;        memory[25698] <=  8'h61;        memory[25699] <=  8'h72;        memory[25700] <=  8'h74;        memory[25701] <=  8'h74;        memory[25702] <=  8'h62;        memory[25703] <=  8'h61;        memory[25704] <=  8'h72;        memory[25705] <=  8'h74;        memory[25706] <=  8'h78;        memory[25707] <=  8'h61;        memory[25708] <=  8'h74;        memory[25709] <=  8'h6b;        memory[25710] <=  8'h73;        memory[25711] <=  8'h68;        memory[25712] <=  8'h63;        memory[25713] <=  8'h66;        memory[25714] <=  8'h69;        memory[25715] <=  8'h77;        memory[25716] <=  8'h68;        memory[25717] <=  8'h61;        memory[25718] <=  8'h74;        memory[25719] <=  8'h61;        memory[25720] <=  8'h6e;        memory[25721] <=  8'h61;        memory[25722] <=  8'h62;        memory[25723] <=  8'h61;        memory[25724] <=  8'h63;        memory[25725] <=  8'h61;        memory[25726] <=  8'h74;        memory[25727] <=  8'h61;        memory[25728] <=  8'h62;        memory[25729] <=  8'h61;        memory[25730] <=  8'h72;        memory[25731] <=  8'h63;        memory[25732] <=  8'h61;        memory[25733] <=  8'h68;        memory[25734] <=  8'h64;        memory[25735] <=  8'h75;        memory[25736] <=  8'h63;        memory[25737] <=  8'h74;        memory[25738] <=  8'h61;        memory[25739] <=  8'h64;        memory[25740] <=  8'h61;        memory[25741] <=  8'h61;        memory[25742] <=  8'h63;        memory[25743] <=  8'h61;        memory[25744] <=  8'h72;        memory[25745] <=  8'h63;        memory[25746] <=  8'h74;        memory[25747] <=  8'h72;        memory[25748] <=  8'h63;        memory[25749] <=  8'h61;        memory[25750] <=  8'h74;        memory[25751] <=  8'h72;        memory[25752] <=  8'h63;        memory[25753] <=  8'h61;        memory[25754] <=  8'h74;        memory[25755] <=  8'h63;        memory[25756] <=  8'h62;        memory[25757] <=  8'h61;        memory[25758] <=  8'h74;        memory[25759] <=  8'h62;        memory[25760] <=  8'h72;        memory[25761] <=  8'h63;        memory[25762] <=  8'h61;        memory[25763] <=  8'h74;        memory[25764] <=  8'h72;        memory[25765] <=  8'h6e;        memory[25766] <=  8'h62;        memory[25767] <=  8'h61;        memory[25768] <=  8'h63;        memory[25769] <=  8'h61;        memory[25770] <=  8'h74;        memory[25771] <=  8'h79;        memory[25772] <=  8'h73;        memory[25773] <=  8'h6e;        memory[25774] <=  8'h63;        memory[25775] <=  8'h74;        memory[25776] <=  8'h61;        memory[25777] <=  8'h6e;        memory[25778] <=  8'h62;        memory[25779] <=  8'h61;        memory[25780] <=  8'h63;        memory[25781] <=  8'h72;        memory[25782] <=  8'h6e;        memory[25783] <=  8'h74;        memory[25784] <=  8'h61;        memory[25785] <=  8'h62;        memory[25786] <=  8'h74;        memory[25787] <=  8'h6e;        memory[25788] <=  8'h61;        memory[25789] <=  8'h72;        memory[25790] <=  8'h62;        memory[25791] <=  8'h78;        memory[25792] <=  8'h74;        memory[25793] <=  8'h61;        memory[25794] <=  8'h72;        memory[25795] <=  8'h62;        memory[25796] <=  8'h61;        memory[25797] <=  8'h72;        memory[25798] <=  8'h74;        memory[25799] <=  8'h74;        memory[25800] <=  8'h62;        memory[25801] <=  8'h61;        memory[25802] <=  8'h72;        memory[25803] <=  8'h74;        memory[25804] <=  8'h78;        memory[25805] <=  8'h61;        memory[25806] <=  8'h74;        memory[25807] <=  8'h6b;        memory[25808] <=  8'h73;        memory[25809] <=  8'h68;        memory[25810] <=  8'h63;        memory[25811] <=  8'h66;        memory[25812] <=  8'h69;        memory[25813] <=  8'h77;        memory[25814] <=  8'h68;        memory[25815] <=  8'h61;        memory[25816] <=  8'h74;        memory[25817] <=  8'h61;        memory[25818] <=  8'h6e;        memory[25819] <=  8'h61;        memory[25820] <=  8'h62;        memory[25821] <=  8'h61;        memory[25822] <=  8'h63;        memory[25823] <=  8'h61;        memory[25824] <=  8'h74;        memory[25825] <=  8'h61;        memory[25826] <=  8'h62;        memory[25827] <=  8'h61;        memory[25828] <=  8'h72;        memory[25829] <=  8'h63;        memory[25830] <=  8'h61;        memory[25831] <=  8'h68;        memory[25832] <=  8'h64;        memory[25833] <=  8'h75;        memory[25834] <=  8'h63;        memory[25835] <=  8'h74;        memory[25836] <=  8'h61;        memory[25837] <=  8'h64;        memory[25838] <=  8'h61;        memory[25839] <=  8'h61;        memory[25840] <=  8'h63;        memory[25841] <=  8'h61;        memory[25842] <=  8'h72;        memory[25843] <=  8'h63;        memory[25844] <=  8'h74;        memory[25845] <=  8'h72;        memory[25846] <=  8'h63;        memory[25847] <=  8'h61;        memory[25848] <=  8'h74;        memory[25849] <=  8'h72;        memory[25850] <=  8'h63;        memory[25851] <=  8'h61;        memory[25852] <=  8'h74;        memory[25853] <=  8'h63;        memory[25854] <=  8'h62;        memory[25855] <=  8'h61;        memory[25856] <=  8'h74;        memory[25857] <=  8'h62;        memory[25858] <=  8'h72;        memory[25859] <=  8'h63;        memory[25860] <=  8'h61;        memory[25861] <=  8'h74;        memory[25862] <=  8'h72;        memory[25863] <=  8'h6e;        memory[25864] <=  8'h62;        memory[25865] <=  8'h61;        memory[25866] <=  8'h63;        memory[25867] <=  8'h61;        memory[25868] <=  8'h74;        memory[25869] <=  8'h79;        memory[25870] <=  8'h73;        memory[25871] <=  8'h6e;        memory[25872] <=  8'h63;        memory[25873] <=  8'h74;        memory[25874] <=  8'h61;        memory[25875] <=  8'h6e;        memory[25876] <=  8'h62;        memory[25877] <=  8'h61;        memory[25878] <=  8'h63;        memory[25879] <=  8'h72;        memory[25880] <=  8'h6e;        memory[25881] <=  8'h74;        memory[25882] <=  8'h61;        memory[25883] <=  8'h62;        memory[25884] <=  8'h74;        memory[25885] <=  8'h6e;        memory[25886] <=  8'h61;        memory[25887] <=  8'h72;        memory[25888] <=  8'h62;        memory[25889] <=  8'h78;        memory[25890] <=  8'h74;        memory[25891] <=  8'h61;        memory[25892] <=  8'h72;        memory[25893] <=  8'h64;        memory[25894] <=  8'h66;        memory[25895] <=  8'h73;        memory[25896] <=  8'h67;        memory[25897] <=  8'h76;        memory[25898] <=  8'h68;        memory[25899] <=  8'h62;        memory[25900] <=  8'h6b;        memory[25901] <=  8'h6a;        memory[25902] <=  8'h6e;        memory[25903] <=  8'h6d;        memory[25904] <=  8'h62;        memory[25905] <=  8'h76;        memory[25906] <=  8'h78;        memory[25907] <=  8'h63;        memory[25908] <=  8'h73;        memory[25909] <=  8'h66;        memory[25910] <=  8'h72;        memory[25911] <=  8'h74;        memory[25912] <=  8'h79;        memory[25913] <=  8'h75;        memory[25914] <=  8'h6a;        memory[25915] <=  8'h6e;        memory[25916] <=  8'h62;        memory[25917] <=  8'h76;        memory[25918] <=  8'h63;        memory[25919] <=  8'h64;        memory[25920] <=  8'h74;        memory[25921] <=  8'h79;        memory[25922] <=  8'h75;        memory[25923] <=  8'h69;        memory[25924] <=  8'h6b;        memory[25925] <=  8'h6d;        memory[25926] <=  8'h6e;        memory[25927] <=  8'h62;        memory[25928] <=  8'h76;        memory[25929] <=  8'h63;        memory[25930] <=  8'h78;        memory[25931] <=  8'h73;        memory[25932] <=  8'h64;        memory[25933] <=  8'h72;        memory[25934] <=  8'h74;        memory[25935] <=  8'h79;        memory[25936] <=  8'h75;        memory[25937] <=  8'h69;        memory[25938] <=  8'h6b;        memory[25939] <=  8'h6d;        memory[25940] <=  8'h6e;        memory[25941] <=  8'h62;        memory[25942] <=  8'h76;        memory[25943] <=  8'h63;        memory[25944] <=  8'h73;        memory[25945] <=  8'h77;        memory[25946] <=  8'h33;        memory[25947] <=  8'h34;        memory[25948] <=  8'h35;        memory[25949] <=  8'h36;        memory[25950] <=  8'h37;        memory[25951] <=  8'h38;        memory[25952] <=  8'h69;        memory[25953] <=  8'h6b;        memory[25954] <=  8'h6d;        memory[25955] <=  8'h6e;        memory[25956] <=  8'h62;        memory[25957] <=  8'h76;        memory[25958] <=  8'h63;        memory[25959] <=  8'h64;        memory[25960] <=  8'h65;        memory[25961] <=  8'h72;        memory[25962] <=  8'h36;        memory[25963] <=  8'h37;        memory[25964] <=  8'h38;        memory[25965] <=  8'h69;        memory[25966] <=  8'h6f;        memory[25967] <=  8'h6b;        memory[25968] <=  8'h6a;        memory[25969] <=  8'h6e;        memory[25970] <=  8'h62;        memory[25971] <=  8'h76;        memory[25972] <=  8'h63;        memory[25973] <=  8'h64;        memory[25974] <=  8'h72;        memory[25975] <=  8'h74;        memory[25976] <=  8'h79;        memory[25977] <=  8'h75;        memory[25978] <=  8'h73;        memory[25979] <=  8'h6a;        memory[25980] <=  8'h63;        memory[25981] <=  8'h6e;        memory[25982] <=  8'h62;        memory[25983] <=  8'h64;        memory[25984] <=  8'h66;        memory[25985] <=  8'h73;        memory[25986] <=  8'h74;        memory[25987] <=  8'h79;        memory[25988] <=  8'h75;        memory[25989] <=  8'h61;        memory[25990] <=  8'h69;        memory[25991] <=  8'h6b;        memory[25992] <=  8'h78;        memory[25993] <=  8'h6d;        memory[25994] <=  8'h6e;        memory[25995] <=  8'h73;        memory[25996] <=  8'h6a;        memory[25997] <=  8'h6f;        memory[25998] <=  8'h64;        memory[25999] <=  8'h6c;        memory[26000] <=  8'h63;        memory[26001] <=  8'h78;        memory[26002] <=  8'h62;        memory[26003] <=  8'h61;        memory[26004] <=  8'h72;        memory[26005] <=  8'h74;        memory[26006] <=  8'h78;        memory[26007] <=  8'h61;        memory[26008] <=  8'h74;        memory[26009] <=  8'h6b;        memory[26010] <=  8'h73;        memory[26011] <=  8'h68;        memory[26012] <=  8'h63;        memory[26013] <=  8'h66;        memory[26014] <=  8'h69;        memory[26015] <=  8'h77;        memory[26016] <=  8'h68;        memory[26017] <=  8'h61;        memory[26018] <=  8'h74;        memory[26019] <=  8'h61;        memory[26020] <=  8'h6e;        memory[26021] <=  8'h61;        memory[26022] <=  8'h62;        memory[26023] <=  8'h61;        memory[26024] <=  8'h63;        memory[26025] <=  8'h61;        memory[26026] <=  8'h74;        memory[26027] <=  8'h61;        memory[26028] <=  8'h62;        memory[26029] <=  8'h61;        memory[26030] <=  8'h72;        memory[26031] <=  8'h63;        memory[26032] <=  8'h61;        memory[26033] <=  8'h68;        memory[26034] <=  8'h64;        memory[26035] <=  8'h75;        memory[26036] <=  8'h63;        memory[26037] <=  8'h74;        memory[26038] <=  8'h61;        memory[26039] <=  8'h64;        memory[26040] <=  8'h61;        memory[26041] <=  8'h61;        memory[26042] <=  8'h63;        memory[26043] <=  8'h61;        memory[26044] <=  8'h72;        memory[26045] <=  8'h62;        memory[26046] <=  8'h61;        memory[26047] <=  8'h72;        memory[26048] <=  8'h74;        memory[26049] <=  8'h78;        memory[26050] <=  8'h61;        memory[26051] <=  8'h74;        memory[26052] <=  8'h6b;        memory[26053] <=  8'h73;        memory[26054] <=  8'h68;        memory[26055] <=  8'h63;        memory[26056] <=  8'h66;        memory[26057] <=  8'h69;        memory[26058] <=  8'h77;        memory[26059] <=  8'h68;        memory[26060] <=  8'h61;        memory[26061] <=  8'h74;        memory[26062] <=  8'h61;        memory[26063] <=  8'h6e;        memory[26064] <=  8'h61;        memory[26065] <=  8'h62;        memory[26066] <=  8'h61;        memory[26067] <=  8'h63;        memory[26068] <=  8'h61;        memory[26069] <=  8'h74;        memory[26070] <=  8'h61;        memory[26071] <=  8'h62;        memory[26072] <=  8'h61;        memory[26073] <=  8'h72;        memory[26074] <=  8'h63;        memory[26075] <=  8'h61;        memory[26076] <=  8'h68;        memory[26077] <=  8'h64;        memory[26078] <=  8'h75;        memory[26079] <=  8'h63;        memory[26080] <=  8'h74;        memory[26081] <=  8'h61;        memory[26082] <=  8'h64;        memory[26083] <=  8'h61;        memory[26084] <=  8'h61;        memory[26085] <=  8'h63;        memory[26086] <=  8'h61;        memory[26087] <=  8'h72;        memory[26088] <=  8'h62;        memory[26089] <=  8'h61;        memory[26090] <=  8'h72;        memory[26091] <=  8'h74;        memory[26092] <=  8'h78;        memory[26093] <=  8'h61;        memory[26094] <=  8'h74;        memory[26095] <=  8'h6b;        memory[26096] <=  8'h73;        memory[26097] <=  8'h68;        memory[26098] <=  8'h63;        memory[26099] <=  8'h66;        memory[26100] <=  8'h69;        memory[26101] <=  8'h77;        memory[26102] <=  8'h68;        memory[26103] <=  8'h61;        memory[26104] <=  8'h74;        memory[26105] <=  8'h61;        memory[26106] <=  8'h6e;        memory[26107] <=  8'h61;        memory[26108] <=  8'h62;        memory[26109] <=  8'h61;        memory[26110] <=  8'h63;        memory[26111] <=  8'h61;        memory[26112] <=  8'h74;        memory[26113] <=  8'h61;        memory[26114] <=  8'h62;        memory[26115] <=  8'h61;        memory[26116] <=  8'h72;        memory[26117] <=  8'h63;        memory[26118] <=  8'h61;        memory[26119] <=  8'h68;        memory[26120] <=  8'h64;        memory[26121] <=  8'h75;        memory[26122] <=  8'h63;        memory[26123] <=  8'h74;        memory[26124] <=  8'h61;        memory[26125] <=  8'h64;        memory[26126] <=  8'h61;        memory[26127] <=  8'h61;        memory[26128] <=  8'h63;        memory[26129] <=  8'h61;        memory[26130] <=  8'h72;        memory[26131] <=  8'h62;        memory[26132] <=  8'h61;        memory[26133] <=  8'h72;        memory[26134] <=  8'h74;        memory[26135] <=  8'h78;        memory[26136] <=  8'h61;        memory[26137] <=  8'h74;        memory[26138] <=  8'h6b;        memory[26139] <=  8'h73;        memory[26140] <=  8'h68;        memory[26141] <=  8'h63;        memory[26142] <=  8'h66;        memory[26143] <=  8'h69;        memory[26144] <=  8'h77;        memory[26145] <=  8'h68;        memory[26146] <=  8'h61;        memory[26147] <=  8'h74;        memory[26148] <=  8'h61;        memory[26149] <=  8'h6e;        memory[26150] <=  8'h61;        memory[26151] <=  8'h62;        memory[26152] <=  8'h61;        memory[26153] <=  8'h63;        memory[26154] <=  8'h61;        memory[26155] <=  8'h74;        memory[26156] <=  8'h61;        memory[26157] <=  8'h62;        memory[26158] <=  8'h61;        memory[26159] <=  8'h72;        memory[26160] <=  8'h63;        memory[26161] <=  8'h61;        memory[26162] <=  8'h68;        memory[26163] <=  8'h64;        memory[26164] <=  8'h75;        memory[26165] <=  8'h63;        memory[26166] <=  8'h74;        memory[26167] <=  8'h61;        memory[26168] <=  8'h64;        memory[26169] <=  8'h61;        memory[26170] <=  8'h61;        memory[26171] <=  8'h63;        memory[26172] <=  8'h61;        memory[26173] <=  8'h72;        memory[26174] <=  8'h62;        memory[26175] <=  8'h61;        memory[26176] <=  8'h72;        memory[26177] <=  8'h74;        memory[26178] <=  8'h78;        memory[26179] <=  8'h61;        memory[26180] <=  8'h74;        memory[26181] <=  8'h6b;        memory[26182] <=  8'h73;        memory[26183] <=  8'h68;        memory[26184] <=  8'h63;        memory[26185] <=  8'h66;        memory[26186] <=  8'h69;        memory[26187] <=  8'h77;        memory[26188] <=  8'h68;        memory[26189] <=  8'h61;        memory[26190] <=  8'h74;        memory[26191] <=  8'h61;        memory[26192] <=  8'h6e;        memory[26193] <=  8'h61;        memory[26194] <=  8'h62;        memory[26195] <=  8'h61;        memory[26196] <=  8'h63;        memory[26197] <=  8'h61;        memory[26198] <=  8'h74;        memory[26199] <=  8'h61;        memory[26200] <=  8'h62;        memory[26201] <=  8'h61;        memory[26202] <=  8'h72;        memory[26203] <=  8'h63;        memory[26204] <=  8'h61;        memory[26205] <=  8'h68;        memory[26206] <=  8'h64;        memory[26207] <=  8'h75;        memory[26208] <=  8'h63;        memory[26209] <=  8'h74;        memory[26210] <=  8'h61;        memory[26211] <=  8'h64;        memory[26212] <=  8'h61;        memory[26213] <=  8'h61;        memory[26214] <=  8'h63;        memory[26215] <=  8'h61;        memory[26216] <=  8'h72;        memory[26217] <=  8'h62;        memory[26218] <=  8'h61;        memory[26219] <=  8'h72;        memory[26220] <=  8'h74;        memory[26221] <=  8'h78;        memory[26222] <=  8'h61;        memory[26223] <=  8'h74;        memory[26224] <=  8'h6b;        memory[26225] <=  8'h73;        memory[26226] <=  8'h68;        memory[26227] <=  8'h63;        memory[26228] <=  8'h66;        memory[26229] <=  8'h69;        memory[26230] <=  8'h77;        memory[26231] <=  8'h68;        memory[26232] <=  8'h61;        memory[26233] <=  8'h74;        memory[26234] <=  8'h61;        memory[26235] <=  8'h6e;        memory[26236] <=  8'h61;        memory[26237] <=  8'h62;        memory[26238] <=  8'h61;        memory[26239] <=  8'h63;        memory[26240] <=  8'h61;        memory[26241] <=  8'h74;        memory[26242] <=  8'h61;        memory[26243] <=  8'h62;        memory[26244] <=  8'h61;        memory[26245] <=  8'h72;        memory[26246] <=  8'h63;        memory[26247] <=  8'h61;        memory[26248] <=  8'h68;        memory[26249] <=  8'h64;        memory[26250] <=  8'h75;        memory[26251] <=  8'h63;        memory[26252] <=  8'h74;        memory[26253] <=  8'h61;        memory[26254] <=  8'h64;        memory[26255] <=  8'h61;        memory[26256] <=  8'h61;        memory[26257] <=  8'h63;        memory[26258] <=  8'h61;        memory[26259] <=  8'h72;        memory[26260] <=  8'h62;        memory[26261] <=  8'h61;        memory[26262] <=  8'h72;        memory[26263] <=  8'h74;        memory[26264] <=  8'h78;        memory[26265] <=  8'h61;        memory[26266] <=  8'h74;        memory[26267] <=  8'h6b;        memory[26268] <=  8'h73;        memory[26269] <=  8'h68;        memory[26270] <=  8'h63;        memory[26271] <=  8'h66;        memory[26272] <=  8'h69;        memory[26273] <=  8'h77;        memory[26274] <=  8'h68;        memory[26275] <=  8'h61;        memory[26276] <=  8'h74;        memory[26277] <=  8'h61;        memory[26278] <=  8'h6e;        memory[26279] <=  8'h61;        memory[26280] <=  8'h62;        memory[26281] <=  8'h61;        memory[26282] <=  8'h63;        memory[26283] <=  8'h61;        memory[26284] <=  8'h74;        memory[26285] <=  8'h61;        memory[26286] <=  8'h62;        memory[26287] <=  8'h61;        memory[26288] <=  8'h72;        memory[26289] <=  8'h63;        memory[26290] <=  8'h61;        memory[26291] <=  8'h68;        memory[26292] <=  8'h64;        memory[26293] <=  8'h75;        memory[26294] <=  8'h63;        memory[26295] <=  8'h74;        memory[26296] <=  8'h61;        memory[26297] <=  8'h64;        memory[26298] <=  8'h61;        memory[26299] <=  8'h61;        memory[26300] <=  8'h63;        memory[26301] <=  8'h61;        memory[26302] <=  8'h72;        memory[26303] <=  8'h62;        memory[26304] <=  8'h61;        memory[26305] <=  8'h72;        memory[26306] <=  8'h74;        memory[26307] <=  8'h78;        memory[26308] <=  8'h61;        memory[26309] <=  8'h74;        memory[26310] <=  8'h6b;        memory[26311] <=  8'h73;        memory[26312] <=  8'h68;        memory[26313] <=  8'h63;        memory[26314] <=  8'h66;        memory[26315] <=  8'h69;        memory[26316] <=  8'h77;        memory[26317] <=  8'h68;        memory[26318] <=  8'h61;        memory[26319] <=  8'h74;        memory[26320] <=  8'h61;        memory[26321] <=  8'h6e;        memory[26322] <=  8'h61;        memory[26323] <=  8'h62;        memory[26324] <=  8'h61;        memory[26325] <=  8'h63;        memory[26326] <=  8'h61;        memory[26327] <=  8'h74;        memory[26328] <=  8'h61;        memory[26329] <=  8'h62;        memory[26330] <=  8'h61;        memory[26331] <=  8'h72;        memory[26332] <=  8'h63;        memory[26333] <=  8'h61;        memory[26334] <=  8'h68;        memory[26335] <=  8'h64;        memory[26336] <=  8'h75;        memory[26337] <=  8'h63;        memory[26338] <=  8'h74;        memory[26339] <=  8'h61;        memory[26340] <=  8'h64;        memory[26341] <=  8'h61;        memory[26342] <=  8'h61;        memory[26343] <=  8'h63;        memory[26344] <=  8'h61;        memory[26345] <=  8'h72;        memory[26346] <=  8'h62;        memory[26347] <=  8'h61;        memory[26348] <=  8'h72;        memory[26349] <=  8'h74;        memory[26350] <=  8'h78;        memory[26351] <=  8'h61;        memory[26352] <=  8'h74;        memory[26353] <=  8'h6b;        memory[26354] <=  8'h73;        memory[26355] <=  8'h68;        memory[26356] <=  8'h63;        memory[26357] <=  8'h66;        memory[26358] <=  8'h69;        memory[26359] <=  8'h77;        memory[26360] <=  8'h68;        memory[26361] <=  8'h61;        memory[26362] <=  8'h74;        memory[26363] <=  8'h61;        memory[26364] <=  8'h6e;        memory[26365] <=  8'h61;        memory[26366] <=  8'h62;        memory[26367] <=  8'h61;        memory[26368] <=  8'h63;        memory[26369] <=  8'h61;        memory[26370] <=  8'h74;        memory[26371] <=  8'h61;        memory[26372] <=  8'h62;        memory[26373] <=  8'h61;        memory[26374] <=  8'h72;        memory[26375] <=  8'h63;        memory[26376] <=  8'h61;        memory[26377] <=  8'h68;        memory[26378] <=  8'h64;        memory[26379] <=  8'h75;        memory[26380] <=  8'h63;        memory[26381] <=  8'h74;        memory[26382] <=  8'h61;        memory[26383] <=  8'h64;        memory[26384] <=  8'h61;        memory[26385] <=  8'h61;        memory[26386] <=  8'h63;        memory[26387] <=  8'h61;        memory[26388] <=  8'h72;        memory[26389] <=  8'h62;        memory[26390] <=  8'h61;        memory[26391] <=  8'h72;        memory[26392] <=  8'h74;        memory[26393] <=  8'h74;        memory[26394] <=  8'h62;        memory[26395] <=  8'h61;        memory[26396] <=  8'h72;        memory[26397] <=  8'h74;        memory[26398] <=  8'h78;        memory[26399] <=  8'h61;        memory[26400] <=  8'h74;        memory[26401] <=  8'h6b;        memory[26402] <=  8'h73;        memory[26403] <=  8'h68;        memory[26404] <=  8'h63;        memory[26405] <=  8'h66;        memory[26406] <=  8'h69;        memory[26407] <=  8'h77;        memory[26408] <=  8'h68;        memory[26409] <=  8'h61;        memory[26410] <=  8'h74;        memory[26411] <=  8'h61;        memory[26412] <=  8'h6e;        memory[26413] <=  8'h61;        memory[26414] <=  8'h62;        memory[26415] <=  8'h61;        memory[26416] <=  8'h63;        memory[26417] <=  8'h61;        memory[26418] <=  8'h74;        memory[26419] <=  8'h61;        memory[26420] <=  8'h62;        memory[26421] <=  8'h61;        memory[26422] <=  8'h72;        memory[26423] <=  8'h63;        memory[26424] <=  8'h61;        memory[26425] <=  8'h68;        memory[26426] <=  8'h64;        memory[26427] <=  8'h75;        memory[26428] <=  8'h63;        memory[26429] <=  8'h74;        memory[26430] <=  8'h61;        memory[26431] <=  8'h64;        memory[26432] <=  8'h61;        memory[26433] <=  8'h61;        memory[26434] <=  8'h63;        memory[26435] <=  8'h61;        memory[26436] <=  8'h72;        memory[26437] <=  8'h63;        memory[26438] <=  8'h74;        memory[26439] <=  8'h72;        memory[26440] <=  8'h63;        memory[26441] <=  8'h61;        memory[26442] <=  8'h74;        memory[26443] <=  8'h72;        memory[26444] <=  8'h63;        memory[26445] <=  8'h61;        memory[26446] <=  8'h74;        memory[26447] <=  8'h63;        memory[26448] <=  8'h62;        memory[26449] <=  8'h61;        memory[26450] <=  8'h74;        memory[26451] <=  8'h62;        memory[26452] <=  8'h72;        memory[26453] <=  8'h63;        memory[26454] <=  8'h61;        memory[26455] <=  8'h72;        memory[26456] <=  8'h62;        memory[26457] <=  8'h78;        memory[26458] <=  8'h74;        memory[26459] <=  8'h61;        memory[26460] <=  8'h72;        memory[26461] <=  8'h64;        memory[26462] <=  8'h66;        memory[26463] <=  8'h73;        memory[26464] <=  8'h67;        memory[26465] <=  8'h76;        memory[26466] <=  8'h68;        memory[26467] <=  8'h62;        memory[26468] <=  8'h6b;        memory[26469] <=  8'h6a;        memory[26470] <=  8'h6e;        memory[26471] <=  8'h6d;        memory[26472] <=  8'h62;        memory[26473] <=  8'h76;        memory[26474] <=  8'h78;        memory[26475] <=  8'h63;        memory[26476] <=  8'h73;        memory[26477] <=  8'h66;        memory[26478] <=  8'h72;        memory[26479] <=  8'h74;        memory[26480] <=  8'h79;        memory[26481] <=  8'h75;        memory[26482] <=  8'h6a;        memory[26483] <=  8'h6e;        memory[26484] <=  8'h62;        memory[26485] <=  8'h76;        memory[26486] <=  8'h63;        memory[26487] <=  8'h64;        memory[26488] <=  8'h74;        memory[26489] <=  8'h79;        memory[26490] <=  8'h75;        memory[26491] <=  8'h69;        memory[26492] <=  8'h6b;        memory[26493] <=  8'h6d;        memory[26494] <=  8'h6e;        memory[26495] <=  8'h62;        memory[26496] <=  8'h76;        memory[26497] <=  8'h63;        memory[26498] <=  8'h78;        memory[26499] <=  8'h73;        memory[26500] <=  8'h64;        memory[26501] <=  8'h72;        memory[26502] <=  8'h74;        memory[26503] <=  8'h79;        memory[26504] <=  8'h75;        memory[26505] <=  8'h69;        memory[26506] <=  8'h6b;        memory[26507] <=  8'h6d;        memory[26508] <=  8'h6e;        memory[26509] <=  8'h62;        memory[26510] <=  8'h76;        memory[26511] <=  8'h63;        memory[26512] <=  8'h73;        memory[26513] <=  8'h77;        memory[26514] <=  8'h33;        memory[26515] <=  8'h34;        memory[26516] <=  8'h35;        memory[26517] <=  8'h36;        memory[26518] <=  8'h37;        memory[26519] <=  8'h38;        memory[26520] <=  8'h69;        memory[26521] <=  8'h6b;        memory[26522] <=  8'h6d;        memory[26523] <=  8'h6e;        memory[26524] <=  8'h62;        memory[26525] <=  8'h76;        memory[26526] <=  8'h63;        memory[26527] <=  8'h64;        memory[26528] <=  8'h65;        memory[26529] <=  8'h72;        memory[26530] <=  8'h36;        memory[26531] <=  8'h37;        memory[26532] <=  8'h38;        memory[26533] <=  8'h69;        memory[26534] <=  8'h6f;        memory[26535] <=  8'h6b;        memory[26536] <=  8'h6a;        memory[26537] <=  8'h6e;        memory[26538] <=  8'h62;        memory[26539] <=  8'h76;        memory[26540] <=  8'h63;        memory[26541] <=  8'h64;        memory[26542] <=  8'h72;        memory[26543] <=  8'h74;        memory[26544] <=  8'h79;        memory[26545] <=  8'h75;        memory[26546] <=  8'h73;        memory[26547] <=  8'h6a;        memory[26548] <=  8'h63;        memory[26549] <=  8'h6e;        memory[26550] <=  8'h62;        memory[26551] <=  8'h64;        memory[26552] <=  8'h66;        memory[26553] <=  8'h73;        memory[26554] <=  8'h74;        memory[26555] <=  8'h79;        memory[26556] <=  8'h75;        memory[26557] <=  8'h61;        memory[26558] <=  8'h69;        memory[26559] <=  8'h6b;        memory[26560] <=  8'h78;        memory[26561] <=  8'h6d;        memory[26562] <=  8'h6e;        memory[26563] <=  8'h73;        memory[26564] <=  8'h6a;        memory[26565] <=  8'h6f;        memory[26566] <=  8'h64;        memory[26567] <=  8'h6c;        memory[26568] <=  8'h63;        memory[26569] <=  8'h78;        memory[26570] <=  8'h2c;        memory[26571] <=  8'h6d;        memory[26572] <=  8'h73;        memory[26573] <=  8'h6b;        memory[26574] <=  8'h64;        memory[26575] <=  8'h6c;        memory[26576] <=  8'h70;        memory[26577] <=  8'h5b;        memory[26578] <=  8'h3b;        memory[26579] <=  8'h73;        memory[26580] <=  8'h6c;        memory[26581] <=  8'h64;        memory[26582] <=  8'h70;        memory[26583] <=  8'h76;        memory[26584] <=  8'h63;        memory[26585] <=  8'h5b;        memory[26586] <=  8'h78;        memory[26587] <=  8'h76;        memory[26588] <=  8'h63;        memory[26589] <=  8'h5b;        memory[26590] <=  8'h78;        memory[26591] <=  8'h70;        memory[26592] <=  8'h6f;        memory[26593] <=  8'h20;        memory[26594] <=  8'h62;        memory[26595] <=  8'h61;        memory[26596] <=  8'h72;        memory[26597] <=  8'h74;        memory[26598] <=  8'h74;        memory[26599] <=  8'h62;        memory[26600] <=  8'h61;        memory[26601] <=  8'h72;        memory[26602] <=  8'h74;        memory[26603] <=  8'h78;        memory[26604] <=  8'h61;        memory[26605] <=  8'h74;        memory[26606] <=  8'h6b;        memory[26607] <=  8'h73;        memory[26608] <=  8'h68;        memory[26609] <=  8'h63;        memory[26610] <=  8'h66;        memory[26611] <=  8'h69;        memory[26612] <=  8'h77;        memory[26613] <=  8'h68;        memory[26614] <=  8'h61;        memory[26615] <=  8'h69;        memory[26616] <=  8'h6a;        memory[26617] <=  8'h78;        memory[26618] <=  8'h5d;        memory[26619] <=  8'h65;        memory[26620] <=  8'h6b;        memory[26621] <=  8'h6f;        memory[26622] <=  8'h39;        memory[26623] <=  8'h64;        memory[26624] <=  8'h75;        memory[26625] <=  8'h38;        memory[26626] <=  8'h79;        memory[26627] <=  8'h20;        memory[26628] <=  8'h37;        memory[26629] <=  8'h63;        memory[26630] <=  8'h67;        memory[26631] <=  8'h78;        memory[26632] <=  8'h63;        memory[26633] <=  8'h75;        memory[26634] <=  8'h68;        memory[26635] <=  8'h69;        memory[26636] <=  8'h6a;        memory[26637] <=  8'h77;        memory[26638] <=  8'h69;        memory[26639] <=  8'h64;        memory[26640] <=  8'h66;        memory[26641] <=  8'h68;        memory[26642] <=  8'h75;        memory[26643] <=  8'h76;        memory[26644] <=  8'h64;        memory[26645] <=  8'h62;        memory[26646] <=  8'h66;        memory[26647] <=  8'h6a;        memory[26648] <=  8'h6e;        memory[26649] <=  8'h6b;        memory[26650] <=  8'h6a;        memory[26651] <=  8'h65;        memory[26652] <=  8'h38;        memory[26653] <=  8'h66;        memory[26654] <=  8'h37;        memory[26655] <=  8'h67;        memory[26656] <=  8'h79;        memory[26657] <=  8'h76;        memory[26658] <=  8'h63;        memory[26659] <=  8'h68;        memory[26660] <=  8'h69;        memory[26661] <=  8'h6a;        memory[26662] <=  8'h33;        memory[26663] <=  8'h65;        memory[26664] <=  8'h67;        memory[26665] <=  8'h79;        memory[26666] <=  8'h72;        memory[26667] <=  8'h64;        memory[26668] <=  8'h62;        memory[26669] <=  8'h6e;        memory[26670] <=  8'h63;        memory[26671] <=  8'h7a;        memory[26672] <=  8'h6a;        memory[26673] <=  8'h6f;        memory[26674] <=  8'h66;        memory[26675] <=  8'h78;        memory[26676] <=  8'h6a;        memory[26677] <=  8'h69;        memory[26678] <=  8'h63;        memory[26679] <=  8'h68;        memory[26680] <=  8'h62;        memory[26681] <=  8'h6e;        memory[26682] <=  8'h6d;        memory[26683] <=  8'h63;        memory[26684] <=  8'h73;        memory[26685] <=  8'h6c;        memory[26686] <=  8'h6b;        memory[26687] <=  8'h6a;        memory[26688] <=  8'h69;        memory[26689] <=  8'h68;        memory[26690] <=  8'h76;        memory[26691] <=  8'h75;        memory[26692] <=  8'h69;        memory[26693] <=  8'h64;        memory[26694] <=  8'h68;        memory[26695] <=  8'h75;        memory[26696] <=  8'h67;        memory[26697] <=  8'h79;        memory[26698] <=  8'h62;        memory[26699] <=  8'h68;        memory[26700] <=  8'h65;        memory[26701] <=  8'h6a;        memory[26702] <=  8'h72;        memory[26703] <=  8'h6b;        memory[26704] <=  8'h6a;        memory[26705] <=  8'h6f;        memory[26706] <=  8'h64;        memory[26707] <=  8'h67;        memory[26708] <=  8'h69;        memory[26709] <=  8'h75;        memory[26710] <=  8'h69;        memory[26711] <=  8'h67;        memory[26712] <=  8'h76;        memory[26713] <=  8'h79;        memory[26714] <=  8'h75;        memory[26715] <=  8'h67;        memory[26716] <=  8'h78;        memory[26717] <=  8'h68;        memory[26718] <=  8'h63;        memory[26719] <=  8'h20;        memory[26720] <=  8'h20;        memory[26721] <=  8'h20;        memory[26722] <=  8'h78;        memory[26723] <=  8'h76;        memory[26724] <=  8'h20;        memory[26725] <=  8'h63;        memory[26726] <=  8'h78;        memory[26727] <=  8'h67;        memory[26728] <=  8'h79;        memory[26729] <=  8'h63;        memory[26730] <=  8'h75;        memory[26731] <=  8'h68;        memory[26732] <=  8'h6a;        memory[26733] <=  8'h6b;        memory[26734] <=  8'h61;        memory[26735] <=  8'h6c;        memory[26736] <=  8'h78;        memory[26737] <=  8'h76;        memory[26738] <=  8'h70;        memory[26739] <=  8'h6f;        memory[26740] <=  8'h69;        memory[26741] <=  8'h6a;        memory[26742] <=  8'h69;        memory[26743] <=  8'h68;        memory[26744] <=  8'h6a;        memory[26745] <=  8'h62;        memory[26746] <=  8'h77;        memory[26747] <=  8'h65;        memory[26748] <=  8'h6e;        memory[26749] <=  8'h61;        memory[26750] <=  8'h66;        memory[26751] <=  8'h6d;        memory[26752] <=  8'h64;        memory[26753] <=  8'h6b;        memory[26754] <=  8'h6d;        memory[26755] <=  8'h76;        memory[26756] <=  8'h6c;        memory[26757] <=  8'h63;        memory[26758] <=  8'h6f;        memory[26759] <=  8'h64;        memory[26760] <=  8'h69;        memory[26761] <=  8'h75;        memory[26762] <=  8'h68;        memory[26763] <=  8'h73;        memory[26764] <=  8'h66;        memory[26765] <=  8'h65;        memory[26766] <=  8'h62;        memory[26767] <=  8'h6e;        memory[26768] <=  8'h64;        memory[26769] <=  8'h73;        memory[26770] <=  8'h63;        memory[26771] <=  8'h6b;        memory[26772] <=  8'h20;        memory[26773] <=  8'h78;        memory[26774] <=  8'h6a;        memory[26775] <=  8'h78;        memory[26776] <=  8'h63;        memory[26777] <=  8'h73;        memory[26778] <=  8'h64;        memory[26779] <=  8'h66;        memory[26780] <=  8'h6b;        memory[26781] <=  8'h64;        memory[26782] <=  8'h6e;        memory[26783] <=  8'h6d;        memory[26784] <=  8'h64;        memory[26785] <=  8'h73;        memory[26786] <=  8'h63;        memory[26787] <=  8'h6b;        memory[26788] <=  8'h78;        memory[26789] <=  8'h6c;        memory[26790] <=  8'h6f;        memory[26791] <=  8'h66;        memory[26792] <=  8'h6a;        memory[26793] <=  8'h69;        memory[26794] <=  8'h61;        memory[26795] <=  8'h62;        memory[26796] <=  8'h6e;        memory[26797] <=  8'h20;        memory[26798] <=  8'h78;        memory[26799] <=  8'h6b;        memory[26800] <=  8'h6d;        memory[26801] <=  8'h20;        memory[26802] <=  8'h6f;        memory[26803] <=  8'h63;        memory[26804] <=  8'h76;        memory[26805] <=  8'h73;        memory[26806] <=  8'h64;        memory[26807] <=  8'h69;        memory[26808] <=  8'h66;        memory[26809] <=  8'h68;        memory[26810] <=  8'h65;        memory[26811] <=  8'h71;        memory[26812] <=  8'h6a;        memory[26813] <=  8'h77;        memory[26814] <=  8'h62;        memory[26815] <=  8'h65;        memory[26816] <=  8'h6e;        memory[26817] <=  8'h20;        memory[26818] <=  8'h6d;        memory[26819] <=  8'h64;        memory[26820] <=  8'h73;        memory[26821] <=  8'h6c;        memory[26822] <=  8'h76;        memory[26823] <=  8'h6b;        memory[26824] <=  8'h63;        memory[26825] <=  8'h78;        memory[26826] <=  8'h20;        memory[26827] <=  8'h6f;        memory[26828] <=  8'h78;        memory[26829] <=  8'h69;        memory[26830] <=  8'h63;        memory[26831] <=  8'h6a;        memory[26832] <=  8'h76;        memory[26833] <=  8'h64;        memory[26834] <=  8'h66;        memory[26835] <=  8'h65;        memory[26836] <=  8'h71;        memory[26837] <=  8'h6e;        memory[26838] <=  8'h20;        memory[26839] <=  8'h64;        memory[26840] <=  8'h6d;        memory[26841] <=  8'h73;        memory[26842] <=  8'h6c;        memory[26843] <=  8'h63;        memory[26844] <=  8'h78;        memory[26845] <=  8'h6b;        memory[26846] <=  8'h20;        memory[26847] <=  8'h6f;        memory[26848] <=  8'h78;        memory[26849] <=  8'h63;        memory[26850] <=  8'h76;        memory[26851] <=  8'h6a;        memory[26852] <=  8'h64;        memory[26853] <=  8'h62;        memory[26854] <=  8'h71;        memory[26855] <=  8'h77;        memory[26856] <=  8'h65;        memory[26857] <=  8'h6e;        memory[26858] <=  8'h6d;        memory[26859] <=  8'h64;        memory[26860] <=  8'h6c;        memory[26861] <=  8'h73;        memory[26862] <=  8'h2c;        memory[26863] <=  8'h76;        memory[26864] <=  8'h63;        memory[26865] <=  8'h78;        memory[26866] <=  8'h20;        memory[26867] <=  8'h63;        memory[26868] <=  8'h6f;        memory[26869] <=  8'h69;        memory[26870] <=  8'h76;        memory[26871] <=  8'h68;        memory[26872] <=  8'h73;        memory[26873] <=  8'h64;        memory[26874] <=  8'h62;        memory[26875] <=  8'h71;        memory[26876] <=  8'h77;        memory[26877] <=  8'h65;        memory[26878] <=  8'h6e;        memory[26879] <=  8'h64;        memory[26880] <=  8'h6b;        memory[26881] <=  8'h73;        memory[26882] <=  8'h76;        memory[26883] <=  8'h6f;        memory[26884] <=  8'h63;        memory[26885] <=  8'h20;        memory[26886] <=  8'h76;        memory[26887] <=  8'h69;        memory[26888] <=  8'h75;        memory[26889] <=  8'h69;        memory[26890] <=  8'h68;        memory[26891] <=  8'h63;        memory[26892] <=  8'h78;        memory[26893] <=  8'h69;        memory[26894] <=  8'h6f;        memory[26895] <=  8'h76;        memory[26896] <=  8'h73;        memory[26897] <=  8'h64;        memory[26898] <=  8'h61;        memory[26899] <=  8'h64;        memory[26900] <=  8'h6e;        memory[26901] <=  8'h77;        memory[26902] <=  8'h71;        memory[26903] <=  8'h6b;        memory[26904] <=  8'h6c;        memory[26905] <=  8'h73;        memory[26906] <=  8'h76;        memory[26907] <=  8'h6e;        memory[26908] <=  8'h62;        memory[26909] <=  8'h20;        memory[26910] <=  8'h64;        memory[26911] <=  8'h66;        memory[26912] <=  8'h6a;        memory[26913] <=  8'h6b;        memory[26914] <=  8'h71;        memory[26915] <=  8'h64;        memory[26916] <=  8'h77;        memory[26917] <=  8'h65;        memory[26918] <=  8'h6e;        memory[26919] <=  8'h62;        memory[26920] <=  8'h20;        memory[26921] <=  8'h64;        memory[26922] <=  8'h73;        memory[26923] <=  8'h76;        memory[26924] <=  8'h68;        memory[26925] <=  8'h64;        memory[26926] <=  8'h61;        memory[26927] <=  8'h71;        memory[26928] <=  8'h77;        memory[26929] <=  8'h6a;        memory[26930] <=  8'h65;        memory[26931] <=  8'h6e;        memory[26932] <=  8'h64;        memory[26933] <=  8'h20;        memory[26934] <=  8'h61;        memory[26935] <=  8'h63;        memory[26936] <=  8'h62;        memory[26937] <=  8'h68;        memory[26938] <=  8'h64;        memory[26939] <=  8'h61;        memory[26940] <=  8'h77;        memory[26941] <=  8'h71;        memory[26942] <=  8'h6e;        memory[26943] <=  8'h20;        memory[26944] <=  8'h62;        memory[26945] <=  8'h73;        memory[26946] <=  8'h76;        memory[26947] <=  8'h61;        memory[26948] <=  8'h67;        memory[26949] <=  8'h76;        memory[26950] <=  8'h68;        memory[26951] <=  8'h67;        memory[26952] <=  8'h61;        memory[26953] <=  8'h73;        memory[26954] <=  8'h6a;        memory[26955] <=  8'h6b;        memory[26956] <=  8'h63;        memory[26957] <=  8'h78;        memory[26958] <=  8'h76;        memory[26959] <=  8'h6e;        memory[26960] <=  8'h73;        memory[26961] <=  8'h64;        memory[26962] <=  8'h20;        memory[26963] <=  8'h66;        memory[26964] <=  8'h62;        memory[26965] <=  8'h64;        memory[26966] <=  8'h61;        memory[26967] <=  8'h73;        memory[26968] <=  8'h76;        memory[26969] <=  8'h67;        memory[26970] <=  8'h63;        memory[26971] <=  8'h79;        memory[26972] <=  8'h7a;        memory[26973] <=  8'h78;        memory[26974] <=  8'h79;        memory[26975] <=  8'h75;        memory[26976] <=  8'h20;        memory[26977] <=  8'h69;        memory[26978] <=  8'h6a;        memory[26979] <=  8'h64;        memory[26980] <=  8'h66;        memory[26981] <=  8'h6b;        memory[26982] <=  8'h61;        memory[26983] <=  8'h64;        memory[26984] <=  8'h63;        memory[26985] <=  8'h78;        memory[26986] <=  8'h68;        memory[26987] <=  8'h20;        memory[26988] <=  8'h67;        memory[26989] <=  8'h61;        memory[26990] <=  8'h68;        memory[26991] <=  8'h75;        memory[26992] <=  8'h64;        memory[26993] <=  8'h73;        memory[26994] <=  8'h69;        memory[26995] <=  8'h6a;        memory[26996] <=  8'h61;        memory[26997] <=  8'h6b;        memory[26998] <=  8'h63;        memory[26999] <=  8'h62;        memory[27000] <=  8'h61;        memory[27001] <=  8'h72;        memory[27002] <=  8'h73;        memory[27003] <=  8'h68;        memory[27004] <=  8'h64;        memory[27005] <=  8'h66;        memory[27006] <=  8'h67;        memory[27007] <=  8'h73;        memory[27008] <=  8'h68;        memory[27009] <=  8'h64;        memory[27010] <=  8'h66;        memory[27011] <=  8'h68;        memory[27012] <=  8'h64;        memory[27013] <=  8'h6a;        memory[27014] <=  8'h68;        memory[27015] <=  8'h62;        memory[27016] <=  8'h67;        memory[27017] <=  8'h63;        memory[27018] <=  8'h61;        memory[27019] <=  8'h66;        memory[27020] <=  8'h73;        memory[27021] <=  8'h79;        memory[27022] <=  8'h67;        memory[27023] <=  8'h6b;        memory[27024] <=  8'h75;        memory[27025] <=  8'h64;        memory[27026] <=  8'h68;        memory[27027] <=  8'h62;        memory[27028] <=  8'h77;        memory[27029] <=  8'h76;        memory[27030] <=  8'h67;        memory[27031] <=  8'h61;        memory[27032] <=  8'h66;        memory[27033] <=  8'h64;        memory[27034] <=  8'h74;        memory[27035] <=  8'h75;        memory[27036] <=  8'h66;        memory[27037] <=  8'h79;        memory[27038] <=  8'h67;        memory[27039] <=  8'h69;        memory[27040] <=  8'h75;        memory[27041] <=  8'h68;        memory[27042] <=  8'h6c;        memory[27043] <=  8'h6a;        memory[27044] <=  8'h62;        memory[27045] <=  8'h6b;        memory[27046] <=  8'h68;        memory[27047] <=  8'h76;        memory[27048] <=  8'h67;        memory[27049] <=  8'h63;        memory[27050] <=  8'h66;        memory[27051] <=  8'h78;        memory[27052] <=  8'h64;        memory[27053] <=  8'h74;        memory[27054] <=  8'h75;        memory[27055] <=  8'h79;        memory[27056] <=  8'h69;        memory[27057] <=  8'h75;        memory[27058] <=  8'h68;        memory[27059] <=  8'h6c;        memory[27060] <=  8'h6a;        memory[27061] <=  8'h6b;        memory[27062] <=  8'h67;        memory[27063] <=  8'h6a;        memory[27064] <=  8'h63;        memory[27065] <=  8'h66;        memory[27066] <=  8'h68;        memory[27067] <=  8'h64;        memory[27068] <=  8'h67;        memory[27069] <=  8'h72;        memory[27070] <=  8'h79;        memory[27071] <=  8'h74;        memory[27072] <=  8'h66;        memory[27073] <=  8'h75;        memory[27074] <=  8'h79;        memory[27075] <=  8'h69;        memory[27076] <=  8'h68;        memory[27077] <=  8'h6c;        memory[27078] <=  8'h62;        memory[27079] <=  8'h6d;        memory[27080] <=  8'h76;        memory[27081] <=  8'h6e;        memory[27082] <=  8'h63;        memory[27083] <=  8'h66;        memory[27084] <=  8'h68;        memory[27085] <=  8'h64;        memory[27086] <=  8'h74;        memory[27087] <=  8'h75;        memory[27088] <=  8'h67;        memory[27089] <=  8'h79;        memory[27090] <=  8'h69;        memory[27091] <=  8'h68;        memory[27092] <=  8'h75;        memory[27093] <=  8'h6a;        memory[27094] <=  8'h6c;        memory[27095] <=  8'h62;        memory[27096] <=  8'h6d;        memory[27097] <=  8'h76;        memory[27098] <=  8'h6e;        memory[27099] <=  8'h63;        memory[27100] <=  8'h66;        memory[27101] <=  8'h68;        memory[27102] <=  8'h67;        memory[27103] <=  8'h79;        memory[27104] <=  8'h68;        memory[27105] <=  8'h75;        memory[27106] <=  8'h6a;        memory[27107] <=  8'h6e;        memory[27108] <=  8'h2c;        memory[27109] <=  8'h62;        memory[27110] <=  8'h6e;        memory[27111] <=  8'h6d;        memory[27112] <=  8'h76;        memory[27113] <=  8'h6e;        memory[27114] <=  8'h63;        memory[27115] <=  8'h66;        memory[27116] <=  8'h68;        memory[27117] <=  8'h74;        memory[27118] <=  8'h79;        memory[27119] <=  8'h69;        memory[27120] <=  8'h75;        memory[27121] <=  8'h6c;        memory[27122] <=  8'h6a;        memory[27123] <=  8'h62;        memory[27124] <=  8'h6d;        memory[27125] <=  8'h76;        memory[27126] <=  8'h6e;        memory[27127] <=  8'h63;        memory[27128] <=  8'h66;        memory[27129] <=  8'h74;        memory[27130] <=  8'h75;        memory[27131] <=  8'h79;        memory[27132] <=  8'h69;        memory[27133] <=  8'h68;        memory[27134] <=  8'h6b;        memory[27135] <=  8'h62;        memory[27136] <=  8'h76;        memory[27137] <=  8'h63;        memory[27138] <=  8'h66;        memory[27139] <=  8'h67;        memory[27140] <=  8'h74;        memory[27141] <=  8'h75;        memory[27142] <=  8'h79;        memory[27143] <=  8'h69;        memory[27144] <=  8'h75;        memory[27145] <=  8'h68;        memory[27146] <=  8'h6a;        memory[27147] <=  8'h6b;        memory[27148] <=  8'h62;        memory[27149] <=  8'h76;        memory[27150] <=  8'h63;        memory[27151] <=  8'h66;        memory[27152] <=  8'h74;        memory[27153] <=  8'h75;        memory[27154] <=  8'h79;        memory[27155] <=  8'h69;        memory[27156] <=  8'h75;        memory[27157] <=  8'h6a;        memory[27158] <=  8'h6b;        memory[27159] <=  8'h6e;        memory[27160] <=  8'h62;        memory[27161] <=  8'h76;        memory[27162] <=  8'h67;        memory[27163] <=  8'h66;        memory[27164] <=  8'h74;        memory[27165] <=  8'h79;        memory[27166] <=  8'h75;        memory[27167] <=  8'h75;        memory[27168] <=  8'h69;        memory[27169] <=  8'h6a;        memory[27170] <=  8'h6b;        memory[27171] <=  8'h68;        memory[27172] <=  8'h62;        memory[27173] <=  8'h6a;        memory[27174] <=  8'h67;        memory[27175] <=  8'h68;        memory[27176] <=  8'h66;        memory[27177] <=  8'h79;        memory[27178] <=  8'h74;        memory[27179] <=  8'h79;        memory[27180] <=  8'h69;        memory[27181] <=  8'h75;        memory[27182] <=  8'h64;        memory[27183] <=  8'h6a;        memory[27184] <=  8'h6b;        memory[27185] <=  8'h68;        memory[27186] <=  8'h63;        memory[27187] <=  8'h7a;        memory[27188] <=  8'h67;        memory[27189] <=  8'h68;        memory[27190] <=  8'h74;        memory[27191] <=  8'h75;        memory[27192] <=  8'h79;        memory[27193] <=  8'h69;        memory[27194] <=  8'h61;        memory[27195] <=  8'h73;        memory[27196] <=  8'h75;        memory[27197] <=  8'h6a;        memory[27198] <=  8'h6b;        memory[27199] <=  8'h62;        memory[27200] <=  8'h6e;        memory[27201] <=  8'h61;        memory[27202] <=  8'h76;        memory[27203] <=  8'h63;        memory[27204] <=  8'h66;        memory[27205] <=  8'h68;        memory[27206] <=  8'h75;        memory[27207] <=  8'h61;        memory[27208] <=  8'h73;        memory[27209] <=  8'h79;        memory[27210] <=  8'h64;        memory[27211] <=  8'h75;        memory[27212] <=  8'h69;        memory[27213] <=  8'h6a;        memory[27214] <=  8'h61;        memory[27215] <=  8'h6b;        memory[27216] <=  8'h62;        memory[27217] <=  8'h63;        memory[27218] <=  8'h78;        memory[27219] <=  8'h68;        memory[27220] <=  8'h67;        memory[27221] <=  8'h79;        memory[27222] <=  8'h75;        memory[27223] <=  8'h7a;        memory[27224] <=  8'h63;        memory[27225] <=  8'h61;        memory[27226] <=  8'h73;        memory[27227] <=  8'h69;        memory[27228] <=  8'h75;        memory[27229] <=  8'h6f;        memory[27230] <=  8'h69;        memory[27231] <=  8'h6a;        memory[27232] <=  8'h61;        memory[27233] <=  8'h6c;        memory[27234] <=  8'h63;        memory[27235] <=  8'h78;        memory[27236] <=  8'h62;        memory[27237] <=  8'h63;        memory[27238] <=  8'h20;        memory[27239] <=  8'h6e;        memory[27240] <=  8'h76;        memory[27241] <=  8'h63;        memory[27242] <=  8'h61;        memory[27243] <=  8'h64;        memory[27244] <=  8'h73;        memory[27245] <=  8'h67;        memory[27246] <=  8'h79;        memory[27247] <=  8'h68;        memory[27248] <=  8'h75;        memory[27249] <=  8'h61;        memory[27250] <=  8'h6a;        memory[27251] <=  8'h6b;        memory[27252] <=  8'h78;        memory[27253] <=  8'h62;        memory[27254] <=  8'h20;        memory[27255] <=  8'h6e;        memory[27256] <=  8'h76;        memory[27257] <=  8'h63;        memory[27258] <=  8'h61;        memory[27259] <=  8'h73;        memory[27260] <=  8'h67;        memory[27261] <=  8'h68;        memory[27262] <=  8'h75;        memory[27263] <=  8'h6a;        memory[27264] <=  8'h6c;        memory[27265] <=  8'h6b;        memory[27266] <=  8'h63;        memory[27267] <=  8'h78;        memory[27268] <=  8'h20;        memory[27269] <=  8'h6a;        memory[27270] <=  8'h6b;        memory[27271] <=  8'h68;        memory[27272] <=  8'h61;        memory[27273] <=  8'h73;        memory[27274] <=  8'h76;        memory[27275] <=  8'h64;        memory[27276] <=  8'h6e;        memory[27277] <=  8'h20;        memory[27278] <=  8'h62;        memory[27279] <=  8'h6e;        memory[27280] <=  8'h6d;        memory[27281] <=  8'h6b;        memory[27282] <=  8'h77;        memory[27283] <=  8'h64;        memory[27284] <=  8'h6f;        memory[27285] <=  8'h77;        memory[27286] <=  8'h69;        memory[27287] <=  8'h6f;        memory[27288] <=  8'h75;        memory[27289] <=  8'h69;        memory[27290] <=  8'h68;        memory[27291] <=  8'h62;        memory[27292] <=  8'h6e;        memory[27293] <=  8'h6b;        memory[27294] <=  8'h77;        memory[27295] <=  8'h69;        memory[27296] <=  8'h6f;        memory[27297] <=  8'h75;        memory[27298] <=  8'h71;        memory[27299] <=  8'h69;        memory[27300] <=  8'h79;        memory[27301] <=  8'h67;        memory[27302] <=  8'h6a;        memory[27303] <=  8'h64;        memory[27304] <=  8'h61;        memory[27305] <=  8'h76;        memory[27306] <=  8'h62;        memory[27307] <=  8'h6e;        memory[27308] <=  8'h6b;        memory[27309] <=  8'h6f;        memory[27310] <=  8'h70;        memory[27311] <=  8'h64;        memory[27312] <=  8'h76;        memory[27313] <=  8'h69;        memory[27314] <=  8'h6f;        memory[27315] <=  8'h75;        memory[27316] <=  8'h69;        memory[27317] <=  8'h48;        memory[27318] <=  8'h42;        memory[27319] <=  8'h6b;        memory[27320] <=  8'h64;        memory[27321] <=  8'h6e;        memory[27322] <=  8'h6c;        memory[27323] <=  8'h71;        memory[27324] <=  8'h6b;        memory[27325] <=  8'h6d;        memory[27326] <=  8'h6a;        memory[27327] <=  8'h70;        memory[27328] <=  8'h69;        memory[27329] <=  8'h6f;        memory[27330] <=  8'h68;        memory[27331] <=  8'h65;        memory[27332] <=  8'h66;        memory[27333] <=  8'h75;        memory[27334] <=  8'h67;        memory[27335] <=  8'h69;        memory[27336] <=  8'h73;        memory[27337] <=  8'h61;        memory[27338] <=  8'h62;        memory[27339] <=  8'h64;        memory[27340] <=  8'h6b;        memory[27341] <=  8'h6a;        memory[27342] <=  8'h6b;        memory[27343] <=  8'h6c;        memory[27344] <=  8'h6a;        memory[27345] <=  8'h69;        memory[27346] <=  8'h73;        memory[27347] <=  8'h6f;        memory[27348] <=  8'h71;        memory[27349] <=  8'h68;        memory[27350] <=  8'h77;        memory[27351] <=  8'h67;        memory[27352] <=  8'h69;        memory[27353] <=  8'h79;        memory[27354] <=  8'h6a;        memory[27355] <=  8'h64;        memory[27356] <=  8'h76;        memory[27357] <=  8'h62;        memory[27358] <=  8'h6e;        memory[27359] <=  8'h61;        memory[27360] <=  8'h73;        memory[27361] <=  8'h66;        memory[27362] <=  8'h6c;        memory[27363] <=  8'h6b;        memory[27364] <=  8'h64;        memory[27365] <=  8'h6a;        memory[27366] <=  8'h68;        memory[27367] <=  8'h63;        memory[27368] <=  8'h67;        memory[27369] <=  8'h6a;        memory[27370] <=  8'h76;        memory[27371] <=  8'h73;        memory[27372] <=  8'h64;        memory[27373] <=  8'h62;        memory[27374] <=  8'h62;        memory[27375] <=  8'h61;        memory[27376] <=  8'h72;        memory[27377] <=  8'h62;        memory[27378] <=  8'h62;        memory[27379] <=  8'h73;        memory[27380] <=  8'h62;        memory[27381] <=  8'h67;        memory[27382] <=  8'h73;        memory[27383] <=  8'h66;        memory[27384] <=  8'h67;        memory[27385] <=  8'h61;        memory[27386] <=  8'h68;        memory[27387] <=  8'h66;        memory[27388] <=  8'h73;        memory[27389] <=  8'h68;        memory[27390] <=  8'h61;        memory[27391] <=  8'h66;        memory[27392] <=  8'h73;        memory[27393] <=  8'h66;        memory[27394] <=  8'h68;        memory[27395] <=  8'h61;        memory[27396] <=  8'h69;        memory[27397] <=  8'h64;        memory[27398] <=  8'h75;        memory[27399] <=  8'h67;        memory[27400] <=  8'h64;        memory[27401] <=  8'h77;        memory[27402] <=  8'h62;        memory[27403] <=  8'h61;        memory[27404] <=  8'h62;        memory[27405] <=  8'h72;        memory[27406] <=  8'h62;        memory[27407] <=  8'h61;        memory[27408] <=  8'h62;        memory[27409] <=  8'h62;        memory[27410] <=  8'h74;        memory[27411] <=  8'h62;        memory[27412] <=  8'h62;        memory[27413] <=  8'h62;        memory[27414] <=  8'h62;        memory[27415] <=  8'h62;        memory[27416] <=  8'h62;        memory[27417] <=  8'h62;        memory[27418] <=  8'h62;        memory[27419] <=  8'h61;        memory[27420] <=  8'h62;        memory[27421] <=  8'h62;        memory[27422] <=  8'h72;        memory[27423] <=  8'h74;        memory[27424] <=  8'h62;        memory[27425] <=  8'h62;        memory[27426] <=  8'h61;        memory[27427] <=  8'h62;        memory[27428] <=  8'h72;        memory[27429] <=  8'h62;        memory[27430] <=  8'h74;        memory[27431] <=  8'h62;        memory[27432] <=  8'h62;        memory[27433] <=  8'h62;        memory[27434] <=  8'h63;        memory[27435] <=  8'h61;        memory[27436] <=  8'h72;        memory[27437] <=  8'h74;        memory[27438] <=  8'h73;        memory[27439] <=  8'h62;        memory[27440] <=  8'h61;        memory[27441] <=  8'h72;        memory[27442] <=  8'h74;        memory[27443] <=  8'h74;        memory[27444] <=  8'h62;        memory[27445] <=  8'h61;        memory[27446] <=  8'h72;        memory[27447] <=  8'h74;        memory[27448] <=  8'h78;        memory[27449] <=  8'h61;        memory[27450] <=  8'h74;        memory[27451] <=  8'h6b;        memory[27452] <=  8'h73;        memory[27453] <=  8'h68;        memory[27454] <=  8'h63;        memory[27455] <=  8'h66;        memory[27456] <=  8'h69;        memory[27457] <=  8'h77;        memory[27458] <=  8'h68;        memory[27459] <=  8'h61;        memory[27460] <=  8'h74;        memory[27461] <=  8'h61;        memory[27462] <=  8'h6e;        memory[27463] <=  8'h61;        memory[27464] <=  8'h62;        memory[27465] <=  8'h61;        memory[27466] <=  8'h63;        memory[27467] <=  8'h61;        memory[27468] <=  8'h74;        memory[27469] <=  8'h61;        memory[27470] <=  8'h62;        memory[27471] <=  8'h61;        memory[27472] <=  8'h72;        memory[27473] <=  8'h63;        memory[27474] <=  8'h61;        memory[27475] <=  8'h68;        memory[27476] <=  8'h64;        memory[27477] <=  8'h75;        memory[27478] <=  8'h63;        memory[27479] <=  8'h74;        memory[27480] <=  8'h61;        memory[27481] <=  8'h64;        memory[27482] <=  8'h61;        memory[27483] <=  8'h61;        memory[27484] <=  8'h63;        memory[27485] <=  8'h61;        memory[27486] <=  8'h72;        memory[27487] <=  8'h63;        memory[27488] <=  8'h74;        memory[27489] <=  8'h72;        memory[27490] <=  8'h63;        memory[27491] <=  8'h61;        memory[27492] <=  8'h74;        memory[27493] <=  8'h72;        memory[27494] <=  8'h63;        memory[27495] <=  8'h61;        memory[27496] <=  8'h74;        memory[27497] <=  8'h63;        memory[27498] <=  8'h62;        memory[27499] <=  8'h61;        memory[27500] <=  8'h74;        memory[27501] <=  8'h62;        memory[27502] <=  8'h72;        memory[27503] <=  8'h63;        memory[27504] <=  8'h61;        memory[27505] <=  8'h74;        memory[27506] <=  8'h72;        memory[27507] <=  8'h6e;        memory[27508] <=  8'h62;        memory[27509] <=  8'h61;        memory[27510] <=  8'h63;        memory[27511] <=  8'h61;        memory[27512] <=  8'h74;        memory[27513] <=  8'h79;        memory[27514] <=  8'h73;        memory[27515] <=  8'h6e;        memory[27516] <=  8'h63;        memory[27517] <=  8'h74;        memory[27518] <=  8'h61;        memory[27519] <=  8'h6e;        memory[27520] <=  8'h62;        memory[27521] <=  8'h61;        memory[27522] <=  8'h63;        memory[27523] <=  8'h72;        memory[27524] <=  8'h6e;        memory[27525] <=  8'h74;        memory[27526] <=  8'h61;        memory[27527] <=  8'h62;        memory[27528] <=  8'h74;        memory[27529] <=  8'h6e;        memory[27530] <=  8'h61;        memory[27531] <=  8'h72;        memory[27532] <=  8'h62;        memory[27533] <=  8'h78;        memory[27534] <=  8'h74;        memory[27535] <=  8'h61;        memory[27536] <=  8'h72;        memory[27537] <=  8'h62;        memory[27538] <=  8'h61;        memory[27539] <=  8'h72;        memory[27540] <=  8'h74;        memory[27541] <=  8'h74;        memory[27542] <=  8'h62;        memory[27543] <=  8'h61;        memory[27544] <=  8'h72;        memory[27545] <=  8'h74;        memory[27546] <=  8'h78;        memory[27547] <=  8'h61;        memory[27548] <=  8'h74;        memory[27549] <=  8'h6b;        memory[27550] <=  8'h73;        memory[27551] <=  8'h68;        memory[27552] <=  8'h63;        memory[27553] <=  8'h66;        memory[27554] <=  8'h69;        memory[27555] <=  8'h77;        memory[27556] <=  8'h68;        memory[27557] <=  8'h61;        memory[27558] <=  8'h74;        memory[27559] <=  8'h61;        memory[27560] <=  8'h6e;        memory[27561] <=  8'h61;        memory[27562] <=  8'h62;        memory[27563] <=  8'h61;        memory[27564] <=  8'h63;        memory[27565] <=  8'h61;        memory[27566] <=  8'h74;        memory[27567] <=  8'h61;        memory[27568] <=  8'h62;        memory[27569] <=  8'h61;        memory[27570] <=  8'h72;        memory[27571] <=  8'h63;        memory[27572] <=  8'h61;        memory[27573] <=  8'h68;        memory[27574] <=  8'h64;        memory[27575] <=  8'h75;        memory[27576] <=  8'h63;        memory[27577] <=  8'h74;        memory[27578] <=  8'h61;        memory[27579] <=  8'h64;        memory[27580] <=  8'h61;        memory[27581] <=  8'h61;        memory[27582] <=  8'h63;        memory[27583] <=  8'h61;        memory[27584] <=  8'h72;        memory[27585] <=  8'h63;        memory[27586] <=  8'h74;        memory[27587] <=  8'h72;        memory[27588] <=  8'h63;        memory[27589] <=  8'h61;        memory[27590] <=  8'h74;        memory[27591] <=  8'h72;        memory[27592] <=  8'h63;        memory[27593] <=  8'h61;        memory[27594] <=  8'h74;        memory[27595] <=  8'h63;        memory[27596] <=  8'h62;        memory[27597] <=  8'h61;        memory[27598] <=  8'h74;        memory[27599] <=  8'h62;        memory[27600] <=  8'h72;        memory[27601] <=  8'h63;        memory[27602] <=  8'h61;        memory[27603] <=  8'h74;        memory[27604] <=  8'h72;        memory[27605] <=  8'h6e;        memory[27606] <=  8'h62;        memory[27607] <=  8'h61;        memory[27608] <=  8'h63;        memory[27609] <=  8'h61;        memory[27610] <=  8'h74;        memory[27611] <=  8'h79;        memory[27612] <=  8'h73;        memory[27613] <=  8'h6e;        memory[27614] <=  8'h63;        memory[27615] <=  8'h74;        memory[27616] <=  8'h61;        memory[27617] <=  8'h6e;        memory[27618] <=  8'h62;        memory[27619] <=  8'h61;        memory[27620] <=  8'h63;        memory[27621] <=  8'h72;        memory[27622] <=  8'h6e;        memory[27623] <=  8'h74;        memory[27624] <=  8'h61;        memory[27625] <=  8'h62;        memory[27626] <=  8'h74;        memory[27627] <=  8'h6e;        memory[27628] <=  8'h61;        memory[27629] <=  8'h72;        memory[27630] <=  8'h62;        memory[27631] <=  8'h78;        memory[27632] <=  8'h74;        memory[27633] <=  8'h61;        memory[27634] <=  8'h72;        memory[27635] <=  8'h62;        memory[27636] <=  8'h61;        memory[27637] <=  8'h72;        memory[27638] <=  8'h74;        memory[27639] <=  8'h74;        memory[27640] <=  8'h62;        memory[27641] <=  8'h61;        memory[27642] <=  8'h72;        memory[27643] <=  8'h74;        memory[27644] <=  8'h78;        memory[27645] <=  8'h61;        memory[27646] <=  8'h74;        memory[27647] <=  8'h6b;        memory[27648] <=  8'h73;        memory[27649] <=  8'h68;        memory[27650] <=  8'h63;        memory[27651] <=  8'h66;        memory[27652] <=  8'h69;        memory[27653] <=  8'h77;        memory[27654] <=  8'h68;        memory[27655] <=  8'h61;        memory[27656] <=  8'h74;        memory[27657] <=  8'h61;        memory[27658] <=  8'h6e;        memory[27659] <=  8'h61;        memory[27660] <=  8'h62;        memory[27661] <=  8'h61;        memory[27662] <=  8'h63;        memory[27663] <=  8'h61;        memory[27664] <=  8'h74;        memory[27665] <=  8'h61;        memory[27666] <=  8'h62;        memory[27667] <=  8'h61;        memory[27668] <=  8'h72;        memory[27669] <=  8'h63;        memory[27670] <=  8'h61;        memory[27671] <=  8'h68;        memory[27672] <=  8'h64;        memory[27673] <=  8'h75;        memory[27674] <=  8'h63;        memory[27675] <=  8'h74;        memory[27676] <=  8'h61;        memory[27677] <=  8'h64;        memory[27678] <=  8'h61;        memory[27679] <=  8'h61;        memory[27680] <=  8'h63;        memory[27681] <=  8'h61;        memory[27682] <=  8'h72;        memory[27683] <=  8'h63;        memory[27684] <=  8'h74;        memory[27685] <=  8'h72;        memory[27686] <=  8'h63;        memory[27687] <=  8'h61;        memory[27688] <=  8'h74;        memory[27689] <=  8'h72;        memory[27690] <=  8'h63;        memory[27691] <=  8'h61;        memory[27692] <=  8'h74;        memory[27693] <=  8'h63;        memory[27694] <=  8'h62;        memory[27695] <=  8'h61;        memory[27696] <=  8'h74;        memory[27697] <=  8'h62;        memory[27698] <=  8'h72;        memory[27699] <=  8'h63;        memory[27700] <=  8'h61;        memory[27701] <=  8'h74;        memory[27702] <=  8'h72;        memory[27703] <=  8'h6e;        memory[27704] <=  8'h62;        memory[27705] <=  8'h61;        memory[27706] <=  8'h63;        memory[27707] <=  8'h61;        memory[27708] <=  8'h74;        memory[27709] <=  8'h79;        memory[27710] <=  8'h73;        memory[27711] <=  8'h6e;        memory[27712] <=  8'h63;        memory[27713] <=  8'h74;        memory[27714] <=  8'h61;        memory[27715] <=  8'h6e;        memory[27716] <=  8'h62;        memory[27717] <=  8'h61;        memory[27718] <=  8'h63;        memory[27719] <=  8'h72;        memory[27720] <=  8'h6e;        memory[27721] <=  8'h74;        memory[27722] <=  8'h61;        memory[27723] <=  8'h62;        memory[27724] <=  8'h74;        memory[27725] <=  8'h6e;        memory[27726] <=  8'h61;        memory[27727] <=  8'h72;        memory[27728] <=  8'h62;        memory[27729] <=  8'h78;        memory[27730] <=  8'h74;        memory[27731] <=  8'h61;        memory[27732] <=  8'h72;        memory[27733] <=  8'h5d;        memory[27734] <=  8'h5d;        memory[27735] <=  8'h65;        memory[27736] <=  8'h66;        memory[27737] <=  8'h77;        memory[27738] <=  8'h65;        memory[27739] <=  8'h5d;        memory[27740] <=  8'h65;        memory[27741] <=  8'h67;        memory[27742] <=  8'h73;        memory[27743] <=  8'h67;        memory[27744] <=  8'h66;        memory[27745] <=  8'h62;        memory[27746] <=  8'h61;        memory[27747] <=  8'h72;        memory[27748] <=  8'h74;        memory[27749] <=  8'h74;        memory[27750] <=  8'h62;        memory[27751] <=  8'h61;        memory[27752] <=  8'h72;        memory[27753] <=  8'h74;        memory[27754] <=  8'h78;        memory[27755] <=  8'h61;        memory[27756] <=  8'h74;        memory[27757] <=  8'h6b;        memory[27758] <=  8'h73;        memory[27759] <=  8'h68;        memory[27760] <=  8'h63;        memory[27761] <=  8'h66;        memory[27762] <=  8'h69;        memory[27763] <=  8'h77;        memory[27764] <=  8'h68;        memory[27765] <=  8'h61;        memory[27766] <=  8'h74;        memory[27767] <=  8'h61;        memory[27768] <=  8'h6e;        memory[27769] <=  8'h61;        memory[27770] <=  8'h62;        memory[27771] <=  8'h61;        memory[27772] <=  8'h63;        memory[27773] <=  8'h61;        memory[27774] <=  8'h74;        memory[27775] <=  8'h61;        memory[27776] <=  8'h62;        memory[27777] <=  8'h61;        memory[27778] <=  8'h72;        memory[27779] <=  8'h63;        memory[27780] <=  8'h61;        memory[27781] <=  8'h68;        memory[27782] <=  8'h64;        memory[27783] <=  8'h75;        memory[27784] <=  8'h63;        memory[27785] <=  8'h74;        memory[27786] <=  8'h61;        memory[27787] <=  8'h64;        memory[27788] <=  8'h61;        memory[27789] <=  8'h61;        memory[27790] <=  8'h63;        memory[27791] <=  8'h61;        memory[27792] <=  8'h72;        memory[27793] <=  8'h63;        memory[27794] <=  8'h74;        memory[27795] <=  8'h72;        memory[27796] <=  8'h63;        memory[27797] <=  8'h61;        memory[27798] <=  8'h74;        memory[27799] <=  8'h72;        memory[27800] <=  8'h63;        memory[27801] <=  8'h61;        memory[27802] <=  8'h74;        memory[27803] <=  8'h63;        memory[27804] <=  8'h62;        memory[27805] <=  8'h61;        memory[27806] <=  8'h74;        memory[27807] <=  8'h62;        memory[27808] <=  8'h72;        memory[27809] <=  8'h63;        memory[27810] <=  8'h61;        memory[27811] <=  8'h74;        memory[27812] <=  8'h72;        memory[27813] <=  8'h6e;        memory[27814] <=  8'h62;        memory[27815] <=  8'h61;        memory[27816] <=  8'h63;        memory[27817] <=  8'h61;        memory[27818] <=  8'h74;        memory[27819] <=  8'h79;        memory[27820] <=  8'h73;        memory[27821] <=  8'h6e;        memory[27822] <=  8'h63;        memory[27823] <=  8'h74;        memory[27824] <=  8'h61;        memory[27825] <=  8'h6e;        memory[27826] <=  8'h62;        memory[27827] <=  8'h61;        memory[27828] <=  8'h63;        memory[27829] <=  8'h72;        memory[27830] <=  8'h6e;        memory[27831] <=  8'h74;        memory[27832] <=  8'h61;        memory[27833] <=  8'h62;        memory[27834] <=  8'h74;        memory[27835] <=  8'h6e;        memory[27836] <=  8'h61;        memory[27837] <=  8'h72;        memory[27838] <=  8'h62;        memory[27839] <=  8'h78;        memory[27840] <=  8'h74;        memory[27841] <=  8'h61;        memory[27842] <=  8'h72;        memory[27843] <=  8'h62;        memory[27844] <=  8'h61;        memory[27845] <=  8'h72;        memory[27846] <=  8'h74;        memory[27847] <=  8'h74;        memory[27848] <=  8'h62;        memory[27849] <=  8'h61;        memory[27850] <=  8'h72;        memory[27851] <=  8'h74;        memory[27852] <=  8'h78;        memory[27853] <=  8'h61;        memory[27854] <=  8'h74;        memory[27855] <=  8'h6b;        memory[27856] <=  8'h73;        memory[27857] <=  8'h68;        memory[27858] <=  8'h63;        memory[27859] <=  8'h66;        memory[27860] <=  8'h69;        memory[27861] <=  8'h77;        memory[27862] <=  8'h68;        memory[27863] <=  8'h61;        memory[27864] <=  8'h74;        memory[27865] <=  8'h61;        memory[27866] <=  8'h6e;        memory[27867] <=  8'h61;        memory[27868] <=  8'h62;        memory[27869] <=  8'h61;        memory[27870] <=  8'h63;        memory[27871] <=  8'h61;        memory[27872] <=  8'h74;        memory[27873] <=  8'h61;        memory[27874] <=  8'h62;        memory[27875] <=  8'h61;        memory[27876] <=  8'h72;        memory[27877] <=  8'h63;        memory[27878] <=  8'h61;        memory[27879] <=  8'h68;        memory[27880] <=  8'h64;        memory[27881] <=  8'h75;        memory[27882] <=  8'h63;        memory[27883] <=  8'h74;        memory[27884] <=  8'h61;        memory[27885] <=  8'h64;        memory[27886] <=  8'h61;        memory[27887] <=  8'h61;        memory[27888] <=  8'h63;        memory[27889] <=  8'h61;        memory[27890] <=  8'h72;        memory[27891] <=  8'h63;        memory[27892] <=  8'h74;        memory[27893] <=  8'h72;        memory[27894] <=  8'h63;        memory[27895] <=  8'h61;        memory[27896] <=  8'h74;        memory[27897] <=  8'h72;        memory[27898] <=  8'h63;        memory[27899] <=  8'h61;        memory[27900] <=  8'h74;        memory[27901] <=  8'h63;        memory[27902] <=  8'h62;        memory[27903] <=  8'h61;        memory[27904] <=  8'h74;        memory[27905] <=  8'h62;        memory[27906] <=  8'h72;        memory[27907] <=  8'h63;        memory[27908] <=  8'h61;        memory[27909] <=  8'h74;        memory[27910] <=  8'h72;        memory[27911] <=  8'h6e;        memory[27912] <=  8'h62;        memory[27913] <=  8'h61;        memory[27914] <=  8'h63;        memory[27915] <=  8'h61;        memory[27916] <=  8'h74;        memory[27917] <=  8'h79;        memory[27918] <=  8'h73;        memory[27919] <=  8'h6e;        memory[27920] <=  8'h63;        memory[27921] <=  8'h74;        memory[27922] <=  8'h61;        memory[27923] <=  8'h6e;        memory[27924] <=  8'h62;        memory[27925] <=  8'h61;        memory[27926] <=  8'h63;        memory[27927] <=  8'h72;        memory[27928] <=  8'h6e;        memory[27929] <=  8'h74;        memory[27930] <=  8'h61;        memory[27931] <=  8'h62;        memory[27932] <=  8'h74;        memory[27933] <=  8'h6e;        memory[27934] <=  8'h61;        memory[27935] <=  8'h72;        memory[27936] <=  8'h62;        memory[27937] <=  8'h78;        memory[27938] <=  8'h74;        memory[27939] <=  8'h61;        memory[27940] <=  8'h72;        memory[27941] <=  8'h64;        memory[27942] <=  8'h66;        memory[27943] <=  8'h73;        memory[27944] <=  8'h67;        memory[27945] <=  8'h76;        memory[27946] <=  8'h68;        memory[27947] <=  8'h62;        memory[27948] <=  8'h6b;        memory[27949] <=  8'h6a;        memory[27950] <=  8'h6e;        memory[27951] <=  8'h6d;        memory[27952] <=  8'h62;        memory[27953] <=  8'h76;        memory[27954] <=  8'h78;        memory[27955] <=  8'h63;        memory[27956] <=  8'h73;        memory[27957] <=  8'h66;        memory[27958] <=  8'h72;        memory[27959] <=  8'h74;        memory[27960] <=  8'h79;        memory[27961] <=  8'h75;        memory[27962] <=  8'h6a;        memory[27963] <=  8'h6e;        memory[27964] <=  8'h62;        memory[27965] <=  8'h76;        memory[27966] <=  8'h63;        memory[27967] <=  8'h64;        memory[27968] <=  8'h74;        memory[27969] <=  8'h79;        memory[27970] <=  8'h75;        memory[27971] <=  8'h69;        memory[27972] <=  8'h6b;        memory[27973] <=  8'h6d;        memory[27974] <=  8'h6e;        memory[27975] <=  8'h62;        memory[27976] <=  8'h76;        memory[27977] <=  8'h63;        memory[27978] <=  8'h78;        memory[27979] <=  8'h73;        memory[27980] <=  8'h64;        memory[27981] <=  8'h72;        memory[27982] <=  8'h74;        memory[27983] <=  8'h79;        memory[27984] <=  8'h75;        memory[27985] <=  8'h69;        memory[27986] <=  8'h6b;        memory[27987] <=  8'h6d;        memory[27988] <=  8'h6e;        memory[27989] <=  8'h62;        memory[27990] <=  8'h76;        memory[27991] <=  8'h63;        memory[27992] <=  8'h73;        memory[27993] <=  8'h77;        memory[27994] <=  8'h33;        memory[27995] <=  8'h34;        memory[27996] <=  8'h35;        memory[27997] <=  8'h36;        memory[27998] <=  8'h37;        memory[27999] <=  8'h38;        memory[28000] <=  8'h69;        memory[28001] <=  8'h6b;        memory[28002] <=  8'h6d;        memory[28003] <=  8'h6e;        memory[28004] <=  8'h62;        memory[28005] <=  8'h76;        memory[28006] <=  8'h63;        memory[28007] <=  8'h64;        memory[28008] <=  8'h65;        memory[28009] <=  8'h72;        memory[28010] <=  8'h36;        memory[28011] <=  8'h37;        memory[28012] <=  8'h38;        memory[28013] <=  8'h69;        memory[28014] <=  8'h6f;        memory[28015] <=  8'h6b;        memory[28016] <=  8'h6a;        memory[28017] <=  8'h6e;        memory[28018] <=  8'h62;        memory[28019] <=  8'h76;        memory[28020] <=  8'h63;        memory[28021] <=  8'h64;        memory[28022] <=  8'h72;        memory[28023] <=  8'h74;        memory[28024] <=  8'h79;        memory[28025] <=  8'h75;        memory[28026] <=  8'h73;        memory[28027] <=  8'h6a;        memory[28028] <=  8'h63;        memory[28029] <=  8'h6e;        memory[28030] <=  8'h62;        memory[28031] <=  8'h64;        memory[28032] <=  8'h66;        memory[28033] <=  8'h73;        memory[28034] <=  8'h74;        memory[28035] <=  8'h79;        memory[28036] <=  8'h75;        memory[28037] <=  8'h61;        memory[28038] <=  8'h69;        memory[28039] <=  8'h6b;        memory[28040] <=  8'h78;        memory[28041] <=  8'h6d;        memory[28042] <=  8'h6e;        memory[28043] <=  8'h73;        memory[28044] <=  8'h6a;        memory[28045] <=  8'h6f;        memory[28046] <=  8'h64;        memory[28047] <=  8'h6c;        memory[28048] <=  8'h63;        memory[28049] <=  8'h78;        memory[28050] <=  8'h62;        memory[28051] <=  8'h61;        memory[28052] <=  8'h72;        memory[28053] <=  8'h74;        memory[28054] <=  8'h78;        memory[28055] <=  8'h61;        memory[28056] <=  8'h74;        memory[28057] <=  8'h6b;        memory[28058] <=  8'h73;        memory[28059] <=  8'h68;        memory[28060] <=  8'h63;        memory[28061] <=  8'h66;        memory[28062] <=  8'h69;        memory[28063] <=  8'h77;        memory[28064] <=  8'h68;        memory[28065] <=  8'h61;        memory[28066] <=  8'h74;        memory[28067] <=  8'h61;        memory[28068] <=  8'h6e;        memory[28069] <=  8'h61;        memory[28070] <=  8'h62;        memory[28071] <=  8'h61;        memory[28072] <=  8'h63;        memory[28073] <=  8'h61;        memory[28074] <=  8'h74;        memory[28075] <=  8'h61;        memory[28076] <=  8'h62;        memory[28077] <=  8'h61;        memory[28078] <=  8'h72;        memory[28079] <=  8'h63;        memory[28080] <=  8'h61;        memory[28081] <=  8'h68;        memory[28082] <=  8'h64;        memory[28083] <=  8'h75;        memory[28084] <=  8'h63;        memory[28085] <=  8'h74;        memory[28086] <=  8'h61;        memory[28087] <=  8'h64;        memory[28088] <=  8'h61;        memory[28089] <=  8'h61;        memory[28090] <=  8'h63;        memory[28091] <=  8'h61;        memory[28092] <=  8'h72;        memory[28093] <=  8'h62;        memory[28094] <=  8'h61;        memory[28095] <=  8'h72;        memory[28096] <=  8'h74;        memory[28097] <=  8'h78;        memory[28098] <=  8'h61;        memory[28099] <=  8'h74;        memory[28100] <=  8'h6b;        memory[28101] <=  8'h73;        memory[28102] <=  8'h68;        memory[28103] <=  8'h63;        memory[28104] <=  8'h66;        memory[28105] <=  8'h69;        memory[28106] <=  8'h77;        memory[28107] <=  8'h68;        memory[28108] <=  8'h61;        memory[28109] <=  8'h74;        memory[28110] <=  8'h61;        memory[28111] <=  8'h6e;        memory[28112] <=  8'h61;        memory[28113] <=  8'h62;        memory[28114] <=  8'h61;        memory[28115] <=  8'h63;        memory[28116] <=  8'h61;        memory[28117] <=  8'h74;        memory[28118] <=  8'h61;        memory[28119] <=  8'h62;        memory[28120] <=  8'h61;        memory[28121] <=  8'h72;        memory[28122] <=  8'h63;        memory[28123] <=  8'h61;        memory[28124] <=  8'h68;        memory[28125] <=  8'h64;        memory[28126] <=  8'h75;        memory[28127] <=  8'h63;        memory[28128] <=  8'h74;        memory[28129] <=  8'h61;        memory[28130] <=  8'h64;        memory[28131] <=  8'h61;        memory[28132] <=  8'h61;        memory[28133] <=  8'h63;        memory[28134] <=  8'h61;        memory[28135] <=  8'h72;        memory[28136] <=  8'h62;        memory[28137] <=  8'h61;        memory[28138] <=  8'h72;        memory[28139] <=  8'h74;        memory[28140] <=  8'h78;        memory[28141] <=  8'h61;        memory[28142] <=  8'h74;        memory[28143] <=  8'h6b;        memory[28144] <=  8'h73;        memory[28145] <=  8'h68;        memory[28146] <=  8'h63;        memory[28147] <=  8'h66;        memory[28148] <=  8'h69;        memory[28149] <=  8'h77;        memory[28150] <=  8'h68;        memory[28151] <=  8'h61;        memory[28152] <=  8'h74;        memory[28153] <=  8'h61;        memory[28154] <=  8'h6e;        memory[28155] <=  8'h61;        memory[28156] <=  8'h62;        memory[28157] <=  8'h61;        memory[28158] <=  8'h63;        memory[28159] <=  8'h61;        memory[28160] <=  8'h74;        memory[28161] <=  8'h61;        memory[28162] <=  8'h62;        memory[28163] <=  8'h61;        memory[28164] <=  8'h72;        memory[28165] <=  8'h63;        memory[28166] <=  8'h61;        memory[28167] <=  8'h68;        memory[28168] <=  8'h64;        memory[28169] <=  8'h75;        memory[28170] <=  8'h63;        memory[28171] <=  8'h74;        memory[28172] <=  8'h61;        memory[28173] <=  8'h64;        memory[28174] <=  8'h61;        memory[28175] <=  8'h61;        memory[28176] <=  8'h63;        memory[28177] <=  8'h61;        memory[28178] <=  8'h72;        memory[28179] <=  8'h62;        memory[28180] <=  8'h61;        memory[28181] <=  8'h72;        memory[28182] <=  8'h74;        memory[28183] <=  8'h78;        memory[28184] <=  8'h61;        memory[28185] <=  8'h74;        memory[28186] <=  8'h6b;        memory[28187] <=  8'h73;        memory[28188] <=  8'h68;        memory[28189] <=  8'h63;        memory[28190] <=  8'h66;        memory[28191] <=  8'h69;        memory[28192] <=  8'h77;        memory[28193] <=  8'h68;        memory[28194] <=  8'h61;        memory[28195] <=  8'h74;        memory[28196] <=  8'h61;        memory[28197] <=  8'h6e;        memory[28198] <=  8'h61;        memory[28199] <=  8'h62;        memory[28200] <=  8'h61;        memory[28201] <=  8'h63;        memory[28202] <=  8'h61;        memory[28203] <=  8'h74;        memory[28204] <=  8'h61;        memory[28205] <=  8'h62;        memory[28206] <=  8'h61;        memory[28207] <=  8'h72;        memory[28208] <=  8'h63;        memory[28209] <=  8'h61;        memory[28210] <=  8'h68;        memory[28211] <=  8'h64;        memory[28212] <=  8'h75;        memory[28213] <=  8'h63;        memory[28214] <=  8'h74;        memory[28215] <=  8'h61;        memory[28216] <=  8'h64;        memory[28217] <=  8'h61;        memory[28218] <=  8'h61;        memory[28219] <=  8'h63;        memory[28220] <=  8'h61;        memory[28221] <=  8'h72;        memory[28222] <=  8'h62;        memory[28223] <=  8'h61;        memory[28224] <=  8'h72;        memory[28225] <=  8'h74;        memory[28226] <=  8'h78;        memory[28227] <=  8'h61;        memory[28228] <=  8'h74;        memory[28229] <=  8'h6b;        memory[28230] <=  8'h73;        memory[28231] <=  8'h68;        memory[28232] <=  8'h63;        memory[28233] <=  8'h66;        memory[28234] <=  8'h69;        memory[28235] <=  8'h77;        memory[28236] <=  8'h68;        memory[28237] <=  8'h61;        memory[28238] <=  8'h74;        memory[28239] <=  8'h61;        memory[28240] <=  8'h6e;        memory[28241] <=  8'h61;        memory[28242] <=  8'h62;        memory[28243] <=  8'h61;        memory[28244] <=  8'h63;        memory[28245] <=  8'h61;        memory[28246] <=  8'h74;        memory[28247] <=  8'h61;        memory[28248] <=  8'h62;        memory[28249] <=  8'h61;        memory[28250] <=  8'h72;        memory[28251] <=  8'h63;        memory[28252] <=  8'h61;        memory[28253] <=  8'h68;        memory[28254] <=  8'h64;        memory[28255] <=  8'h75;        memory[28256] <=  8'h63;        memory[28257] <=  8'h74;        memory[28258] <=  8'h61;        memory[28259] <=  8'h64;        memory[28260] <=  8'h61;        memory[28261] <=  8'h61;        memory[28262] <=  8'h63;        memory[28263] <=  8'h61;        memory[28264] <=  8'h72;        memory[28265] <=  8'h62;        memory[28266] <=  8'h61;        memory[28267] <=  8'h72;        memory[28268] <=  8'h74;        memory[28269] <=  8'h78;        memory[28270] <=  8'h61;        memory[28271] <=  8'h74;        memory[28272] <=  8'h6b;        memory[28273] <=  8'h73;        memory[28274] <=  8'h68;        memory[28275] <=  8'h63;        memory[28276] <=  8'h66;        memory[28277] <=  8'h69;        memory[28278] <=  8'h77;        memory[28279] <=  8'h68;        memory[28280] <=  8'h61;        memory[28281] <=  8'h74;        memory[28282] <=  8'h61;        memory[28283] <=  8'h6e;        memory[28284] <=  8'h61;        memory[28285] <=  8'h62;        memory[28286] <=  8'h61;        memory[28287] <=  8'h63;        memory[28288] <=  8'h61;        memory[28289] <=  8'h74;        memory[28290] <=  8'h61;        memory[28291] <=  8'h62;        memory[28292] <=  8'h61;        memory[28293] <=  8'h72;        memory[28294] <=  8'h63;        memory[28295] <=  8'h61;        memory[28296] <=  8'h68;        memory[28297] <=  8'h64;        memory[28298] <=  8'h75;        memory[28299] <=  8'h63;        memory[28300] <=  8'h74;        memory[28301] <=  8'h61;        memory[28302] <=  8'h64;        memory[28303] <=  8'h61;        memory[28304] <=  8'h61;        memory[28305] <=  8'h63;        memory[28306] <=  8'h61;        memory[28307] <=  8'h72;        memory[28308] <=  8'h62;        memory[28309] <=  8'h61;        memory[28310] <=  8'h72;        memory[28311] <=  8'h74;        memory[28312] <=  8'h78;        memory[28313] <=  8'h61;        memory[28314] <=  8'h74;        memory[28315] <=  8'h6b;        memory[28316] <=  8'h73;        memory[28317] <=  8'h68;        memory[28318] <=  8'h63;        memory[28319] <=  8'h66;        memory[28320] <=  8'h69;        memory[28321] <=  8'h77;        memory[28322] <=  8'h68;        memory[28323] <=  8'h61;        memory[28324] <=  8'h74;        memory[28325] <=  8'h61;        memory[28326] <=  8'h6e;        memory[28327] <=  8'h61;        memory[28328] <=  8'h62;        memory[28329] <=  8'h61;        memory[28330] <=  8'h63;        memory[28331] <=  8'h61;        memory[28332] <=  8'h74;        memory[28333] <=  8'h61;        memory[28334] <=  8'h62;        memory[28335] <=  8'h61;        memory[28336] <=  8'h72;        memory[28337] <=  8'h63;        memory[28338] <=  8'h61;        memory[28339] <=  8'h68;        memory[28340] <=  8'h64;        memory[28341] <=  8'h75;        memory[28342] <=  8'h63;        memory[28343] <=  8'h74;        memory[28344] <=  8'h61;        memory[28345] <=  8'h64;        memory[28346] <=  8'h61;        memory[28347] <=  8'h61;        memory[28348] <=  8'h63;        memory[28349] <=  8'h61;        memory[28350] <=  8'h72;        memory[28351] <=  8'h62;        memory[28352] <=  8'h61;        memory[28353] <=  8'h72;        memory[28354] <=  8'h74;        memory[28355] <=  8'h78;        memory[28356] <=  8'h61;        memory[28357] <=  8'h74;        memory[28358] <=  8'h6b;        memory[28359] <=  8'h73;        memory[28360] <=  8'h68;        memory[28361] <=  8'h63;        memory[28362] <=  8'h66;        memory[28363] <=  8'h69;        memory[28364] <=  8'h77;        memory[28365] <=  8'h68;        memory[28366] <=  8'h61;        memory[28367] <=  8'h74;        memory[28368] <=  8'h61;        memory[28369] <=  8'h6e;        memory[28370] <=  8'h61;        memory[28371] <=  8'h62;        memory[28372] <=  8'h61;        memory[28373] <=  8'h63;        memory[28374] <=  8'h61;        memory[28375] <=  8'h74;        memory[28376] <=  8'h61;        memory[28377] <=  8'h62;        memory[28378] <=  8'h61;        memory[28379] <=  8'h72;        memory[28380] <=  8'h63;        memory[28381] <=  8'h61;        memory[28382] <=  8'h68;        memory[28383] <=  8'h64;        memory[28384] <=  8'h75;        memory[28385] <=  8'h63;        memory[28386] <=  8'h74;        memory[28387] <=  8'h61;        memory[28388] <=  8'h64;        memory[28389] <=  8'h61;        memory[28390] <=  8'h61;        memory[28391] <=  8'h63;        memory[28392] <=  8'h61;        memory[28393] <=  8'h72;        memory[28394] <=  8'h62;        memory[28395] <=  8'h61;        memory[28396] <=  8'h72;        memory[28397] <=  8'h74;        memory[28398] <=  8'h78;        memory[28399] <=  8'h61;        memory[28400] <=  8'h74;        memory[28401] <=  8'h6b;        memory[28402] <=  8'h73;        memory[28403] <=  8'h68;        memory[28404] <=  8'h63;        memory[28405] <=  8'h66;        memory[28406] <=  8'h69;        memory[28407] <=  8'h77;        memory[28408] <=  8'h68;        memory[28409] <=  8'h61;        memory[28410] <=  8'h74;        memory[28411] <=  8'h61;        memory[28412] <=  8'h6e;        memory[28413] <=  8'h61;        memory[28414] <=  8'h62;        memory[28415] <=  8'h61;        memory[28416] <=  8'h63;        memory[28417] <=  8'h61;        memory[28418] <=  8'h74;        memory[28419] <=  8'h61;        memory[28420] <=  8'h62;        memory[28421] <=  8'h61;        memory[28422] <=  8'h72;        memory[28423] <=  8'h63;        memory[28424] <=  8'h61;        memory[28425] <=  8'h68;        memory[28426] <=  8'h64;        memory[28427] <=  8'h75;        memory[28428] <=  8'h63;        memory[28429] <=  8'h74;        memory[28430] <=  8'h61;        memory[28431] <=  8'h64;        memory[28432] <=  8'h61;        memory[28433] <=  8'h61;        memory[28434] <=  8'h63;        memory[28435] <=  8'h61;        memory[28436] <=  8'h72;        memory[28437] <=  8'h62;        memory[28438] <=  8'h61;        memory[28439] <=  8'h72;        memory[28440] <=  8'h74;        memory[28441] <=  8'h74;        memory[28442] <=  8'h62;        memory[28443] <=  8'h61;        memory[28444] <=  8'h72;        memory[28445] <=  8'h74;        memory[28446] <=  8'h78;        memory[28447] <=  8'h61;        memory[28448] <=  8'h74;        memory[28449] <=  8'h6b;        memory[28450] <=  8'h73;        memory[28451] <=  8'h68;        memory[28452] <=  8'h63;        memory[28453] <=  8'h66;        memory[28454] <=  8'h69;        memory[28455] <=  8'h77;        memory[28456] <=  8'h68;        memory[28457] <=  8'h61;        memory[28458] <=  8'h74;        memory[28459] <=  8'h61;        memory[28460] <=  8'h6e;        memory[28461] <=  8'h61;        memory[28462] <=  8'h62;        memory[28463] <=  8'h61;        memory[28464] <=  8'h63;        memory[28465] <=  8'h61;        memory[28466] <=  8'h74;        memory[28467] <=  8'h61;        memory[28468] <=  8'h62;        memory[28469] <=  8'h61;        memory[28470] <=  8'h72;        memory[28471] <=  8'h63;        memory[28472] <=  8'h61;        memory[28473] <=  8'h68;        memory[28474] <=  8'h64;        memory[28475] <=  8'h75;        memory[28476] <=  8'h63;        memory[28477] <=  8'h74;        memory[28478] <=  8'h61;        memory[28479] <=  8'h64;        memory[28480] <=  8'h61;        memory[28481] <=  8'h61;        memory[28482] <=  8'h63;        memory[28483] <=  8'h61;        memory[28484] <=  8'h72;        memory[28485] <=  8'h63;        memory[28486] <=  8'h74;        memory[28487] <=  8'h72;        memory[28488] <=  8'h63;        memory[28489] <=  8'h61;        memory[28490] <=  8'h74;        memory[28491] <=  8'h72;        memory[28492] <=  8'h63;        memory[28493] <=  8'h61;        memory[28494] <=  8'h74;        memory[28495] <=  8'h63;        memory[28496] <=  8'h62;        memory[28497] <=  8'h61;        memory[28498] <=  8'h74;        memory[28499] <=  8'h62;        memory[28500] <=  8'h72;        memory[28501] <=  8'h63;        memory[28502] <=  8'h61;        memory[28503] <=  8'h72;        memory[28504] <=  8'h62;        memory[28505] <=  8'h78;        memory[28506] <=  8'h74;        memory[28507] <=  8'h61;        memory[28508] <=  8'h72;        memory[28509] <=  8'h64;        memory[28510] <=  8'h66;        memory[28511] <=  8'h73;        memory[28512] <=  8'h67;        memory[28513] <=  8'h76;        memory[28514] <=  8'h68;        memory[28515] <=  8'h62;        memory[28516] <=  8'h6b;        memory[28517] <=  8'h6a;        memory[28518] <=  8'h6e;        memory[28519] <=  8'h6d;        memory[28520] <=  8'h62;        memory[28521] <=  8'h76;        memory[28522] <=  8'h78;        memory[28523] <=  8'h63;        memory[28524] <=  8'h73;        memory[28525] <=  8'h66;        memory[28526] <=  8'h72;        memory[28527] <=  8'h74;        memory[28528] <=  8'h79;        memory[28529] <=  8'h75;        memory[28530] <=  8'h6a;        memory[28531] <=  8'h6e;        memory[28532] <=  8'h62;        memory[28533] <=  8'h76;        memory[28534] <=  8'h63;        memory[28535] <=  8'h64;        memory[28536] <=  8'h74;        memory[28537] <=  8'h79;        memory[28538] <=  8'h75;        memory[28539] <=  8'h69;        memory[28540] <=  8'h6b;        memory[28541] <=  8'h6d;        memory[28542] <=  8'h6e;        memory[28543] <=  8'h62;        memory[28544] <=  8'h76;        memory[28545] <=  8'h63;        memory[28546] <=  8'h78;        memory[28547] <=  8'h73;        memory[28548] <=  8'h64;        memory[28549] <=  8'h72;        memory[28550] <=  8'h74;        memory[28551] <=  8'h79;        memory[28552] <=  8'h75;        memory[28553] <=  8'h69;        memory[28554] <=  8'h6b;        memory[28555] <=  8'h6d;        memory[28556] <=  8'h6e;        memory[28557] <=  8'h62;        memory[28558] <=  8'h76;        memory[28559] <=  8'h63;        memory[28560] <=  8'h73;        memory[28561] <=  8'h77;        memory[28562] <=  8'h33;        memory[28563] <=  8'h34;        memory[28564] <=  8'h35;        memory[28565] <=  8'h36;        memory[28566] <=  8'h37;        memory[28567] <=  8'h38;        memory[28568] <=  8'h69;        memory[28569] <=  8'h6b;        memory[28570] <=  8'h6d;        memory[28571] <=  8'h6e;        memory[28572] <=  8'h62;        memory[28573] <=  8'h76;        memory[28574] <=  8'h63;        memory[28575] <=  8'h64;        memory[28576] <=  8'h65;        memory[28577] <=  8'h72;        memory[28578] <=  8'h36;        memory[28579] <=  8'h37;        memory[28580] <=  8'h38;        memory[28581] <=  8'h69;        memory[28582] <=  8'h6f;        memory[28583] <=  8'h6b;        memory[28584] <=  8'h6a;        memory[28585] <=  8'h6e;        memory[28586] <=  8'h62;        memory[28587] <=  8'h76;        memory[28588] <=  8'h63;        memory[28589] <=  8'h64;        memory[28590] <=  8'h72;        memory[28591] <=  8'h74;        memory[28592] <=  8'h79;        memory[28593] <=  8'h75;        memory[28594] <=  8'h73;        memory[28595] <=  8'h6a;        memory[28596] <=  8'h63;        memory[28597] <=  8'h6e;        memory[28598] <=  8'h62;        memory[28599] <=  8'h64;        memory[28600] <=  8'h66;        memory[28601] <=  8'h73;        memory[28602] <=  8'h74;        memory[28603] <=  8'h79;        memory[28604] <=  8'h75;        memory[28605] <=  8'h61;        memory[28606] <=  8'h69;        memory[28607] <=  8'h6b;        memory[28608] <=  8'h78;        memory[28609] <=  8'h6d;        memory[28610] <=  8'h6e;        memory[28611] <=  8'h73;        memory[28612] <=  8'h6a;        memory[28613] <=  8'h6f;        memory[28614] <=  8'h64;        memory[28615] <=  8'h6c;        memory[28616] <=  8'h63;        memory[28617] <=  8'h78;        memory[28618] <=  8'h2c;        memory[28619] <=  8'h6d;        memory[28620] <=  8'h73;        memory[28621] <=  8'h6b;        memory[28622] <=  8'h64;        memory[28623] <=  8'h6c;        memory[28624] <=  8'h70;        memory[28625] <=  8'h5b;        memory[28626] <=  8'h3b;        memory[28627] <=  8'h73;        memory[28628] <=  8'h6c;        memory[28629] <=  8'h64;        memory[28630] <=  8'h70;        memory[28631] <=  8'h76;        memory[28632] <=  8'h63;        memory[28633] <=  8'h5b;        memory[28634] <=  8'h78;        memory[28635] <=  8'h76;        memory[28636] <=  8'h63;        memory[28637] <=  8'h5b;        memory[28638] <=  8'h78;        memory[28639] <=  8'h70;        memory[28640] <=  8'h6f;        memory[28641] <=  8'h20;        memory[28642] <=  8'h62;        memory[28643] <=  8'h61;        memory[28644] <=  8'h72;        memory[28645] <=  8'h74;        memory[28646] <=  8'h74;        memory[28647] <=  8'h62;        memory[28648] <=  8'h61;        memory[28649] <=  8'h72;        memory[28650] <=  8'h74;        memory[28651] <=  8'h78;        memory[28652] <=  8'h61;        memory[28653] <=  8'h74;        memory[28654] <=  8'h6b;        memory[28655] <=  8'h73;        memory[28656] <=  8'h68;        memory[28657] <=  8'h63;        memory[28658] <=  8'h66;        memory[28659] <=  8'h69;        memory[28660] <=  8'h77;        memory[28661] <=  8'h68;        memory[28662] <=  8'h61;        memory[28663] <=  8'h69;        memory[28664] <=  8'h6a;        memory[28665] <=  8'h78;        memory[28666] <=  8'h5d;        memory[28667] <=  8'h65;        memory[28668] <=  8'h6b;        memory[28669] <=  8'h6f;        memory[28670] <=  8'h39;        memory[28671] <=  8'h64;        memory[28672] <=  8'h75;        memory[28673] <=  8'h38;        memory[28674] <=  8'h79;        memory[28675] <=  8'h20;        memory[28676] <=  8'h37;        memory[28677] <=  8'h63;        memory[28678] <=  8'h67;        memory[28679] <=  8'h78;        memory[28680] <=  8'h63;        memory[28681] <=  8'h75;        memory[28682] <=  8'h68;        memory[28683] <=  8'h69;        memory[28684] <=  8'h6a;        memory[28685] <=  8'h77;        memory[28686] <=  8'h69;        memory[28687] <=  8'h64;        memory[28688] <=  8'h66;        memory[28689] <=  8'h68;        memory[28690] <=  8'h75;        memory[28691] <=  8'h76;        memory[28692] <=  8'h64;        memory[28693] <=  8'h62;        memory[28694] <=  8'h66;        memory[28695] <=  8'h6a;        memory[28696] <=  8'h6e;        memory[28697] <=  8'h6b;        memory[28698] <=  8'h6a;        memory[28699] <=  8'h65;        memory[28700] <=  8'h38;        memory[28701] <=  8'h66;        memory[28702] <=  8'h37;        memory[28703] <=  8'h67;        memory[28704] <=  8'h79;        memory[28705] <=  8'h76;        memory[28706] <=  8'h63;        memory[28707] <=  8'h68;        memory[28708] <=  8'h69;        memory[28709] <=  8'h6a;        memory[28710] <=  8'h33;        memory[28711] <=  8'h65;        memory[28712] <=  8'h67;        memory[28713] <=  8'h79;        memory[28714] <=  8'h72;        memory[28715] <=  8'h64;        memory[28716] <=  8'h62;        memory[28717] <=  8'h6e;        memory[28718] <=  8'h63;        memory[28719] <=  8'h7a;        memory[28720] <=  8'h6a;        memory[28721] <=  8'h6f;        memory[28722] <=  8'h66;        memory[28723] <=  8'h78;        memory[28724] <=  8'h6a;        memory[28725] <=  8'h69;        memory[28726] <=  8'h63;        memory[28727] <=  8'h68;        memory[28728] <=  8'h62;        memory[28729] <=  8'h6e;        memory[28730] <=  8'h6d;        memory[28731] <=  8'h63;        memory[28732] <=  8'h73;        memory[28733] <=  8'h6c;        memory[28734] <=  8'h6b;        memory[28735] <=  8'h6a;        memory[28736] <=  8'h69;        memory[28737] <=  8'h68;        memory[28738] <=  8'h76;        memory[28739] <=  8'h75;        memory[28740] <=  8'h69;        memory[28741] <=  8'h64;        memory[28742] <=  8'h68;        memory[28743] <=  8'h75;        memory[28744] <=  8'h67;        memory[28745] <=  8'h79;        memory[28746] <=  8'h62;        memory[28747] <=  8'h68;        memory[28748] <=  8'h65;        memory[28749] <=  8'h6a;        memory[28750] <=  8'h72;        memory[28751] <=  8'h6b;        memory[28752] <=  8'h6a;        memory[28753] <=  8'h6f;        memory[28754] <=  8'h64;        memory[28755] <=  8'h67;        memory[28756] <=  8'h69;        memory[28757] <=  8'h75;        memory[28758] <=  8'h69;        memory[28759] <=  8'h67;        memory[28760] <=  8'h76;        memory[28761] <=  8'h79;        memory[28762] <=  8'h75;        memory[28763] <=  8'h67;        memory[28764] <=  8'h78;        memory[28765] <=  8'h68;        memory[28766] <=  8'h63;        memory[28767] <=  8'h20;        memory[28768] <=  8'h20;        memory[28769] <=  8'h20;        memory[28770] <=  8'h78;        memory[28771] <=  8'h76;        memory[28772] <=  8'h20;        memory[28773] <=  8'h63;        memory[28774] <=  8'h78;        memory[28775] <=  8'h67;        memory[28776] <=  8'h79;        memory[28777] <=  8'h63;        memory[28778] <=  8'h75;        memory[28779] <=  8'h68;        memory[28780] <=  8'h6a;        memory[28781] <=  8'h6b;        memory[28782] <=  8'h61;        memory[28783] <=  8'h6c;        memory[28784] <=  8'h78;        memory[28785] <=  8'h76;        memory[28786] <=  8'h70;        memory[28787] <=  8'h6f;        memory[28788] <=  8'h69;        memory[28789] <=  8'h6a;        memory[28790] <=  8'h69;        memory[28791] <=  8'h68;        memory[28792] <=  8'h6a;        memory[28793] <=  8'h62;        memory[28794] <=  8'h77;        memory[28795] <=  8'h65;        memory[28796] <=  8'h6e;        memory[28797] <=  8'h61;        memory[28798] <=  8'h66;        memory[28799] <=  8'h6d;        memory[28800] <=  8'h64;        memory[28801] <=  8'h6b;        memory[28802] <=  8'h6d;        memory[28803] <=  8'h76;        memory[28804] <=  8'h6c;        memory[28805] <=  8'h63;        memory[28806] <=  8'h6f;        memory[28807] <=  8'h64;        memory[28808] <=  8'h69;        memory[28809] <=  8'h75;        memory[28810] <=  8'h68;        memory[28811] <=  8'h73;        memory[28812] <=  8'h66;        memory[28813] <=  8'h65;        memory[28814] <=  8'h62;        memory[28815] <=  8'h6e;        memory[28816] <=  8'h64;        memory[28817] <=  8'h73;        memory[28818] <=  8'h63;        memory[28819] <=  8'h6b;        memory[28820] <=  8'h20;        memory[28821] <=  8'h78;        memory[28822] <=  8'h6a;        memory[28823] <=  8'h78;        memory[28824] <=  8'h63;        memory[28825] <=  8'h73;        memory[28826] <=  8'h64;        memory[28827] <=  8'h66;        memory[28828] <=  8'h6b;        memory[28829] <=  8'h64;        memory[28830] <=  8'h6e;        memory[28831] <=  8'h6d;        memory[28832] <=  8'h64;        memory[28833] <=  8'h73;        memory[28834] <=  8'h63;        memory[28835] <=  8'h6b;        memory[28836] <=  8'h78;        memory[28837] <=  8'h6c;        memory[28838] <=  8'h6f;        memory[28839] <=  8'h66;        memory[28840] <=  8'h6a;        memory[28841] <=  8'h69;        memory[28842] <=  8'h61;        memory[28843] <=  8'h62;        memory[28844] <=  8'h6e;        memory[28845] <=  8'h20;        memory[28846] <=  8'h78;        memory[28847] <=  8'h6b;        memory[28848] <=  8'h6d;        memory[28849] <=  8'h20;        memory[28850] <=  8'h6f;        memory[28851] <=  8'h63;        memory[28852] <=  8'h76;        memory[28853] <=  8'h73;        memory[28854] <=  8'h64;        memory[28855] <=  8'h69;        memory[28856] <=  8'h66;        memory[28857] <=  8'h68;        memory[28858] <=  8'h65;        memory[28859] <=  8'h71;        memory[28860] <=  8'h6a;        memory[28861] <=  8'h77;        memory[28862] <=  8'h62;        memory[28863] <=  8'h65;        memory[28864] <=  8'h6e;        memory[28865] <=  8'h20;        memory[28866] <=  8'h6d;        memory[28867] <=  8'h64;        memory[28868] <=  8'h73;        memory[28869] <=  8'h6c;        memory[28870] <=  8'h76;        memory[28871] <=  8'h6b;        memory[28872] <=  8'h63;        memory[28873] <=  8'h78;        memory[28874] <=  8'h20;        memory[28875] <=  8'h6f;        memory[28876] <=  8'h78;        memory[28877] <=  8'h69;        memory[28878] <=  8'h63;        memory[28879] <=  8'h6a;        memory[28880] <=  8'h76;        memory[28881] <=  8'h64;        memory[28882] <=  8'h66;        memory[28883] <=  8'h65;        memory[28884] <=  8'h71;        memory[28885] <=  8'h6e;        memory[28886] <=  8'h20;        memory[28887] <=  8'h64;        memory[28888] <=  8'h6d;        memory[28889] <=  8'h73;        memory[28890] <=  8'h6c;        memory[28891] <=  8'h63;        memory[28892] <=  8'h78;        memory[28893] <=  8'h6b;        memory[28894] <=  8'h20;        memory[28895] <=  8'h6f;        memory[28896] <=  8'h78;        memory[28897] <=  8'h63;        memory[28898] <=  8'h76;        memory[28899] <=  8'h6a;        memory[28900] <=  8'h64;        memory[28901] <=  8'h62;        memory[28902] <=  8'h71;        memory[28903] <=  8'h77;        memory[28904] <=  8'h65;        memory[28905] <=  8'h6e;        memory[28906] <=  8'h6d;        memory[28907] <=  8'h64;        memory[28908] <=  8'h6c;        memory[28909] <=  8'h73;        memory[28910] <=  8'h2c;        memory[28911] <=  8'h76;        memory[28912] <=  8'h63;        memory[28913] <=  8'h78;        memory[28914] <=  8'h20;        memory[28915] <=  8'h63;        memory[28916] <=  8'h6f;        memory[28917] <=  8'h69;        memory[28918] <=  8'h76;        memory[28919] <=  8'h68;        memory[28920] <=  8'h73;        memory[28921] <=  8'h64;        memory[28922] <=  8'h62;        memory[28923] <=  8'h71;        memory[28924] <=  8'h77;        memory[28925] <=  8'h65;        memory[28926] <=  8'h6e;        memory[28927] <=  8'h64;        memory[28928] <=  8'h6b;        memory[28929] <=  8'h73;        memory[28930] <=  8'h76;        memory[28931] <=  8'h6f;        memory[28932] <=  8'h63;        memory[28933] <=  8'h20;        memory[28934] <=  8'h76;        memory[28935] <=  8'h69;        memory[28936] <=  8'h75;        memory[28937] <=  8'h69;        memory[28938] <=  8'h68;        memory[28939] <=  8'h63;        memory[28940] <=  8'h78;        memory[28941] <=  8'h69;        memory[28942] <=  8'h6f;        memory[28943] <=  8'h76;        memory[28944] <=  8'h73;        memory[28945] <=  8'h64;        memory[28946] <=  8'h61;        memory[28947] <=  8'h64;        memory[28948] <=  8'h6e;        memory[28949] <=  8'h77;        memory[28950] <=  8'h71;        memory[28951] <=  8'h6b;        memory[28952] <=  8'h6c;        memory[28953] <=  8'h73;        memory[28954] <=  8'h76;        memory[28955] <=  8'h6e;        memory[28956] <=  8'h62;        memory[28957] <=  8'h20;        memory[28958] <=  8'h64;        memory[28959] <=  8'h66;        memory[28960] <=  8'h6a;        memory[28961] <=  8'h6b;        memory[28962] <=  8'h71;        memory[28963] <=  8'h64;        memory[28964] <=  8'h77;        memory[28965] <=  8'h65;        memory[28966] <=  8'h6e;        memory[28967] <=  8'h62;        memory[28968] <=  8'h20;        memory[28969] <=  8'h64;        memory[28970] <=  8'h73;        memory[28971] <=  8'h76;        memory[28972] <=  8'h68;        memory[28973] <=  8'h64;        memory[28974] <=  8'h61;        memory[28975] <=  8'h71;        memory[28976] <=  8'h77;        memory[28977] <=  8'h6a;        memory[28978] <=  8'h65;        memory[28979] <=  8'h6e;        memory[28980] <=  8'h64;        memory[28981] <=  8'h20;        memory[28982] <=  8'h61;        memory[28983] <=  8'h63;        memory[28984] <=  8'h62;        memory[28985] <=  8'h68;        memory[28986] <=  8'h64;        memory[28987] <=  8'h61;        memory[28988] <=  8'h77;        memory[28989] <=  8'h71;        memory[28990] <=  8'h6e;        memory[28991] <=  8'h20;        memory[28992] <=  8'h62;        memory[28993] <=  8'h73;        memory[28994] <=  8'h76;        memory[28995] <=  8'h61;        memory[28996] <=  8'h67;        memory[28997] <=  8'h76;        memory[28998] <=  8'h68;        memory[28999] <=  8'h67;        memory[29000] <=  8'h61;        memory[29001] <=  8'h73;        memory[29002] <=  8'h6a;        memory[29003] <=  8'h6b;        memory[29004] <=  8'h63;        memory[29005] <=  8'h78;        memory[29006] <=  8'h76;        memory[29007] <=  8'h6e;        memory[29008] <=  8'h73;        memory[29009] <=  8'h64;        memory[29010] <=  8'h20;        memory[29011] <=  8'h66;        memory[29012] <=  8'h62;        memory[29013] <=  8'h64;        memory[29014] <=  8'h61;        memory[29015] <=  8'h73;        memory[29016] <=  8'h76;        memory[29017] <=  8'h67;        memory[29018] <=  8'h63;        memory[29019] <=  8'h79;        memory[29020] <=  8'h7a;        memory[29021] <=  8'h78;        memory[29022] <=  8'h79;        memory[29023] <=  8'h75;        memory[29024] <=  8'h20;        memory[29025] <=  8'h69;        memory[29026] <=  8'h6a;        memory[29027] <=  8'h64;        memory[29028] <=  8'h66;        memory[29029] <=  8'h6b;        memory[29030] <=  8'h61;        memory[29031] <=  8'h64;        memory[29032] <=  8'h63;        memory[29033] <=  8'h78;        memory[29034] <=  8'h68;        memory[29035] <=  8'h20;        memory[29036] <=  8'h67;        memory[29037] <=  8'h61;        memory[29038] <=  8'h68;        memory[29039] <=  8'h75;        memory[29040] <=  8'h64;        memory[29041] <=  8'h73;        memory[29042] <=  8'h69;        memory[29043] <=  8'h6a;        memory[29044] <=  8'h61;        memory[29045] <=  8'h6b;        memory[29046] <=  8'h63;        memory[29047] <=  8'h62;        memory[29048] <=  8'h61;        memory[29049] <=  8'h72;        memory[29050] <=  8'h73;        memory[29051] <=  8'h68;        memory[29052] <=  8'h64;        memory[29053] <=  8'h66;        memory[29054] <=  8'h67;        memory[29055] <=  8'h73;        memory[29056] <=  8'h68;        memory[29057] <=  8'h64;        memory[29058] <=  8'h66;        memory[29059] <=  8'h68;        memory[29060] <=  8'h64;        memory[29061] <=  8'h6a;        memory[29062] <=  8'h68;        memory[29063] <=  8'h62;        memory[29064] <=  8'h67;        memory[29065] <=  8'h63;        memory[29066] <=  8'h61;        memory[29067] <=  8'h66;        memory[29068] <=  8'h73;        memory[29069] <=  8'h79;        memory[29070] <=  8'h67;        memory[29071] <=  8'h6b;        memory[29072] <=  8'h75;        memory[29073] <=  8'h64;        memory[29074] <=  8'h68;        memory[29075] <=  8'h62;        memory[29076] <=  8'h77;        memory[29077] <=  8'h76;        memory[29078] <=  8'h67;        memory[29079] <=  8'h61;        memory[29080] <=  8'h66;        memory[29081] <=  8'h64;        memory[29082] <=  8'h74;        memory[29083] <=  8'h75;        memory[29084] <=  8'h66;        memory[29085] <=  8'h79;        memory[29086] <=  8'h67;        memory[29087] <=  8'h69;        memory[29088] <=  8'h75;        memory[29089] <=  8'h68;        memory[29090] <=  8'h6c;        memory[29091] <=  8'h6a;        memory[29092] <=  8'h62;        memory[29093] <=  8'h6b;        memory[29094] <=  8'h68;        memory[29095] <=  8'h76;        memory[29096] <=  8'h67;        memory[29097] <=  8'h63;        memory[29098] <=  8'h66;        memory[29099] <=  8'h78;        memory[29100] <=  8'h64;        memory[29101] <=  8'h74;        memory[29102] <=  8'h75;        memory[29103] <=  8'h79;        memory[29104] <=  8'h69;        memory[29105] <=  8'h75;        memory[29106] <=  8'h68;        memory[29107] <=  8'h6c;        memory[29108] <=  8'h6a;        memory[29109] <=  8'h6b;        memory[29110] <=  8'h67;        memory[29111] <=  8'h6a;        memory[29112] <=  8'h63;        memory[29113] <=  8'h66;        memory[29114] <=  8'h68;        memory[29115] <=  8'h64;        memory[29116] <=  8'h67;        memory[29117] <=  8'h72;        memory[29118] <=  8'h79;        memory[29119] <=  8'h74;        memory[29120] <=  8'h66;        memory[29121] <=  8'h75;        memory[29122] <=  8'h79;        memory[29123] <=  8'h69;        memory[29124] <=  8'h68;        memory[29125] <=  8'h6c;        memory[29126] <=  8'h62;        memory[29127] <=  8'h6d;        memory[29128] <=  8'h76;        memory[29129] <=  8'h6e;        memory[29130] <=  8'h63;        memory[29131] <=  8'h66;        memory[29132] <=  8'h68;        memory[29133] <=  8'h64;        memory[29134] <=  8'h74;        memory[29135] <=  8'h75;        memory[29136] <=  8'h67;        memory[29137] <=  8'h79;        memory[29138] <=  8'h69;        memory[29139] <=  8'h68;        memory[29140] <=  8'h75;        memory[29141] <=  8'h6a;        memory[29142] <=  8'h6c;        memory[29143] <=  8'h62;        memory[29144] <=  8'h6d;        memory[29145] <=  8'h76;        memory[29146] <=  8'h6e;        memory[29147] <=  8'h63;        memory[29148] <=  8'h66;        memory[29149] <=  8'h68;        memory[29150] <=  8'h67;        memory[29151] <=  8'h79;        memory[29152] <=  8'h68;        memory[29153] <=  8'h75;        memory[29154] <=  8'h6a;        memory[29155] <=  8'h6e;        memory[29156] <=  8'h2c;        memory[29157] <=  8'h62;        memory[29158] <=  8'h6e;        memory[29159] <=  8'h6d;        memory[29160] <=  8'h76;        memory[29161] <=  8'h6e;        memory[29162] <=  8'h63;        memory[29163] <=  8'h66;        memory[29164] <=  8'h68;        memory[29165] <=  8'h74;        memory[29166] <=  8'h79;        memory[29167] <=  8'h69;        memory[29168] <=  8'h75;        memory[29169] <=  8'h6c;        memory[29170] <=  8'h6a;        memory[29171] <=  8'h62;        memory[29172] <=  8'h6d;        memory[29173] <=  8'h76;        memory[29174] <=  8'h6e;        memory[29175] <=  8'h63;        memory[29176] <=  8'h66;        memory[29177] <=  8'h74;        memory[29178] <=  8'h75;        memory[29179] <=  8'h79;        memory[29180] <=  8'h69;        memory[29181] <=  8'h68;        memory[29182] <=  8'h6b;        memory[29183] <=  8'h62;        memory[29184] <=  8'h76;        memory[29185] <=  8'h63;        memory[29186] <=  8'h66;        memory[29187] <=  8'h67;        memory[29188] <=  8'h74;        memory[29189] <=  8'h75;        memory[29190] <=  8'h79;        memory[29191] <=  8'h69;        memory[29192] <=  8'h75;        memory[29193] <=  8'h68;        memory[29194] <=  8'h6a;        memory[29195] <=  8'h6b;        memory[29196] <=  8'h62;        memory[29197] <=  8'h76;        memory[29198] <=  8'h63;        memory[29199] <=  8'h66;        memory[29200] <=  8'h74;        memory[29201] <=  8'h75;        memory[29202] <=  8'h79;        memory[29203] <=  8'h69;        memory[29204] <=  8'h75;        memory[29205] <=  8'h6a;        memory[29206] <=  8'h6b;        memory[29207] <=  8'h6e;        memory[29208] <=  8'h62;        memory[29209] <=  8'h76;        memory[29210] <=  8'h67;        memory[29211] <=  8'h66;        memory[29212] <=  8'h74;        memory[29213] <=  8'h79;        memory[29214] <=  8'h75;        memory[29215] <=  8'h75;        memory[29216] <=  8'h69;        memory[29217] <=  8'h6a;        memory[29218] <=  8'h6b;        memory[29219] <=  8'h68;        memory[29220] <=  8'h62;        memory[29221] <=  8'h6a;        memory[29222] <=  8'h67;        memory[29223] <=  8'h68;        memory[29224] <=  8'h66;        memory[29225] <=  8'h79;        memory[29226] <=  8'h74;        memory[29227] <=  8'h79;        memory[29228] <=  8'h69;        memory[29229] <=  8'h75;        memory[29230] <=  8'h64;        memory[29231] <=  8'h6a;        memory[29232] <=  8'h6b;        memory[29233] <=  8'h68;        memory[29234] <=  8'h63;        memory[29235] <=  8'h7a;        memory[29236] <=  8'h67;        memory[29237] <=  8'h68;        memory[29238] <=  8'h74;        memory[29239] <=  8'h75;        memory[29240] <=  8'h79;        memory[29241] <=  8'h69;        memory[29242] <=  8'h61;        memory[29243] <=  8'h73;        memory[29244] <=  8'h75;        memory[29245] <=  8'h6a;        memory[29246] <=  8'h6b;        memory[29247] <=  8'h62;        memory[29248] <=  8'h6e;        memory[29249] <=  8'h61;        memory[29250] <=  8'h76;        memory[29251] <=  8'h63;        memory[29252] <=  8'h66;        memory[29253] <=  8'h68;        memory[29254] <=  8'h75;        memory[29255] <=  8'h61;        memory[29256] <=  8'h73;        memory[29257] <=  8'h79;        memory[29258] <=  8'h64;        memory[29259] <=  8'h75;        memory[29260] <=  8'h69;        memory[29261] <=  8'h6a;        memory[29262] <=  8'h61;        memory[29263] <=  8'h6b;        memory[29264] <=  8'h62;        memory[29265] <=  8'h63;        memory[29266] <=  8'h78;        memory[29267] <=  8'h68;        memory[29268] <=  8'h67;        memory[29269] <=  8'h79;        memory[29270] <=  8'h75;        memory[29271] <=  8'h7a;        memory[29272] <=  8'h63;        memory[29273] <=  8'h61;        memory[29274] <=  8'h73;        memory[29275] <=  8'h69;        memory[29276] <=  8'h75;        memory[29277] <=  8'h6f;        memory[29278] <=  8'h69;        memory[29279] <=  8'h6a;        memory[29280] <=  8'h61;        memory[29281] <=  8'h6c;        memory[29282] <=  8'h63;        memory[29283] <=  8'h78;        memory[29284] <=  8'h62;        memory[29285] <=  8'h63;        memory[29286] <=  8'h20;        memory[29287] <=  8'h6e;        memory[29288] <=  8'h76;        memory[29289] <=  8'h63;        memory[29290] <=  8'h61;        memory[29291] <=  8'h64;        memory[29292] <=  8'h73;        memory[29293] <=  8'h67;        memory[29294] <=  8'h79;        memory[29295] <=  8'h68;        memory[29296] <=  8'h75;        memory[29297] <=  8'h61;        memory[29298] <=  8'h6a;        memory[29299] <=  8'h6b;        memory[29300] <=  8'h78;        memory[29301] <=  8'h62;        memory[29302] <=  8'h20;        memory[29303] <=  8'h6e;        memory[29304] <=  8'h76;        memory[29305] <=  8'h63;        memory[29306] <=  8'h61;        memory[29307] <=  8'h73;        memory[29308] <=  8'h67;        memory[29309] <=  8'h68;        memory[29310] <=  8'h75;        memory[29311] <=  8'h6a;        memory[29312] <=  8'h6c;        memory[29313] <=  8'h6b;        memory[29314] <=  8'h63;        memory[29315] <=  8'h78;        memory[29316] <=  8'h20;        memory[29317] <=  8'h6a;        memory[29318] <=  8'h6b;        memory[29319] <=  8'h68;        memory[29320] <=  8'h61;        memory[29321] <=  8'h73;        memory[29322] <=  8'h76;        memory[29323] <=  8'h64;        memory[29324] <=  8'h6e;        memory[29325] <=  8'h20;        memory[29326] <=  8'h62;        memory[29327] <=  8'h6e;        memory[29328] <=  8'h6d;        memory[29329] <=  8'h6b;        memory[29330] <=  8'h77;        memory[29331] <=  8'h64;        memory[29332] <=  8'h6f;        memory[29333] <=  8'h77;        memory[29334] <=  8'h69;        memory[29335] <=  8'h6f;        memory[29336] <=  8'h75;        memory[29337] <=  8'h69;        memory[29338] <=  8'h68;        memory[29339] <=  8'h62;        memory[29340] <=  8'h6e;        memory[29341] <=  8'h6b;        memory[29342] <=  8'h77;        memory[29343] <=  8'h69;        memory[29344] <=  8'h6f;        memory[29345] <=  8'h75;        memory[29346] <=  8'h71;        memory[29347] <=  8'h69;        memory[29348] <=  8'h79;        memory[29349] <=  8'h67;        memory[29350] <=  8'h6a;        memory[29351] <=  8'h64;        memory[29352] <=  8'h61;        memory[29353] <=  8'h76;        memory[29354] <=  8'h62;        memory[29355] <=  8'h6e;        memory[29356] <=  8'h6b;        memory[29357] <=  8'h6f;        memory[29358] <=  8'h70;        memory[29359] <=  8'h64;        memory[29360] <=  8'h76;        memory[29361] <=  8'h69;        memory[29362] <=  8'h6f;        memory[29363] <=  8'h75;        memory[29364] <=  8'h69;        memory[29365] <=  8'h48;        memory[29366] <=  8'h42;        memory[29367] <=  8'h6b;        memory[29368] <=  8'h64;        memory[29369] <=  8'h6e;        memory[29370] <=  8'h6c;        memory[29371] <=  8'h71;        memory[29372] <=  8'h6b;        memory[29373] <=  8'h6d;        memory[29374] <=  8'h6a;        memory[29375] <=  8'h70;        memory[29376] <=  8'h69;        memory[29377] <=  8'h6f;        memory[29378] <=  8'h68;        memory[29379] <=  8'h65;        memory[29380] <=  8'h66;        memory[29381] <=  8'h75;        memory[29382] <=  8'h67;        memory[29383] <=  8'h69;        memory[29384] <=  8'h73;        memory[29385] <=  8'h61;        memory[29386] <=  8'h62;        memory[29387] <=  8'h64;        memory[29388] <=  8'h6b;        memory[29389] <=  8'h6a;        memory[29390] <=  8'h6b;        memory[29391] <=  8'h6c;        memory[29392] <=  8'h6a;        memory[29393] <=  8'h69;        memory[29394] <=  8'h73;        memory[29395] <=  8'h6f;        memory[29396] <=  8'h71;        memory[29397] <=  8'h68;        memory[29398] <=  8'h77;        memory[29399] <=  8'h67;        memory[29400] <=  8'h69;        memory[29401] <=  8'h79;        memory[29402] <=  8'h6a;        memory[29403] <=  8'h64;        memory[29404] <=  8'h76;        memory[29405] <=  8'h62;        memory[29406] <=  8'h6e;        memory[29407] <=  8'h61;        memory[29408] <=  8'h73;        memory[29409] <=  8'h66;        memory[29410] <=  8'h6c;        memory[29411] <=  8'h6b;        memory[29412] <=  8'h64;        memory[29413] <=  8'h6a;        memory[29414] <=  8'h68;        memory[29415] <=  8'h63;        memory[29416] <=  8'h67;        memory[29417] <=  8'h6a;        memory[29418] <=  8'h76;        memory[29419] <=  8'h73;        memory[29420] <=  8'h64;        memory[29421] <=  8'h62;        memory[29422] <=  8'h62;        memory[29423] <=  8'h61;        memory[29424] <=  8'h72;        memory[29425] <=  8'h62;        memory[29426] <=  8'h62;        memory[29427] <=  8'h73;        memory[29428] <=  8'h62;        memory[29429] <=  8'h67;        memory[29430] <=  8'h73;        memory[29431] <=  8'h66;        memory[29432] <=  8'h67;        memory[29433] <=  8'h61;        memory[29434] <=  8'h68;        memory[29435] <=  8'h66;        memory[29436] <=  8'h73;        memory[29437] <=  8'h68;        memory[29438] <=  8'h61;        memory[29439] <=  8'h66;        memory[29440] <=  8'h73;        memory[29441] <=  8'h66;        memory[29442] <=  8'h68;        memory[29443] <=  8'h61;        memory[29444] <=  8'h69;        memory[29445] <=  8'h64;        memory[29446] <=  8'h75;        memory[29447] <=  8'h67;        memory[29448] <=  8'h64;        memory[29449] <=  8'h77;        memory[29450] <=  8'h62;        memory[29451] <=  8'h61;        memory[29452] <=  8'h62;        memory[29453] <=  8'h72;        memory[29454] <=  8'h62;        memory[29455] <=  8'h61;        memory[29456] <=  8'h62;        memory[29457] <=  8'h62;        memory[29458] <=  8'h74;        memory[29459] <=  8'h62;        memory[29460] <=  8'h62;        memory[29461] <=  8'h62;        memory[29462] <=  8'h62;        memory[29463] <=  8'h62;        memory[29464] <=  8'h62;        memory[29465] <=  8'h62;        memory[29466] <=  8'h62;        memory[29467] <=  8'h61;        memory[29468] <=  8'h62;        memory[29469] <=  8'h62;        memory[29470] <=  8'h72;        memory[29471] <=  8'h74;        memory[29472] <=  8'h62;        memory[29473] <=  8'h62;        memory[29474] <=  8'h61;        memory[29475] <=  8'h62;        memory[29476] <=  8'h72;        memory[29477] <=  8'h62;        memory[29478] <=  8'h74;        memory[29479] <=  8'h62;        memory[29480] <=  8'h62;        memory[29481] <=  8'h62;        memory[29482] <=  8'h63;        memory[29483] <=  8'h61;        memory[29484] <=  8'h72;        memory[29485] <=  8'h74;        memory[29486] <=  8'h73;        memory[29487] <=  8'h62;        memory[29488] <=  8'h61;        memory[29489] <=  8'h72;        memory[29490] <=  8'h74;        memory[29491] <=  8'h74;        memory[29492] <=  8'h62;        memory[29493] <=  8'h61;        memory[29494] <=  8'h72;        memory[29495] <=  8'h74;        memory[29496] <=  8'h78;        memory[29497] <=  8'h61;        memory[29498] <=  8'h74;        memory[29499] <=  8'h6b;        memory[29500] <=  8'h73;        memory[29501] <=  8'h68;        memory[29502] <=  8'h63;        memory[29503] <=  8'h66;        memory[29504] <=  8'h69;        memory[29505] <=  8'h77;        memory[29506] <=  8'h68;        memory[29507] <=  8'h61;        memory[29508] <=  8'h74;        memory[29509] <=  8'h61;        memory[29510] <=  8'h6e;        memory[29511] <=  8'h61;        memory[29512] <=  8'h62;        memory[29513] <=  8'h61;        memory[29514] <=  8'h63;        memory[29515] <=  8'h61;        memory[29516] <=  8'h74;        memory[29517] <=  8'h61;        memory[29518] <=  8'h62;        memory[29519] <=  8'h61;        memory[29520] <=  8'h72;        memory[29521] <=  8'h63;        memory[29522] <=  8'h61;        memory[29523] <=  8'h68;        memory[29524] <=  8'h64;        memory[29525] <=  8'h75;        memory[29526] <=  8'h63;        memory[29527] <=  8'h74;        memory[29528] <=  8'h61;        memory[29529] <=  8'h64;        memory[29530] <=  8'h61;        memory[29531] <=  8'h61;        memory[29532] <=  8'h63;        memory[29533] <=  8'h61;        memory[29534] <=  8'h72;        memory[29535] <=  8'h63;        memory[29536] <=  8'h74;        memory[29537] <=  8'h72;        memory[29538] <=  8'h63;        memory[29539] <=  8'h61;        memory[29540] <=  8'h74;        memory[29541] <=  8'h72;        memory[29542] <=  8'h63;        memory[29543] <=  8'h61;        memory[29544] <=  8'h74;        memory[29545] <=  8'h63;        memory[29546] <=  8'h62;        memory[29547] <=  8'h61;        memory[29548] <=  8'h74;        memory[29549] <=  8'h62;        memory[29550] <=  8'h72;        memory[29551] <=  8'h63;        memory[29552] <=  8'h61;        memory[29553] <=  8'h74;        memory[29554] <=  8'h72;        memory[29555] <=  8'h6e;        memory[29556] <=  8'h62;        memory[29557] <=  8'h61;        memory[29558] <=  8'h63;        memory[29559] <=  8'h61;        memory[29560] <=  8'h74;        memory[29561] <=  8'h79;        memory[29562] <=  8'h73;        memory[29563] <=  8'h6e;        memory[29564] <=  8'h63;        memory[29565] <=  8'h74;        memory[29566] <=  8'h61;        memory[29567] <=  8'h6e;        memory[29568] <=  8'h62;        memory[29569] <=  8'h61;        memory[29570] <=  8'h63;        memory[29571] <=  8'h72;        memory[29572] <=  8'h6e;        memory[29573] <=  8'h74;        memory[29574] <=  8'h61;        memory[29575] <=  8'h62;        memory[29576] <=  8'h74;        memory[29577] <=  8'h6e;        memory[29578] <=  8'h61;        memory[29579] <=  8'h72;        memory[29580] <=  8'h62;        memory[29581] <=  8'h78;        memory[29582] <=  8'h74;        memory[29583] <=  8'h61;        memory[29584] <=  8'h72;        memory[29585] <=  8'h62;        memory[29586] <=  8'h61;        memory[29587] <=  8'h72;        memory[29588] <=  8'h74;        memory[29589] <=  8'h74;        memory[29590] <=  8'h62;        memory[29591] <=  8'h61;        memory[29592] <=  8'h72;        memory[29593] <=  8'h74;        memory[29594] <=  8'h78;        memory[29595] <=  8'h61;        memory[29596] <=  8'h74;        memory[29597] <=  8'h6b;        memory[29598] <=  8'h73;        memory[29599] <=  8'h68;        memory[29600] <=  8'h63;        memory[29601] <=  8'h66;        memory[29602] <=  8'h69;        memory[29603] <=  8'h77;        memory[29604] <=  8'h68;        memory[29605] <=  8'h61;        memory[29606] <=  8'h74;        memory[29607] <=  8'h61;        memory[29608] <=  8'h6e;        memory[29609] <=  8'h61;        memory[29610] <=  8'h62;        memory[29611] <=  8'h61;        memory[29612] <=  8'h63;        memory[29613] <=  8'h61;        memory[29614] <=  8'h74;        memory[29615] <=  8'h61;        memory[29616] <=  8'h62;        memory[29617] <=  8'h61;        memory[29618] <=  8'h72;        memory[29619] <=  8'h63;        memory[29620] <=  8'h61;        memory[29621] <=  8'h68;        memory[29622] <=  8'h64;        memory[29623] <=  8'h75;        memory[29624] <=  8'h63;        memory[29625] <=  8'h74;        memory[29626] <=  8'h61;        memory[29627] <=  8'h64;        memory[29628] <=  8'h61;        memory[29629] <=  8'h61;        memory[29630] <=  8'h63;        memory[29631] <=  8'h61;        memory[29632] <=  8'h72;        memory[29633] <=  8'h63;        memory[29634] <=  8'h74;        memory[29635] <=  8'h72;        memory[29636] <=  8'h63;        memory[29637] <=  8'h61;        memory[29638] <=  8'h74;        memory[29639] <=  8'h72;        memory[29640] <=  8'h63;        memory[29641] <=  8'h61;        memory[29642] <=  8'h74;        memory[29643] <=  8'h63;        memory[29644] <=  8'h62;        memory[29645] <=  8'h61;        memory[29646] <=  8'h74;        memory[29647] <=  8'h62;        memory[29648] <=  8'h72;        memory[29649] <=  8'h63;        memory[29650] <=  8'h61;        memory[29651] <=  8'h74;        memory[29652] <=  8'h72;        memory[29653] <=  8'h6e;        memory[29654] <=  8'h62;        memory[29655] <=  8'h61;        memory[29656] <=  8'h63;        memory[29657] <=  8'h61;        memory[29658] <=  8'h74;        memory[29659] <=  8'h79;        memory[29660] <=  8'h73;        memory[29661] <=  8'h6e;        memory[29662] <=  8'h63;        memory[29663] <=  8'h74;        memory[29664] <=  8'h61;        memory[29665] <=  8'h6e;        memory[29666] <=  8'h62;        memory[29667] <=  8'h61;        memory[29668] <=  8'h63;        memory[29669] <=  8'h72;        memory[29670] <=  8'h6e;        memory[29671] <=  8'h74;        memory[29672] <=  8'h61;        memory[29673] <=  8'h62;        memory[29674] <=  8'h74;        memory[29675] <=  8'h6e;        memory[29676] <=  8'h61;        memory[29677] <=  8'h72;        memory[29678] <=  8'h62;        memory[29679] <=  8'h78;        memory[29680] <=  8'h74;        memory[29681] <=  8'h61;        memory[29682] <=  8'h72;        memory[29683] <=  8'h62;        memory[29684] <=  8'h61;        memory[29685] <=  8'h72;        memory[29686] <=  8'h74;        memory[29687] <=  8'h74;        memory[29688] <=  8'h62;        memory[29689] <=  8'h61;        memory[29690] <=  8'h72;        memory[29691] <=  8'h74;        memory[29692] <=  8'h78;        memory[29693] <=  8'h61;        memory[29694] <=  8'h74;        memory[29695] <=  8'h6b;        memory[29696] <=  8'h73;        memory[29697] <=  8'h68;        memory[29698] <=  8'h63;        memory[29699] <=  8'h66;        memory[29700] <=  8'h69;        memory[29701] <=  8'h77;        memory[29702] <=  8'h68;        memory[29703] <=  8'h61;        memory[29704] <=  8'h74;        memory[29705] <=  8'h61;        memory[29706] <=  8'h6e;        memory[29707] <=  8'h61;        memory[29708] <=  8'h62;        memory[29709] <=  8'h61;        memory[29710] <=  8'h63;        memory[29711] <=  8'h61;        memory[29712] <=  8'h74;        memory[29713] <=  8'h61;        memory[29714] <=  8'h62;        memory[29715] <=  8'h61;        memory[29716] <=  8'h72;        memory[29717] <=  8'h63;        memory[29718] <=  8'h61;        memory[29719] <=  8'h68;        memory[29720] <=  8'h64;        memory[29721] <=  8'h75;        memory[29722] <=  8'h63;        memory[29723] <=  8'h74;        memory[29724] <=  8'h61;        memory[29725] <=  8'h64;        memory[29726] <=  8'h61;        memory[29727] <=  8'h61;        memory[29728] <=  8'h63;        memory[29729] <=  8'h61;        memory[29730] <=  8'h72;        memory[29731] <=  8'h63;        memory[29732] <=  8'h74;        memory[29733] <=  8'h72;        memory[29734] <=  8'h63;        memory[29735] <=  8'h61;        memory[29736] <=  8'h74;        memory[29737] <=  8'h72;        memory[29738] <=  8'h63;        memory[29739] <=  8'h61;        memory[29740] <=  8'h74;        memory[29741] <=  8'h63;        memory[29742] <=  8'h62;        memory[29743] <=  8'h61;        memory[29744] <=  8'h74;        memory[29745] <=  8'h62;        memory[29746] <=  8'h72;        memory[29747] <=  8'h63;        memory[29748] <=  8'h61;        memory[29749] <=  8'h74;        memory[29750] <=  8'h72;        memory[29751] <=  8'h6e;        memory[29752] <=  8'h62;        memory[29753] <=  8'h61;        memory[29754] <=  8'h63;        memory[29755] <=  8'h61;        memory[29756] <=  8'h74;        memory[29757] <=  8'h79;        memory[29758] <=  8'h73;        memory[29759] <=  8'h6e;        memory[29760] <=  8'h63;        memory[29761] <=  8'h74;        memory[29762] <=  8'h61;        memory[29763] <=  8'h6e;        memory[29764] <=  8'h62;        memory[29765] <=  8'h61;        memory[29766] <=  8'h63;        memory[29767] <=  8'h72;        memory[29768] <=  8'h6e;        memory[29769] <=  8'h74;        memory[29770] <=  8'h61;        memory[29771] <=  8'h62;        memory[29772] <=  8'h74;        memory[29773] <=  8'h6e;        memory[29774] <=  8'h61;        memory[29775] <=  8'h72;        memory[29776] <=  8'h62;        memory[29777] <=  8'h78;        memory[29778] <=  8'h74;        memory[29779] <=  8'h61;        memory[29780] <=  8'h72;        memory[29781] <=  8'h5d;        memory[29782] <=  8'h5d;        memory[29783] <=  8'h65;        memory[29784] <=  8'h66;        memory[29785] <=  8'h77;        memory[29786] <=  8'h65;        memory[29787] <=  8'h5d;        memory[29788] <=  8'h65;        memory[29789] <=  8'h67;        memory[29790] <=  8'h73;        memory[29791] <=  8'h67;        memory[29792] <=  8'h66;        memory[29793] <=  8'h62;        memory[29794] <=  8'h61;        memory[29795] <=  8'h72;        memory[29796] <=  8'h74;        memory[29797] <=  8'h74;        memory[29798] <=  8'h62;        memory[29799] <=  8'h61;        memory[29800] <=  8'h72;        memory[29801] <=  8'h74;        memory[29802] <=  8'h78;        memory[29803] <=  8'h61;        memory[29804] <=  8'h74;        memory[29805] <=  8'h6b;        memory[29806] <=  8'h73;        memory[29807] <=  8'h68;        memory[29808] <=  8'h63;        memory[29809] <=  8'h66;        memory[29810] <=  8'h69;        memory[29811] <=  8'h77;        memory[29812] <=  8'h68;        memory[29813] <=  8'h61;        memory[29814] <=  8'h74;        memory[29815] <=  8'h61;        memory[29816] <=  8'h6e;        memory[29817] <=  8'h61;        memory[29818] <=  8'h62;        memory[29819] <=  8'h61;        memory[29820] <=  8'h63;        memory[29821] <=  8'h61;        memory[29822] <=  8'h74;        memory[29823] <=  8'h61;        memory[29824] <=  8'h62;        memory[29825] <=  8'h61;        memory[29826] <=  8'h72;        memory[29827] <=  8'h63;        memory[29828] <=  8'h61;        memory[29829] <=  8'h68;        memory[29830] <=  8'h64;        memory[29831] <=  8'h75;        memory[29832] <=  8'h63;        memory[29833] <=  8'h74;        memory[29834] <=  8'h61;        memory[29835] <=  8'h64;        memory[29836] <=  8'h61;        memory[29837] <=  8'h61;        memory[29838] <=  8'h63;        memory[29839] <=  8'h61;        memory[29840] <=  8'h72;        memory[29841] <=  8'h63;        memory[29842] <=  8'h74;        memory[29843] <=  8'h72;        memory[29844] <=  8'h63;        memory[29845] <=  8'h61;        memory[29846] <=  8'h74;        memory[29847] <=  8'h72;        memory[29848] <=  8'h63;        memory[29849] <=  8'h61;        memory[29850] <=  8'h74;        memory[29851] <=  8'h63;        memory[29852] <=  8'h62;        memory[29853] <=  8'h61;        memory[29854] <=  8'h74;        memory[29855] <=  8'h62;        memory[29856] <=  8'h72;        memory[29857] <=  8'h63;        memory[29858] <=  8'h61;        memory[29859] <=  8'h74;        memory[29860] <=  8'h72;        memory[29861] <=  8'h6e;        memory[29862] <=  8'h62;        memory[29863] <=  8'h61;        memory[29864] <=  8'h63;        memory[29865] <=  8'h61;        memory[29866] <=  8'h74;        memory[29867] <=  8'h79;        memory[29868] <=  8'h73;        memory[29869] <=  8'h6e;        memory[29870] <=  8'h63;        memory[29871] <=  8'h74;        memory[29872] <=  8'h61;        memory[29873] <=  8'h6e;        memory[29874] <=  8'h62;        memory[29875] <=  8'h61;        memory[29876] <=  8'h63;        memory[29877] <=  8'h72;        memory[29878] <=  8'h6e;        memory[29879] <=  8'h74;        memory[29880] <=  8'h61;        memory[29881] <=  8'h62;        memory[29882] <=  8'h74;        memory[29883] <=  8'h6e;        memory[29884] <=  8'h61;        memory[29885] <=  8'h72;        memory[29886] <=  8'h62;        memory[29887] <=  8'h78;        memory[29888] <=  8'h74;        memory[29889] <=  8'h61;        memory[29890] <=  8'h72;        memory[29891] <=  8'h62;        memory[29892] <=  8'h61;        memory[29893] <=  8'h72;        memory[29894] <=  8'h74;        memory[29895] <=  8'h74;        memory[29896] <=  8'h62;        memory[29897] <=  8'h61;        memory[29898] <=  8'h72;        memory[29899] <=  8'h74;        memory[29900] <=  8'h78;        memory[29901] <=  8'h61;        memory[29902] <=  8'h74;        memory[29903] <=  8'h6b;        memory[29904] <=  8'h73;        memory[29905] <=  8'h68;        memory[29906] <=  8'h63;        memory[29907] <=  8'h66;        memory[29908] <=  8'h69;        memory[29909] <=  8'h77;        memory[29910] <=  8'h68;        memory[29911] <=  8'h61;        memory[29912] <=  8'h74;        memory[29913] <=  8'h61;        memory[29914] <=  8'h6e;        memory[29915] <=  8'h61;        memory[29916] <=  8'h62;        memory[29917] <=  8'h61;        memory[29918] <=  8'h63;        memory[29919] <=  8'h61;        memory[29920] <=  8'h74;        memory[29921] <=  8'h61;        memory[29922] <=  8'h62;        memory[29923] <=  8'h61;        memory[29924] <=  8'h72;        memory[29925] <=  8'h63;        memory[29926] <=  8'h61;        memory[29927] <=  8'h68;        memory[29928] <=  8'h64;        memory[29929] <=  8'h75;        memory[29930] <=  8'h63;        memory[29931] <=  8'h74;        memory[29932] <=  8'h61;        memory[29933] <=  8'h64;        memory[29934] <=  8'h61;        memory[29935] <=  8'h61;        memory[29936] <=  8'h63;        memory[29937] <=  8'h61;        memory[29938] <=  8'h72;        memory[29939] <=  8'h63;        memory[29940] <=  8'h74;        memory[29941] <=  8'h72;        memory[29942] <=  8'h63;        memory[29943] <=  8'h61;        memory[29944] <=  8'h74;        memory[29945] <=  8'h72;        memory[29946] <=  8'h63;        memory[29947] <=  8'h61;        memory[29948] <=  8'h74;        memory[29949] <=  8'h63;        memory[29950] <=  8'h62;        memory[29951] <=  8'h61;        memory[29952] <=  8'h74;        memory[29953] <=  8'h62;        memory[29954] <=  8'h72;        memory[29955] <=  8'h63;        memory[29956] <=  8'h61;        memory[29957] <=  8'h74;        memory[29958] <=  8'h72;        memory[29959] <=  8'h6e;        memory[29960] <=  8'h62;        memory[29961] <=  8'h61;        memory[29962] <=  8'h63;        memory[29963] <=  8'h61;        memory[29964] <=  8'h74;        memory[29965] <=  8'h79;        memory[29966] <=  8'h73;        memory[29967] <=  8'h6e;        memory[29968] <=  8'h63;        memory[29969] <=  8'h74;        memory[29970] <=  8'h61;        memory[29971] <=  8'h6e;        memory[29972] <=  8'h62;        memory[29973] <=  8'h61;        memory[29974] <=  8'h63;        memory[29975] <=  8'h72;        memory[29976] <=  8'h6e;        memory[29977] <=  8'h74;        memory[29978] <=  8'h61;        memory[29979] <=  8'h62;        memory[29980] <=  8'h74;        memory[29981] <=  8'h6e;        memory[29982] <=  8'h61;        memory[29983] <=  8'h72;        memory[29984] <=  8'h62;        memory[29985] <=  8'h78;        memory[29986] <=  8'h74;        memory[29987] <=  8'h61;        memory[29988] <=  8'h72;        memory[29989] <=  8'h64;        memory[29990] <=  8'h66;        memory[29991] <=  8'h73;        memory[29992] <=  8'h67;        memory[29993] <=  8'h76;        memory[29994] <=  8'h68;        memory[29995] <=  8'h62;        memory[29996] <=  8'h6b;        memory[29997] <=  8'h6a;        memory[29998] <=  8'h6e;        memory[29999] <=  8'h6d;        memory[30000] <=  8'h62;        memory[30001] <=  8'h76;        memory[30002] <=  8'h78;        memory[30003] <=  8'h63;        memory[30004] <=  8'h73;        memory[30005] <=  8'h66;        memory[30006] <=  8'h72;        memory[30007] <=  8'h74;        memory[30008] <=  8'h79;        memory[30009] <=  8'h75;        memory[30010] <=  8'h6a;        memory[30011] <=  8'h6e;        memory[30012] <=  8'h62;        memory[30013] <=  8'h76;        memory[30014] <=  8'h63;        memory[30015] <=  8'h64;        memory[30016] <=  8'h74;        memory[30017] <=  8'h79;        memory[30018] <=  8'h75;        memory[30019] <=  8'h69;        memory[30020] <=  8'h6b;        memory[30021] <=  8'h6d;        memory[30022] <=  8'h6e;        memory[30023] <=  8'h62;        memory[30024] <=  8'h76;        memory[30025] <=  8'h63;        memory[30026] <=  8'h78;        memory[30027] <=  8'h73;        memory[30028] <=  8'h64;        memory[30029] <=  8'h72;        memory[30030] <=  8'h74;        memory[30031] <=  8'h79;        memory[30032] <=  8'h75;        memory[30033] <=  8'h69;        memory[30034] <=  8'h6b;        memory[30035] <=  8'h6d;        memory[30036] <=  8'h6e;        memory[30037] <=  8'h62;        memory[30038] <=  8'h76;        memory[30039] <=  8'h63;        memory[30040] <=  8'h73;        memory[30041] <=  8'h77;        memory[30042] <=  8'h33;        memory[30043] <=  8'h34;        memory[30044] <=  8'h35;        memory[30045] <=  8'h36;        memory[30046] <=  8'h37;        memory[30047] <=  8'h38;        memory[30048] <=  8'h69;        memory[30049] <=  8'h6b;        memory[30050] <=  8'h6d;        memory[30051] <=  8'h6e;        memory[30052] <=  8'h62;        memory[30053] <=  8'h76;        memory[30054] <=  8'h63;        memory[30055] <=  8'h64;        memory[30056] <=  8'h65;        memory[30057] <=  8'h72;        memory[30058] <=  8'h36;        memory[30059] <=  8'h37;        memory[30060] <=  8'h38;        memory[30061] <=  8'h69;        memory[30062] <=  8'h6f;        memory[30063] <=  8'h6b;        memory[30064] <=  8'h6a;        memory[30065] <=  8'h6e;        memory[30066] <=  8'h62;        memory[30067] <=  8'h76;        memory[30068] <=  8'h63;        memory[30069] <=  8'h64;        memory[30070] <=  8'h72;        memory[30071] <=  8'h74;        memory[30072] <=  8'h79;        memory[30073] <=  8'h75;        memory[30074] <=  8'h73;        memory[30075] <=  8'h6a;        memory[30076] <=  8'h63;        memory[30077] <=  8'h6e;        memory[30078] <=  8'h62;        memory[30079] <=  8'h64;        memory[30080] <=  8'h66;        memory[30081] <=  8'h73;        memory[30082] <=  8'h74;        memory[30083] <=  8'h79;        memory[30084] <=  8'h75;        memory[30085] <=  8'h61;        memory[30086] <=  8'h69;        memory[30087] <=  8'h6b;        memory[30088] <=  8'h78;        memory[30089] <=  8'h6d;        memory[30090] <=  8'h6e;        memory[30091] <=  8'h73;        memory[30092] <=  8'h6a;        memory[30093] <=  8'h6f;        memory[30094] <=  8'h64;        memory[30095] <=  8'h6c;        memory[30096] <=  8'h63;        memory[30097] <=  8'h78;        memory[30098] <=  8'h62;        memory[30099] <=  8'h61;        memory[30100] <=  8'h72;        memory[30101] <=  8'h74;        memory[30102] <=  8'h78;        memory[30103] <=  8'h61;        memory[30104] <=  8'h74;        memory[30105] <=  8'h6b;        memory[30106] <=  8'h73;        memory[30107] <=  8'h68;        memory[30108] <=  8'h63;        memory[30109] <=  8'h66;        memory[30110] <=  8'h69;        memory[30111] <=  8'h77;        memory[30112] <=  8'h68;        memory[30113] <=  8'h61;        memory[30114] <=  8'h74;        memory[30115] <=  8'h61;        memory[30116] <=  8'h6e;        memory[30117] <=  8'h61;        memory[30118] <=  8'h62;        memory[30119] <=  8'h61;        memory[30120] <=  8'h63;        memory[30121] <=  8'h61;        memory[30122] <=  8'h74;        memory[30123] <=  8'h61;        memory[30124] <=  8'h62;        memory[30125] <=  8'h61;        memory[30126] <=  8'h72;        memory[30127] <=  8'h63;        memory[30128] <=  8'h61;        memory[30129] <=  8'h68;        memory[30130] <=  8'h64;        memory[30131] <=  8'h75;        memory[30132] <=  8'h63;        memory[30133] <=  8'h74;        memory[30134] <=  8'h61;        memory[30135] <=  8'h64;        memory[30136] <=  8'h61;        memory[30137] <=  8'h61;        memory[30138] <=  8'h63;        memory[30139] <=  8'h61;        memory[30140] <=  8'h72;        memory[30141] <=  8'h62;        memory[30142] <=  8'h61;        memory[30143] <=  8'h72;        memory[30144] <=  8'h74;        memory[30145] <=  8'h78;        memory[30146] <=  8'h61;        memory[30147] <=  8'h74;        memory[30148] <=  8'h6b;        memory[30149] <=  8'h73;        memory[30150] <=  8'h68;        memory[30151] <=  8'h63;        memory[30152] <=  8'h66;        memory[30153] <=  8'h69;        memory[30154] <=  8'h77;        memory[30155] <=  8'h68;        memory[30156] <=  8'h61;        memory[30157] <=  8'h74;        memory[30158] <=  8'h61;        memory[30159] <=  8'h6e;        memory[30160] <=  8'h61;        memory[30161] <=  8'h62;        memory[30162] <=  8'h61;        memory[30163] <=  8'h63;        memory[30164] <=  8'h61;        memory[30165] <=  8'h74;        memory[30166] <=  8'h61;        memory[30167] <=  8'h62;        memory[30168] <=  8'h61;        memory[30169] <=  8'h72;        memory[30170] <=  8'h63;        memory[30171] <=  8'h61;        memory[30172] <=  8'h68;        memory[30173] <=  8'h64;        memory[30174] <=  8'h75;        memory[30175] <=  8'h63;        memory[30176] <=  8'h74;        memory[30177] <=  8'h61;        memory[30178] <=  8'h64;        memory[30179] <=  8'h61;        memory[30180] <=  8'h61;        memory[30181] <=  8'h63;        memory[30182] <=  8'h61;        memory[30183] <=  8'h72;        memory[30184] <=  8'h62;        memory[30185] <=  8'h61;        memory[30186] <=  8'h72;        memory[30187] <=  8'h74;        memory[30188] <=  8'h78;        memory[30189] <=  8'h61;        memory[30190] <=  8'h74;        memory[30191] <=  8'h6b;        memory[30192] <=  8'h73;        memory[30193] <=  8'h68;        memory[30194] <=  8'h63;        memory[30195] <=  8'h66;        memory[30196] <=  8'h69;        memory[30197] <=  8'h77;        memory[30198] <=  8'h68;        memory[30199] <=  8'h61;        memory[30200] <=  8'h74;        memory[30201] <=  8'h61;        memory[30202] <=  8'h6e;        memory[30203] <=  8'h61;        memory[30204] <=  8'h62;        memory[30205] <=  8'h61;        memory[30206] <=  8'h63;        memory[30207] <=  8'h61;        memory[30208] <=  8'h74;        memory[30209] <=  8'h61;        memory[30210] <=  8'h62;        memory[30211] <=  8'h61;        memory[30212] <=  8'h72;        memory[30213] <=  8'h63;        memory[30214] <=  8'h61;        memory[30215] <=  8'h68;        memory[30216] <=  8'h64;        memory[30217] <=  8'h75;        memory[30218] <=  8'h63;        memory[30219] <=  8'h74;        memory[30220] <=  8'h61;        memory[30221] <=  8'h64;        memory[30222] <=  8'h61;        memory[30223] <=  8'h61;        memory[30224] <=  8'h63;        memory[30225] <=  8'h61;        memory[30226] <=  8'h72;        memory[30227] <=  8'h62;        memory[30228] <=  8'h61;        memory[30229] <=  8'h72;        memory[30230] <=  8'h74;        memory[30231] <=  8'h78;        memory[30232] <=  8'h61;        memory[30233] <=  8'h74;        memory[30234] <=  8'h6b;        memory[30235] <=  8'h73;        memory[30236] <=  8'h68;        memory[30237] <=  8'h63;        memory[30238] <=  8'h66;        memory[30239] <=  8'h69;        memory[30240] <=  8'h77;        memory[30241] <=  8'h68;        memory[30242] <=  8'h61;        memory[30243] <=  8'h74;        memory[30244] <=  8'h61;        memory[30245] <=  8'h6e;        memory[30246] <=  8'h61;        memory[30247] <=  8'h62;        memory[30248] <=  8'h61;        memory[30249] <=  8'h63;        memory[30250] <=  8'h61;        memory[30251] <=  8'h74;        memory[30252] <=  8'h61;        memory[30253] <=  8'h62;        memory[30254] <=  8'h61;        memory[30255] <=  8'h72;        memory[30256] <=  8'h63;        memory[30257] <=  8'h61;        memory[30258] <=  8'h68;        memory[30259] <=  8'h64;        memory[30260] <=  8'h75;        memory[30261] <=  8'h63;        memory[30262] <=  8'h74;        memory[30263] <=  8'h61;        memory[30264] <=  8'h64;        memory[30265] <=  8'h61;        memory[30266] <=  8'h61;        memory[30267] <=  8'h63;        memory[30268] <=  8'h61;        memory[30269] <=  8'h72;        memory[30270] <=  8'h62;        memory[30271] <=  8'h61;        memory[30272] <=  8'h72;        memory[30273] <=  8'h74;        memory[30274] <=  8'h78;        memory[30275] <=  8'h61;        memory[30276] <=  8'h74;        memory[30277] <=  8'h6b;        memory[30278] <=  8'h73;        memory[30279] <=  8'h68;        memory[30280] <=  8'h63;        memory[30281] <=  8'h66;        memory[30282] <=  8'h69;        memory[30283] <=  8'h77;        memory[30284] <=  8'h68;        memory[30285] <=  8'h61;        memory[30286] <=  8'h74;        memory[30287] <=  8'h61;        memory[30288] <=  8'h6e;        memory[30289] <=  8'h61;        memory[30290] <=  8'h62;        memory[30291] <=  8'h61;        memory[30292] <=  8'h63;        memory[30293] <=  8'h61;        memory[30294] <=  8'h74;        memory[30295] <=  8'h61;        memory[30296] <=  8'h62;        memory[30297] <=  8'h61;        memory[30298] <=  8'h72;        memory[30299] <=  8'h63;        memory[30300] <=  8'h61;        memory[30301] <=  8'h68;        memory[30302] <=  8'h64;        memory[30303] <=  8'h75;        memory[30304] <=  8'h63;        memory[30305] <=  8'h74;        memory[30306] <=  8'h61;        memory[30307] <=  8'h64;        memory[30308] <=  8'h61;        memory[30309] <=  8'h61;        memory[30310] <=  8'h63;        memory[30311] <=  8'h61;        memory[30312] <=  8'h72;        memory[30313] <=  8'h62;        memory[30314] <=  8'h61;        memory[30315] <=  8'h72;        memory[30316] <=  8'h74;        memory[30317] <=  8'h78;        memory[30318] <=  8'h61;        memory[30319] <=  8'h74;        memory[30320] <=  8'h6b;        memory[30321] <=  8'h73;        memory[30322] <=  8'h68;        memory[30323] <=  8'h63;        memory[30324] <=  8'h66;        memory[30325] <=  8'h69;        memory[30326] <=  8'h77;        memory[30327] <=  8'h68;        memory[30328] <=  8'h61;        memory[30329] <=  8'h74;        memory[30330] <=  8'h61;        memory[30331] <=  8'h6e;        memory[30332] <=  8'h61;        memory[30333] <=  8'h62;        memory[30334] <=  8'h61;        memory[30335] <=  8'h63;        memory[30336] <=  8'h61;        memory[30337] <=  8'h74;        memory[30338] <=  8'h61;        memory[30339] <=  8'h62;        memory[30340] <=  8'h61;        memory[30341] <=  8'h72;        memory[30342] <=  8'h63;        memory[30343] <=  8'h61;        memory[30344] <=  8'h68;        memory[30345] <=  8'h64;        memory[30346] <=  8'h75;        memory[30347] <=  8'h63;        memory[30348] <=  8'h74;        memory[30349] <=  8'h61;        memory[30350] <=  8'h64;        memory[30351] <=  8'h61;        memory[30352] <=  8'h61;        memory[30353] <=  8'h63;        memory[30354] <=  8'h61;        memory[30355] <=  8'h72;        memory[30356] <=  8'h62;        memory[30357] <=  8'h61;        memory[30358] <=  8'h72;        memory[30359] <=  8'h74;        memory[30360] <=  8'h78;        memory[30361] <=  8'h61;        memory[30362] <=  8'h74;        memory[30363] <=  8'h6b;        memory[30364] <=  8'h73;        memory[30365] <=  8'h68;        memory[30366] <=  8'h63;        memory[30367] <=  8'h66;        memory[30368] <=  8'h69;        memory[30369] <=  8'h77;        memory[30370] <=  8'h68;        memory[30371] <=  8'h61;        memory[30372] <=  8'h74;        memory[30373] <=  8'h61;        memory[30374] <=  8'h6e;        memory[30375] <=  8'h61;        memory[30376] <=  8'h62;        memory[30377] <=  8'h61;        memory[30378] <=  8'h63;        memory[30379] <=  8'h61;        memory[30380] <=  8'h74;        memory[30381] <=  8'h61;        memory[30382] <=  8'h62;        memory[30383] <=  8'h61;        memory[30384] <=  8'h72;        memory[30385] <=  8'h63;        memory[30386] <=  8'h61;        memory[30387] <=  8'h68;        memory[30388] <=  8'h64;        memory[30389] <=  8'h75;        memory[30390] <=  8'h63;        memory[30391] <=  8'h74;        memory[30392] <=  8'h61;        memory[30393] <=  8'h64;        memory[30394] <=  8'h61;        memory[30395] <=  8'h61;        memory[30396] <=  8'h63;        memory[30397] <=  8'h61;        memory[30398] <=  8'h72;        memory[30399] <=  8'h62;        memory[30400] <=  8'h61;        memory[30401] <=  8'h72;        memory[30402] <=  8'h74;        memory[30403] <=  8'h78;        memory[30404] <=  8'h61;        memory[30405] <=  8'h74;        memory[30406] <=  8'h6b;        memory[30407] <=  8'h73;        memory[30408] <=  8'h68;        memory[30409] <=  8'h63;        memory[30410] <=  8'h66;        memory[30411] <=  8'h69;        memory[30412] <=  8'h77;        memory[30413] <=  8'h68;        memory[30414] <=  8'h61;        memory[30415] <=  8'h74;        memory[30416] <=  8'h61;        memory[30417] <=  8'h6e;        memory[30418] <=  8'h61;        memory[30419] <=  8'h62;        memory[30420] <=  8'h61;        memory[30421] <=  8'h63;        memory[30422] <=  8'h61;        memory[30423] <=  8'h74;        memory[30424] <=  8'h61;        memory[30425] <=  8'h62;        memory[30426] <=  8'h61;        memory[30427] <=  8'h72;        memory[30428] <=  8'h63;        memory[30429] <=  8'h61;        memory[30430] <=  8'h68;        memory[30431] <=  8'h64;        memory[30432] <=  8'h75;        memory[30433] <=  8'h63;        memory[30434] <=  8'h74;        memory[30435] <=  8'h61;        memory[30436] <=  8'h64;        memory[30437] <=  8'h61;        memory[30438] <=  8'h61;        memory[30439] <=  8'h63;        memory[30440] <=  8'h61;        memory[30441] <=  8'h72;        memory[30442] <=  8'h62;        memory[30443] <=  8'h61;        memory[30444] <=  8'h72;        memory[30445] <=  8'h74;        memory[30446] <=  8'h78;        memory[30447] <=  8'h61;        memory[30448] <=  8'h74;        memory[30449] <=  8'h6b;        memory[30450] <=  8'h73;        memory[30451] <=  8'h68;        memory[30452] <=  8'h63;        memory[30453] <=  8'h66;        memory[30454] <=  8'h69;        memory[30455] <=  8'h77;        memory[30456] <=  8'h68;        memory[30457] <=  8'h61;        memory[30458] <=  8'h74;        memory[30459] <=  8'h61;        memory[30460] <=  8'h6e;        memory[30461] <=  8'h61;        memory[30462] <=  8'h62;        memory[30463] <=  8'h61;        memory[30464] <=  8'h63;        memory[30465] <=  8'h61;        memory[30466] <=  8'h74;        memory[30467] <=  8'h61;        memory[30468] <=  8'h62;        memory[30469] <=  8'h61;        memory[30470] <=  8'h72;        memory[30471] <=  8'h63;        memory[30472] <=  8'h61;        memory[30473] <=  8'h68;        memory[30474] <=  8'h64;        memory[30475] <=  8'h75;        memory[30476] <=  8'h63;        memory[30477] <=  8'h74;        memory[30478] <=  8'h61;        memory[30479] <=  8'h64;        memory[30480] <=  8'h61;        memory[30481] <=  8'h61;        memory[30482] <=  8'h63;        memory[30483] <=  8'h61;        memory[30484] <=  8'h72;        memory[30485] <=  8'h62;        memory[30486] <=  8'h61;        memory[30487] <=  8'h72;        memory[30488] <=  8'h74;        memory[30489] <=  8'h74;        memory[30490] <=  8'h62;        memory[30491] <=  8'h61;        memory[30492] <=  8'h72;        memory[30493] <=  8'h74;        memory[30494] <=  8'h78;        memory[30495] <=  8'h61;        memory[30496] <=  8'h74;        memory[30497] <=  8'h6b;        memory[30498] <=  8'h73;        memory[30499] <=  8'h68;        memory[30500] <=  8'h63;        memory[30501] <=  8'h66;        memory[30502] <=  8'h69;        memory[30503] <=  8'h77;        memory[30504] <=  8'h68;        memory[30505] <=  8'h61;        memory[30506] <=  8'h74;        memory[30507] <=  8'h61;        memory[30508] <=  8'h6e;        memory[30509] <=  8'h61;        memory[30510] <=  8'h62;        memory[30511] <=  8'h61;        memory[30512] <=  8'h63;        memory[30513] <=  8'h61;        memory[30514] <=  8'h74;        memory[30515] <=  8'h61;        memory[30516] <=  8'h62;        memory[30517] <=  8'h61;        memory[30518] <=  8'h72;        memory[30519] <=  8'h63;        memory[30520] <=  8'h61;        memory[30521] <=  8'h68;        memory[30522] <=  8'h64;        memory[30523] <=  8'h75;        memory[30524] <=  8'h63;        memory[30525] <=  8'h74;        memory[30526] <=  8'h61;        memory[30527] <=  8'h64;        memory[30528] <=  8'h61;        memory[30529] <=  8'h61;        memory[30530] <=  8'h63;        memory[30531] <=  8'h61;        memory[30532] <=  8'h72;        memory[30533] <=  8'h63;        memory[30534] <=  8'h74;        memory[30535] <=  8'h72;        memory[30536] <=  8'h63;        memory[30537] <=  8'h61;        memory[30538] <=  8'h74;        memory[30539] <=  8'h72;        memory[30540] <=  8'h63;        memory[30541] <=  8'h61;        memory[30542] <=  8'h74;        memory[30543] <=  8'h63;        memory[30544] <=  8'h62;        memory[30545] <=  8'h61;        memory[30546] <=  8'h74;        memory[30547] <=  8'h62;        memory[30548] <=  8'h72;        memory[30549] <=  8'h63;        memory[30550] <=  8'h61;        memory[30551] <=  8'h72;        memory[30552] <=  8'h62;        memory[30553] <=  8'h78;        memory[30554] <=  8'h74;        memory[30555] <=  8'h61;        memory[30556] <=  8'h72;        memory[30557] <=  8'h64;        memory[30558] <=  8'h66;        memory[30559] <=  8'h73;        memory[30560] <=  8'h67;        memory[30561] <=  8'h76;        memory[30562] <=  8'h68;        memory[30563] <=  8'h62;        memory[30564] <=  8'h6b;        memory[30565] <=  8'h6a;        memory[30566] <=  8'h6e;        memory[30567] <=  8'h6d;        memory[30568] <=  8'h62;        memory[30569] <=  8'h76;        memory[30570] <=  8'h78;        memory[30571] <=  8'h63;        memory[30572] <=  8'h73;        memory[30573] <=  8'h66;        memory[30574] <=  8'h72;        memory[30575] <=  8'h74;        memory[30576] <=  8'h79;        memory[30577] <=  8'h75;        memory[30578] <=  8'h6a;        memory[30579] <=  8'h6e;        memory[30580] <=  8'h62;        memory[30581] <=  8'h76;        memory[30582] <=  8'h63;        memory[30583] <=  8'h64;        memory[30584] <=  8'h74;        memory[30585] <=  8'h79;        memory[30586] <=  8'h75;        memory[30587] <=  8'h69;        memory[30588] <=  8'h6b;        memory[30589] <=  8'h6d;        memory[30590] <=  8'h6e;        memory[30591] <=  8'h62;        memory[30592] <=  8'h76;        memory[30593] <=  8'h63;        memory[30594] <=  8'h78;        memory[30595] <=  8'h73;        memory[30596] <=  8'h64;        memory[30597] <=  8'h72;        memory[30598] <=  8'h74;        memory[30599] <=  8'h79;        memory[30600] <=  8'h75;        memory[30601] <=  8'h69;        memory[30602] <=  8'h6b;        memory[30603] <=  8'h6d;        memory[30604] <=  8'h6e;        memory[30605] <=  8'h62;        memory[30606] <=  8'h76;        memory[30607] <=  8'h63;        memory[30608] <=  8'h73;        memory[30609] <=  8'h77;        memory[30610] <=  8'h33;        memory[30611] <=  8'h34;        memory[30612] <=  8'h35;        memory[30613] <=  8'h36;        memory[30614] <=  8'h37;        memory[30615] <=  8'h38;        memory[30616] <=  8'h69;        memory[30617] <=  8'h6b;        memory[30618] <=  8'h6d;        memory[30619] <=  8'h6e;        memory[30620] <=  8'h62;        memory[30621] <=  8'h76;        memory[30622] <=  8'h63;        memory[30623] <=  8'h64;        memory[30624] <=  8'h65;        memory[30625] <=  8'h72;        memory[30626] <=  8'h36;        memory[30627] <=  8'h37;        memory[30628] <=  8'h38;        memory[30629] <=  8'h69;        memory[30630] <=  8'h6f;        memory[30631] <=  8'h6b;        memory[30632] <=  8'h6a;        memory[30633] <=  8'h6e;        memory[30634] <=  8'h62;        memory[30635] <=  8'h76;        memory[30636] <=  8'h63;        memory[30637] <=  8'h64;        memory[30638] <=  8'h72;        memory[30639] <=  8'h74;        memory[30640] <=  8'h79;        memory[30641] <=  8'h75;        memory[30642] <=  8'h73;        memory[30643] <=  8'h6a;        memory[30644] <=  8'h63;        memory[30645] <=  8'h6e;        memory[30646] <=  8'h62;        memory[30647] <=  8'h64;        memory[30648] <=  8'h66;        memory[30649] <=  8'h73;        memory[30650] <=  8'h74;        memory[30651] <=  8'h79;        memory[30652] <=  8'h75;        memory[30653] <=  8'h61;        memory[30654] <=  8'h69;        memory[30655] <=  8'h6b;        memory[30656] <=  8'h78;        memory[30657] <=  8'h6d;        memory[30658] <=  8'h6e;        memory[30659] <=  8'h73;        memory[30660] <=  8'h6a;        memory[30661] <=  8'h6f;        memory[30662] <=  8'h64;        memory[30663] <=  8'h6c;        memory[30664] <=  8'h63;        memory[30665] <=  8'h78;        memory[30666] <=  8'h2c;        memory[30667] <=  8'h6d;        memory[30668] <=  8'h73;        memory[30669] <=  8'h6b;        memory[30670] <=  8'h64;        memory[30671] <=  8'h6c;        memory[30672] <=  8'h70;        memory[30673] <=  8'h5b;        memory[30674] <=  8'h3b;        memory[30675] <=  8'h73;        memory[30676] <=  8'h6c;        memory[30677] <=  8'h64;        memory[30678] <=  8'h70;        memory[30679] <=  8'h76;        memory[30680] <=  8'h63;        memory[30681] <=  8'h5b;        memory[30682] <=  8'h78;        memory[30683] <=  8'h76;        memory[30684] <=  8'h63;        memory[30685] <=  8'h5b;        memory[30686] <=  8'h78;        memory[30687] <=  8'h70;        memory[30688] <=  8'h6f;        memory[30689] <=  8'h20;        memory[30690] <=  8'h62;        memory[30691] <=  8'h61;        memory[30692] <=  8'h72;        memory[30693] <=  8'h74;        memory[30694] <=  8'h74;        memory[30695] <=  8'h62;        memory[30696] <=  8'h61;        memory[30697] <=  8'h72;        memory[30698] <=  8'h74;        memory[30699] <=  8'h78;        memory[30700] <=  8'h61;        memory[30701] <=  8'h74;        memory[30702] <=  8'h6b;        memory[30703] <=  8'h73;        memory[30704] <=  8'h68;        memory[30705] <=  8'h63;        memory[30706] <=  8'h66;        memory[30707] <=  8'h69;        memory[30708] <=  8'h77;        memory[30709] <=  8'h68;        memory[30710] <=  8'h61;        memory[30711] <=  8'h69;        memory[30712] <=  8'h6a;        memory[30713] <=  8'h78;        memory[30714] <=  8'h5d;        memory[30715] <=  8'h65;        memory[30716] <=  8'h6b;        memory[30717] <=  8'h6f;        memory[30718] <=  8'h39;        memory[30719] <=  8'h64;        memory[30720] <=  8'h75;        memory[30721] <=  8'h38;        memory[30722] <=  8'h79;        memory[30723] <=  8'h20;        memory[30724] <=  8'h37;        memory[30725] <=  8'h63;        memory[30726] <=  8'h67;        memory[30727] <=  8'h78;        memory[30728] <=  8'h63;        memory[30729] <=  8'h75;        memory[30730] <=  8'h68;        memory[30731] <=  8'h69;        memory[30732] <=  8'h6a;        memory[30733] <=  8'h77;        memory[30734] <=  8'h69;        memory[30735] <=  8'h64;        memory[30736] <=  8'h66;        memory[30737] <=  8'h68;        memory[30738] <=  8'h75;        memory[30739] <=  8'h76;        memory[30740] <=  8'h64;        memory[30741] <=  8'h62;        memory[30742] <=  8'h66;        memory[30743] <=  8'h6a;        memory[30744] <=  8'h6e;        memory[30745] <=  8'h6b;        memory[30746] <=  8'h6a;        memory[30747] <=  8'h65;        memory[30748] <=  8'h38;        memory[30749] <=  8'h66;        memory[30750] <=  8'h37;        memory[30751] <=  8'h67;        memory[30752] <=  8'h79;        memory[30753] <=  8'h76;        memory[30754] <=  8'h63;        memory[30755] <=  8'h68;        memory[30756] <=  8'h69;        memory[30757] <=  8'h6a;        memory[30758] <=  8'h33;        memory[30759] <=  8'h65;        memory[30760] <=  8'h67;        memory[30761] <=  8'h79;        memory[30762] <=  8'h72;        memory[30763] <=  8'h64;        memory[30764] <=  8'h62;        memory[30765] <=  8'h6e;        memory[30766] <=  8'h63;        memory[30767] <=  8'h7a;        memory[30768] <=  8'h6a;        memory[30769] <=  8'h6f;        memory[30770] <=  8'h66;        memory[30771] <=  8'h78;        memory[30772] <=  8'h6a;        memory[30773] <=  8'h69;        memory[30774] <=  8'h63;        memory[30775] <=  8'h68;        memory[30776] <=  8'h62;        memory[30777] <=  8'h6e;        memory[30778] <=  8'h6d;        memory[30779] <=  8'h63;        memory[30780] <=  8'h73;        memory[30781] <=  8'h6c;        memory[30782] <=  8'h6b;        memory[30783] <=  8'h6a;        memory[30784] <=  8'h69;        memory[30785] <=  8'h68;        memory[30786] <=  8'h76;        memory[30787] <=  8'h75;        memory[30788] <=  8'h69;        memory[30789] <=  8'h64;        memory[30790] <=  8'h68;        memory[30791] <=  8'h75;        memory[30792] <=  8'h67;        memory[30793] <=  8'h79;        memory[30794] <=  8'h62;        memory[30795] <=  8'h68;        memory[30796] <=  8'h65;        memory[30797] <=  8'h6a;        memory[30798] <=  8'h72;        memory[30799] <=  8'h6b;        memory[30800] <=  8'h6a;        memory[30801] <=  8'h6f;        memory[30802] <=  8'h64;        memory[30803] <=  8'h67;        memory[30804] <=  8'h69;        memory[30805] <=  8'h75;        memory[30806] <=  8'h69;        memory[30807] <=  8'h67;        memory[30808] <=  8'h76;        memory[30809] <=  8'h79;        memory[30810] <=  8'h75;        memory[30811] <=  8'h67;        memory[30812] <=  8'h78;        memory[30813] <=  8'h68;        memory[30814] <=  8'h63;        memory[30815] <=  8'h20;        memory[30816] <=  8'h20;        memory[30817] <=  8'h20;        memory[30818] <=  8'h78;        memory[30819] <=  8'h76;        memory[30820] <=  8'h20;        memory[30821] <=  8'h63;        memory[30822] <=  8'h78;        memory[30823] <=  8'h67;        memory[30824] <=  8'h79;        memory[30825] <=  8'h63;        memory[30826] <=  8'h75;        memory[30827] <=  8'h68;        memory[30828] <=  8'h6a;        memory[30829] <=  8'h6b;        memory[30830] <=  8'h61;        memory[30831] <=  8'h6c;        memory[30832] <=  8'h78;        memory[30833] <=  8'h76;        memory[30834] <=  8'h70;        memory[30835] <=  8'h6f;        memory[30836] <=  8'h69;        memory[30837] <=  8'h6a;        memory[30838] <=  8'h69;        memory[30839] <=  8'h68;        memory[30840] <=  8'h6a;        memory[30841] <=  8'h62;        memory[30842] <=  8'h77;        memory[30843] <=  8'h65;        memory[30844] <=  8'h6e;        memory[30845] <=  8'h61;        memory[30846] <=  8'h66;        memory[30847] <=  8'h6d;        memory[30848] <=  8'h64;        memory[30849] <=  8'h6b;        memory[30850] <=  8'h6d;        memory[30851] <=  8'h76;        memory[30852] <=  8'h6c;        memory[30853] <=  8'h63;        memory[30854] <=  8'h6f;        memory[30855] <=  8'h64;        memory[30856] <=  8'h69;        memory[30857] <=  8'h75;        memory[30858] <=  8'h68;        memory[30859] <=  8'h73;        memory[30860] <=  8'h66;        memory[30861] <=  8'h65;        memory[30862] <=  8'h62;        memory[30863] <=  8'h6e;        memory[30864] <=  8'h64;        memory[30865] <=  8'h73;        memory[30866] <=  8'h63;        memory[30867] <=  8'h6b;        memory[30868] <=  8'h20;        memory[30869] <=  8'h78;        memory[30870] <=  8'h6a;        memory[30871] <=  8'h78;        memory[30872] <=  8'h63;        memory[30873] <=  8'h73;        memory[30874] <=  8'h64;        memory[30875] <=  8'h66;        memory[30876] <=  8'h6b;        memory[30877] <=  8'h64;        memory[30878] <=  8'h6e;        memory[30879] <=  8'h6d;        memory[30880] <=  8'h64;        memory[30881] <=  8'h73;        memory[30882] <=  8'h63;        memory[30883] <=  8'h6b;        memory[30884] <=  8'h78;        memory[30885] <=  8'h6c;        memory[30886] <=  8'h6f;        memory[30887] <=  8'h66;        memory[30888] <=  8'h6a;        memory[30889] <=  8'h69;        memory[30890] <=  8'h61;        memory[30891] <=  8'h62;        memory[30892] <=  8'h6e;        memory[30893] <=  8'h20;        memory[30894] <=  8'h78;        memory[30895] <=  8'h6b;        memory[30896] <=  8'h6d;        memory[30897] <=  8'h20;        memory[30898] <=  8'h6f;        memory[30899] <=  8'h63;        memory[30900] <=  8'h76;        memory[30901] <=  8'h73;        memory[30902] <=  8'h64;        memory[30903] <=  8'h69;        memory[30904] <=  8'h66;        memory[30905] <=  8'h68;        memory[30906] <=  8'h65;        memory[30907] <=  8'h71;        memory[30908] <=  8'h6a;        memory[30909] <=  8'h77;        memory[30910] <=  8'h62;        memory[30911] <=  8'h65;        memory[30912] <=  8'h6e;        memory[30913] <=  8'h20;        memory[30914] <=  8'h6d;        memory[30915] <=  8'h64;        memory[30916] <=  8'h73;        memory[30917] <=  8'h6c;        memory[30918] <=  8'h76;        memory[30919] <=  8'h6b;        memory[30920] <=  8'h63;        memory[30921] <=  8'h78;        memory[30922] <=  8'h20;        memory[30923] <=  8'h6f;        memory[30924] <=  8'h78;        memory[30925] <=  8'h69;        memory[30926] <=  8'h63;        memory[30927] <=  8'h6a;        memory[30928] <=  8'h76;        memory[30929] <=  8'h64;        memory[30930] <=  8'h66;        memory[30931] <=  8'h65;        memory[30932] <=  8'h71;        memory[30933] <=  8'h6e;        memory[30934] <=  8'h20;        memory[30935] <=  8'h64;        memory[30936] <=  8'h6d;        memory[30937] <=  8'h73;        memory[30938] <=  8'h6c;        memory[30939] <=  8'h63;        memory[30940] <=  8'h78;        memory[30941] <=  8'h6b;        memory[30942] <=  8'h20;        memory[30943] <=  8'h6f;        memory[30944] <=  8'h78;        memory[30945] <=  8'h63;        memory[30946] <=  8'h76;        memory[30947] <=  8'h6a;        memory[30948] <=  8'h64;        memory[30949] <=  8'h62;        memory[30950] <=  8'h71;        memory[30951] <=  8'h77;        memory[30952] <=  8'h65;        memory[30953] <=  8'h6e;        memory[30954] <=  8'h6d;        memory[30955] <=  8'h64;        memory[30956] <=  8'h6c;        memory[30957] <=  8'h73;        memory[30958] <=  8'h2c;        memory[30959] <=  8'h76;        memory[30960] <=  8'h63;        memory[30961] <=  8'h78;        memory[30962] <=  8'h20;        memory[30963] <=  8'h63;        memory[30964] <=  8'h6f;        memory[30965] <=  8'h69;        memory[30966] <=  8'h76;        memory[30967] <=  8'h68;        memory[30968] <=  8'h73;        memory[30969] <=  8'h64;        memory[30970] <=  8'h62;        memory[30971] <=  8'h71;        memory[30972] <=  8'h77;        memory[30973] <=  8'h65;        memory[30974] <=  8'h6e;        memory[30975] <=  8'h64;        memory[30976] <=  8'h6b;        memory[30977] <=  8'h73;        memory[30978] <=  8'h76;        memory[30979] <=  8'h6f;        memory[30980] <=  8'h63;        memory[30981] <=  8'h20;        memory[30982] <=  8'h76;        memory[30983] <=  8'h69;        memory[30984] <=  8'h75;        memory[30985] <=  8'h69;        memory[30986] <=  8'h68;        memory[30987] <=  8'h63;        memory[30988] <=  8'h78;        memory[30989] <=  8'h69;        memory[30990] <=  8'h6f;        memory[30991] <=  8'h76;        memory[30992] <=  8'h73;        memory[30993] <=  8'h64;        memory[30994] <=  8'h61;        memory[30995] <=  8'h64;        memory[30996] <=  8'h6e;        memory[30997] <=  8'h77;        memory[30998] <=  8'h71;        memory[30999] <=  8'h6b;        memory[31000] <=  8'h6c;        memory[31001] <=  8'h73;        memory[31002] <=  8'h76;        memory[31003] <=  8'h6e;        memory[31004] <=  8'h62;        memory[31005] <=  8'h20;        memory[31006] <=  8'h64;        memory[31007] <=  8'h66;        memory[31008] <=  8'h6a;        memory[31009] <=  8'h6b;        memory[31010] <=  8'h71;        memory[31011] <=  8'h64;        memory[31012] <=  8'h77;        memory[31013] <=  8'h65;        memory[31014] <=  8'h6e;        memory[31015] <=  8'h62;        memory[31016] <=  8'h20;        memory[31017] <=  8'h64;        memory[31018] <=  8'h73;        memory[31019] <=  8'h76;        memory[31020] <=  8'h68;        memory[31021] <=  8'h64;        memory[31022] <=  8'h61;        memory[31023] <=  8'h71;        memory[31024] <=  8'h77;        memory[31025] <=  8'h6a;        memory[31026] <=  8'h65;        memory[31027] <=  8'h6e;        memory[31028] <=  8'h64;        memory[31029] <=  8'h20;        memory[31030] <=  8'h61;        memory[31031] <=  8'h63;        memory[31032] <=  8'h62;        memory[31033] <=  8'h68;        memory[31034] <=  8'h64;        memory[31035] <=  8'h61;        memory[31036] <=  8'h77;        memory[31037] <=  8'h71;        memory[31038] <=  8'h6e;        memory[31039] <=  8'h20;        memory[31040] <=  8'h62;        memory[31041] <=  8'h73;        memory[31042] <=  8'h76;        memory[31043] <=  8'h61;        memory[31044] <=  8'h67;        memory[31045] <=  8'h76;        memory[31046] <=  8'h68;        memory[31047] <=  8'h67;        memory[31048] <=  8'h61;        memory[31049] <=  8'h73;        memory[31050] <=  8'h6a;        memory[31051] <=  8'h6b;        memory[31052] <=  8'h63;        memory[31053] <=  8'h78;        memory[31054] <=  8'h76;        memory[31055] <=  8'h6e;        memory[31056] <=  8'h73;        memory[31057] <=  8'h64;        memory[31058] <=  8'h20;        memory[31059] <=  8'h66;        memory[31060] <=  8'h62;        memory[31061] <=  8'h64;        memory[31062] <=  8'h61;        memory[31063] <=  8'h73;        memory[31064] <=  8'h76;        memory[31065] <=  8'h67;        memory[31066] <=  8'h63;        memory[31067] <=  8'h79;        memory[31068] <=  8'h7a;        memory[31069] <=  8'h78;        memory[31070] <=  8'h79;        memory[31071] <=  8'h75;        memory[31072] <=  8'h20;        memory[31073] <=  8'h69;        memory[31074] <=  8'h6a;        memory[31075] <=  8'h64;        memory[31076] <=  8'h66;        memory[31077] <=  8'h6b;        memory[31078] <=  8'h61;        memory[31079] <=  8'h64;        memory[31080] <=  8'h63;        memory[31081] <=  8'h78;        memory[31082] <=  8'h68;        memory[31083] <=  8'h20;        memory[31084] <=  8'h67;        memory[31085] <=  8'h61;        memory[31086] <=  8'h68;        memory[31087] <=  8'h75;        memory[31088] <=  8'h64;        memory[31089] <=  8'h73;        memory[31090] <=  8'h69;        memory[31091] <=  8'h6a;        memory[31092] <=  8'h61;        memory[31093] <=  8'h6b;        memory[31094] <=  8'h63;        memory[31095] <=  8'h62;        memory[31096] <=  8'h61;        memory[31097] <=  8'h72;        memory[31098] <=  8'h73;        memory[31099] <=  8'h68;        memory[31100] <=  8'h64;        memory[31101] <=  8'h66;        memory[31102] <=  8'h67;        memory[31103] <=  8'h73;        memory[31104] <=  8'h68;        memory[31105] <=  8'h64;        memory[31106] <=  8'h66;        memory[31107] <=  8'h68;        memory[31108] <=  8'h64;        memory[31109] <=  8'h6a;        memory[31110] <=  8'h68;        memory[31111] <=  8'h62;        memory[31112] <=  8'h67;        memory[31113] <=  8'h63;        memory[31114] <=  8'h61;        memory[31115] <=  8'h66;        memory[31116] <=  8'h73;        memory[31117] <=  8'h79;        memory[31118] <=  8'h67;        memory[31119] <=  8'h6b;        memory[31120] <=  8'h75;        memory[31121] <=  8'h64;        memory[31122] <=  8'h68;        memory[31123] <=  8'h62;        memory[31124] <=  8'h77;        memory[31125] <=  8'h76;        memory[31126] <=  8'h67;        memory[31127] <=  8'h61;        memory[31128] <=  8'h66;        memory[31129] <=  8'h64;        memory[31130] <=  8'h74;        memory[31131] <=  8'h75;        memory[31132] <=  8'h66;        memory[31133] <=  8'h79;        memory[31134] <=  8'h67;        memory[31135] <=  8'h69;        memory[31136] <=  8'h75;        memory[31137] <=  8'h68;        memory[31138] <=  8'h6c;        memory[31139] <=  8'h6a;        memory[31140] <=  8'h62;        memory[31141] <=  8'h6b;        memory[31142] <=  8'h68;        memory[31143] <=  8'h76;        memory[31144] <=  8'h67;        memory[31145] <=  8'h63;        memory[31146] <=  8'h66;        memory[31147] <=  8'h78;        memory[31148] <=  8'h64;        memory[31149] <=  8'h74;        memory[31150] <=  8'h75;        memory[31151] <=  8'h79;        memory[31152] <=  8'h69;        memory[31153] <=  8'h75;        memory[31154] <=  8'h68;        memory[31155] <=  8'h6c;        memory[31156] <=  8'h6a;        memory[31157] <=  8'h6b;        memory[31158] <=  8'h67;        memory[31159] <=  8'h6a;        memory[31160] <=  8'h63;        memory[31161] <=  8'h66;        memory[31162] <=  8'h68;        memory[31163] <=  8'h64;        memory[31164] <=  8'h67;        memory[31165] <=  8'h72;        memory[31166] <=  8'h79;        memory[31167] <=  8'h74;        memory[31168] <=  8'h66;        memory[31169] <=  8'h75;        memory[31170] <=  8'h79;        memory[31171] <=  8'h69;        memory[31172] <=  8'h68;        memory[31173] <=  8'h6c;        memory[31174] <=  8'h62;        memory[31175] <=  8'h6d;        memory[31176] <=  8'h76;        memory[31177] <=  8'h6e;        memory[31178] <=  8'h63;        memory[31179] <=  8'h66;        memory[31180] <=  8'h68;        memory[31181] <=  8'h64;        memory[31182] <=  8'h74;        memory[31183] <=  8'h75;        memory[31184] <=  8'h67;        memory[31185] <=  8'h79;        memory[31186] <=  8'h69;        memory[31187] <=  8'h68;        memory[31188] <=  8'h75;        memory[31189] <=  8'h6a;        memory[31190] <=  8'h6c;        memory[31191] <=  8'h62;        memory[31192] <=  8'h6d;        memory[31193] <=  8'h76;        memory[31194] <=  8'h6e;        memory[31195] <=  8'h63;        memory[31196] <=  8'h66;        memory[31197] <=  8'h68;        memory[31198] <=  8'h67;        memory[31199] <=  8'h79;        memory[31200] <=  8'h68;        memory[31201] <=  8'h75;        memory[31202] <=  8'h6a;        memory[31203] <=  8'h6e;        memory[31204] <=  8'h2c;        memory[31205] <=  8'h62;        memory[31206] <=  8'h6e;        memory[31207] <=  8'h6d;        memory[31208] <=  8'h76;        memory[31209] <=  8'h6e;        memory[31210] <=  8'h63;        memory[31211] <=  8'h66;        memory[31212] <=  8'h68;        memory[31213] <=  8'h74;        memory[31214] <=  8'h79;        memory[31215] <=  8'h69;        memory[31216] <=  8'h75;        memory[31217] <=  8'h6c;        memory[31218] <=  8'h6a;        memory[31219] <=  8'h62;        memory[31220] <=  8'h6d;        memory[31221] <=  8'h76;        memory[31222] <=  8'h6e;        memory[31223] <=  8'h63;        memory[31224] <=  8'h66;        memory[31225] <=  8'h74;        memory[31226] <=  8'h75;        memory[31227] <=  8'h79;        memory[31228] <=  8'h69;        memory[31229] <=  8'h68;        memory[31230] <=  8'h6b;        memory[31231] <=  8'h62;        memory[31232] <=  8'h76;        memory[31233] <=  8'h63;        memory[31234] <=  8'h66;        memory[31235] <=  8'h67;        memory[31236] <=  8'h74;        memory[31237] <=  8'h75;        memory[31238] <=  8'h79;        memory[31239] <=  8'h69;        memory[31240] <=  8'h75;        memory[31241] <=  8'h68;        memory[31242] <=  8'h6a;        memory[31243] <=  8'h6b;        memory[31244] <=  8'h62;        memory[31245] <=  8'h76;        memory[31246] <=  8'h63;        memory[31247] <=  8'h66;        memory[31248] <=  8'h74;        memory[31249] <=  8'h75;        memory[31250] <=  8'h79;        memory[31251] <=  8'h69;        memory[31252] <=  8'h75;        memory[31253] <=  8'h6a;        memory[31254] <=  8'h6b;        memory[31255] <=  8'h6e;        memory[31256] <=  8'h62;        memory[31257] <=  8'h76;        memory[31258] <=  8'h67;        memory[31259] <=  8'h66;        memory[31260] <=  8'h74;        memory[31261] <=  8'h79;        memory[31262] <=  8'h75;        memory[31263] <=  8'h75;        memory[31264] <=  8'h69;        memory[31265] <=  8'h6a;        memory[31266] <=  8'h6b;        memory[31267] <=  8'h68;        memory[31268] <=  8'h62;        memory[31269] <=  8'h6a;        memory[31270] <=  8'h67;        memory[31271] <=  8'h68;        memory[31272] <=  8'h66;        memory[31273] <=  8'h79;        memory[31274] <=  8'h74;        memory[31275] <=  8'h79;        memory[31276] <=  8'h69;        memory[31277] <=  8'h75;        memory[31278] <=  8'h64;        memory[31279] <=  8'h6a;        memory[31280] <=  8'h6b;        memory[31281] <=  8'h68;        memory[31282] <=  8'h63;        memory[31283] <=  8'h7a;        memory[31284] <=  8'h67;        memory[31285] <=  8'h68;        memory[31286] <=  8'h74;        memory[31287] <=  8'h75;        memory[31288] <=  8'h79;        memory[31289] <=  8'h69;        memory[31290] <=  8'h61;        memory[31291] <=  8'h73;        memory[31292] <=  8'h75;        memory[31293] <=  8'h6a;        memory[31294] <=  8'h6b;        memory[31295] <=  8'h62;        memory[31296] <=  8'h6e;        memory[31297] <=  8'h61;        memory[31298] <=  8'h76;        memory[31299] <=  8'h63;        memory[31300] <=  8'h66;        memory[31301] <=  8'h68;        memory[31302] <=  8'h75;        memory[31303] <=  8'h61;        memory[31304] <=  8'h73;        memory[31305] <=  8'h79;        memory[31306] <=  8'h64;        memory[31307] <=  8'h75;        memory[31308] <=  8'h69;        memory[31309] <=  8'h6a;        memory[31310] <=  8'h61;        memory[31311] <=  8'h6b;        memory[31312] <=  8'h62;        memory[31313] <=  8'h63;        memory[31314] <=  8'h78;        memory[31315] <=  8'h68;        memory[31316] <=  8'h67;        memory[31317] <=  8'h79;        memory[31318] <=  8'h75;        memory[31319] <=  8'h7a;        memory[31320] <=  8'h63;        memory[31321] <=  8'h61;        memory[31322] <=  8'h73;        memory[31323] <=  8'h69;        memory[31324] <=  8'h75;        memory[31325] <=  8'h6f;        memory[31326] <=  8'h69;        memory[31327] <=  8'h6a;        memory[31328] <=  8'h61;        memory[31329] <=  8'h6c;        memory[31330] <=  8'h63;        memory[31331] <=  8'h78;        memory[31332] <=  8'h62;        memory[31333] <=  8'h63;        memory[31334] <=  8'h20;        memory[31335] <=  8'h6e;        memory[31336] <=  8'h76;        memory[31337] <=  8'h63;        memory[31338] <=  8'h61;        memory[31339] <=  8'h64;        memory[31340] <=  8'h73;        memory[31341] <=  8'h67;        memory[31342] <=  8'h79;        memory[31343] <=  8'h68;        memory[31344] <=  8'h75;        memory[31345] <=  8'h61;        memory[31346] <=  8'h6a;        memory[31347] <=  8'h6b;        memory[31348] <=  8'h78;        memory[31349] <=  8'h62;        memory[31350] <=  8'h20;        memory[31351] <=  8'h6e;        memory[31352] <=  8'h76;        memory[31353] <=  8'h63;        memory[31354] <=  8'h61;        memory[31355] <=  8'h73;        memory[31356] <=  8'h67;        memory[31357] <=  8'h68;        memory[31358] <=  8'h75;        memory[31359] <=  8'h6a;        memory[31360] <=  8'h6c;        memory[31361] <=  8'h6b;        memory[31362] <=  8'h63;        memory[31363] <=  8'h78;        memory[31364] <=  8'h20;        memory[31365] <=  8'h6a;        memory[31366] <=  8'h6b;        memory[31367] <=  8'h68;        memory[31368] <=  8'h61;        memory[31369] <=  8'h73;        memory[31370] <=  8'h76;        memory[31371] <=  8'h64;        memory[31372] <=  8'h6e;        memory[31373] <=  8'h20;        memory[31374] <=  8'h62;        memory[31375] <=  8'h6e;        memory[31376] <=  8'h6d;        memory[31377] <=  8'h6b;        memory[31378] <=  8'h77;        memory[31379] <=  8'h64;        memory[31380] <=  8'h6f;        memory[31381] <=  8'h77;        memory[31382] <=  8'h69;        memory[31383] <=  8'h6f;        memory[31384] <=  8'h75;        memory[31385] <=  8'h69;        memory[31386] <=  8'h68;        memory[31387] <=  8'h62;        memory[31388] <=  8'h6e;        memory[31389] <=  8'h6b;        memory[31390] <=  8'h77;        memory[31391] <=  8'h69;        memory[31392] <=  8'h6f;        memory[31393] <=  8'h75;        memory[31394] <=  8'h71;        memory[31395] <=  8'h69;        memory[31396] <=  8'h79;        memory[31397] <=  8'h67;        memory[31398] <=  8'h6a;        memory[31399] <=  8'h64;        memory[31400] <=  8'h61;        memory[31401] <=  8'h76;        memory[31402] <=  8'h62;        memory[31403] <=  8'h6e;        memory[31404] <=  8'h6b;        memory[31405] <=  8'h6f;        memory[31406] <=  8'h70;        memory[31407] <=  8'h64;        memory[31408] <=  8'h76;        memory[31409] <=  8'h69;        memory[31410] <=  8'h6f;        memory[31411] <=  8'h75;        memory[31412] <=  8'h69;        memory[31413] <=  8'h48;        memory[31414] <=  8'h42;        memory[31415] <=  8'h6b;        memory[31416] <=  8'h64;        memory[31417] <=  8'h6e;        memory[31418] <=  8'h6c;        memory[31419] <=  8'h71;        memory[31420] <=  8'h6b;        memory[31421] <=  8'h6d;        memory[31422] <=  8'h6a;        memory[31423] <=  8'h70;        memory[31424] <=  8'h69;        memory[31425] <=  8'h6f;        memory[31426] <=  8'h68;        memory[31427] <=  8'h65;        memory[31428] <=  8'h66;        memory[31429] <=  8'h75;        memory[31430] <=  8'h67;        memory[31431] <=  8'h69;        memory[31432] <=  8'h73;        memory[31433] <=  8'h61;        memory[31434] <=  8'h62;        memory[31435] <=  8'h64;        memory[31436] <=  8'h6b;        memory[31437] <=  8'h6a;        memory[31438] <=  8'h6b;        memory[31439] <=  8'h6c;        memory[31440] <=  8'h6a;        memory[31441] <=  8'h69;        memory[31442] <=  8'h73;        memory[31443] <=  8'h6f;        memory[31444] <=  8'h71;        memory[31445] <=  8'h68;        memory[31446] <=  8'h77;        memory[31447] <=  8'h67;        memory[31448] <=  8'h69;        memory[31449] <=  8'h79;        memory[31450] <=  8'h6a;        memory[31451] <=  8'h64;        memory[31452] <=  8'h76;        memory[31453] <=  8'h62;        memory[31454] <=  8'h6e;        memory[31455] <=  8'h61;        memory[31456] <=  8'h73;        memory[31457] <=  8'h66;        memory[31458] <=  8'h6c;        memory[31459] <=  8'h6b;        memory[31460] <=  8'h64;        memory[31461] <=  8'h6a;        memory[31462] <=  8'h68;        memory[31463] <=  8'h63;        memory[31464] <=  8'h67;        memory[31465] <=  8'h6a;        memory[31466] <=  8'h76;        memory[31467] <=  8'h73;        memory[31468] <=  8'h64;        memory[31469] <=  8'h62;        memory[31470] <=  8'h62;        memory[31471] <=  8'h61;        memory[31472] <=  8'h72;        memory[31473] <=  8'h62;        memory[31474] <=  8'h62;        memory[31475] <=  8'h73;        memory[31476] <=  8'h62;        memory[31477] <=  8'h67;        memory[31478] <=  8'h73;        memory[31479] <=  8'h66;        memory[31480] <=  8'h67;        memory[31481] <=  8'h61;        memory[31482] <=  8'h68;        memory[31483] <=  8'h66;        memory[31484] <=  8'h73;        memory[31485] <=  8'h68;        memory[31486] <=  8'h61;        memory[31487] <=  8'h66;        memory[31488] <=  8'h73;        memory[31489] <=  8'h66;        memory[31490] <=  8'h68;        memory[31491] <=  8'h61;        memory[31492] <=  8'h69;        memory[31493] <=  8'h64;        memory[31494] <=  8'h75;        memory[31495] <=  8'h67;        memory[31496] <=  8'h64;        memory[31497] <=  8'h77;        memory[31498] <=  8'h62;        memory[31499] <=  8'h61;        memory[31500] <=  8'h62;        memory[31501] <=  8'h72;        memory[31502] <=  8'h62;        memory[31503] <=  8'h61;        memory[31504] <=  8'h62;        memory[31505] <=  8'h62;        memory[31506] <=  8'h74;        memory[31507] <=  8'h62;        memory[31508] <=  8'h62;        memory[31509] <=  8'h62;        memory[31510] <=  8'h62;        memory[31511] <=  8'h62;        memory[31512] <=  8'h62;        memory[31513] <=  8'h62;        memory[31514] <=  8'h62;        memory[31515] <=  8'h61;        memory[31516] <=  8'h62;        memory[31517] <=  8'h62;        memory[31518] <=  8'h72;        memory[31519] <=  8'h74;        memory[31520] <=  8'h62;        memory[31521] <=  8'h62;        memory[31522] <=  8'h61;        memory[31523] <=  8'h62;        memory[31524] <=  8'h72;        memory[31525] <=  8'h62;        memory[31526] <=  8'h74;        memory[31527] <=  8'h62;        memory[31528] <=  8'h62;        memory[31529] <=  8'h62;        memory[31530] <=  8'h63;        memory[31531] <=  8'h61;        memory[31532] <=  8'h72;        memory[31533] <=  8'h74;        memory[31534] <=  8'h73;        memory[31535] <=  8'h62;        memory[31536] <=  8'h61;        memory[31537] <=  8'h72;        memory[31538] <=  8'h74;        memory[31539] <=  8'h74;        memory[31540] <=  8'h62;        memory[31541] <=  8'h61;        memory[31542] <=  8'h72;        memory[31543] <=  8'h74;        memory[31544] <=  8'h78;        memory[31545] <=  8'h61;        memory[31546] <=  8'h74;        memory[31547] <=  8'h6b;        memory[31548] <=  8'h73;        memory[31549] <=  8'h68;        memory[31550] <=  8'h63;        memory[31551] <=  8'h66;        memory[31552] <=  8'h69;        memory[31553] <=  8'h77;        memory[31554] <=  8'h68;        memory[31555] <=  8'h61;        memory[31556] <=  8'h74;        memory[31557] <=  8'h61;        memory[31558] <=  8'h6e;        memory[31559] <=  8'h61;        memory[31560] <=  8'h62;        memory[31561] <=  8'h61;        memory[31562] <=  8'h63;        memory[31563] <=  8'h61;        memory[31564] <=  8'h74;        memory[31565] <=  8'h61;        memory[31566] <=  8'h62;        memory[31567] <=  8'h61;        memory[31568] <=  8'h72;        memory[31569] <=  8'h63;        memory[31570] <=  8'h61;        memory[31571] <=  8'h68;        memory[31572] <=  8'h64;        memory[31573] <=  8'h75;        memory[31574] <=  8'h63;        memory[31575] <=  8'h74;        memory[31576] <=  8'h61;        memory[31577] <=  8'h64;        memory[31578] <=  8'h61;        memory[31579] <=  8'h61;        memory[31580] <=  8'h63;        memory[31581] <=  8'h61;        memory[31582] <=  8'h72;        memory[31583] <=  8'h63;        memory[31584] <=  8'h74;        memory[31585] <=  8'h72;        memory[31586] <=  8'h63;        memory[31587] <=  8'h61;        memory[31588] <=  8'h74;        memory[31589] <=  8'h72;        memory[31590] <=  8'h63;        memory[31591] <=  8'h61;        memory[31592] <=  8'h74;        memory[31593] <=  8'h63;        memory[31594] <=  8'h62;        memory[31595] <=  8'h61;        memory[31596] <=  8'h74;        memory[31597] <=  8'h62;        memory[31598] <=  8'h72;        memory[31599] <=  8'h63;        memory[31600] <=  8'h61;        memory[31601] <=  8'h74;        memory[31602] <=  8'h72;        memory[31603] <=  8'h6e;        memory[31604] <=  8'h62;        memory[31605] <=  8'h61;        memory[31606] <=  8'h63;        memory[31607] <=  8'h61;        memory[31608] <=  8'h74;        memory[31609] <=  8'h79;        memory[31610] <=  8'h73;        memory[31611] <=  8'h6e;        memory[31612] <=  8'h63;        memory[31613] <=  8'h74;        memory[31614] <=  8'h61;        memory[31615] <=  8'h6e;        memory[31616] <=  8'h62;        memory[31617] <=  8'h61;        memory[31618] <=  8'h63;        memory[31619] <=  8'h72;        memory[31620] <=  8'h6e;        memory[31621] <=  8'h74;        memory[31622] <=  8'h61;        memory[31623] <=  8'h62;        memory[31624] <=  8'h74;        memory[31625] <=  8'h6e;        memory[31626] <=  8'h61;        memory[31627] <=  8'h72;        memory[31628] <=  8'h62;        memory[31629] <=  8'h78;        memory[31630] <=  8'h74;        memory[31631] <=  8'h61;        memory[31632] <=  8'h72;        memory[31633] <=  8'h62;        memory[31634] <=  8'h61;        memory[31635] <=  8'h72;        memory[31636] <=  8'h74;        memory[31637] <=  8'h74;        memory[31638] <=  8'h62;        memory[31639] <=  8'h61;        memory[31640] <=  8'h72;        memory[31641] <=  8'h74;        memory[31642] <=  8'h78;        memory[31643] <=  8'h61;        memory[31644] <=  8'h74;        memory[31645] <=  8'h6b;        memory[31646] <=  8'h73;        memory[31647] <=  8'h68;        memory[31648] <=  8'h63;        memory[31649] <=  8'h66;        memory[31650] <=  8'h69;        memory[31651] <=  8'h77;        memory[31652] <=  8'h68;        memory[31653] <=  8'h61;        memory[31654] <=  8'h74;        memory[31655] <=  8'h61;        memory[31656] <=  8'h6e;        memory[31657] <=  8'h61;        memory[31658] <=  8'h62;        memory[31659] <=  8'h61;        memory[31660] <=  8'h63;        memory[31661] <=  8'h61;        memory[31662] <=  8'h74;        memory[31663] <=  8'h61;        memory[31664] <=  8'h62;        memory[31665] <=  8'h61;        memory[31666] <=  8'h72;        memory[31667] <=  8'h63;        memory[31668] <=  8'h61;        memory[31669] <=  8'h68;        memory[31670] <=  8'h64;        memory[31671] <=  8'h75;        memory[31672] <=  8'h63;        memory[31673] <=  8'h74;        memory[31674] <=  8'h61;        memory[31675] <=  8'h64;        memory[31676] <=  8'h61;        memory[31677] <=  8'h61;        memory[31678] <=  8'h63;        memory[31679] <=  8'h61;        memory[31680] <=  8'h72;        memory[31681] <=  8'h63;        memory[31682] <=  8'h74;        memory[31683] <=  8'h72;        memory[31684] <=  8'h63;        memory[31685] <=  8'h61;        memory[31686] <=  8'h74;        memory[31687] <=  8'h72;        memory[31688] <=  8'h63;        memory[31689] <=  8'h61;        memory[31690] <=  8'h74;        memory[31691] <=  8'h63;        memory[31692] <=  8'h62;        memory[31693] <=  8'h61;        memory[31694] <=  8'h74;        memory[31695] <=  8'h62;        memory[31696] <=  8'h72;        memory[31697] <=  8'h63;        memory[31698] <=  8'h61;        memory[31699] <=  8'h74;        memory[31700] <=  8'h72;        memory[31701] <=  8'h6e;        memory[31702] <=  8'h62;        memory[31703] <=  8'h61;        memory[31704] <=  8'h63;        memory[31705] <=  8'h61;        memory[31706] <=  8'h74;        memory[31707] <=  8'h79;        memory[31708] <=  8'h73;        memory[31709] <=  8'h6e;        memory[31710] <=  8'h63;        memory[31711] <=  8'h74;        memory[31712] <=  8'h61;        memory[31713] <=  8'h6e;        memory[31714] <=  8'h62;        memory[31715] <=  8'h61;        memory[31716] <=  8'h63;        memory[31717] <=  8'h72;        memory[31718] <=  8'h6e;        memory[31719] <=  8'h74;        memory[31720] <=  8'h61;        memory[31721] <=  8'h62;        memory[31722] <=  8'h74;        memory[31723] <=  8'h6e;        memory[31724] <=  8'h61;        memory[31725] <=  8'h72;        memory[31726] <=  8'h62;        memory[31727] <=  8'h78;        memory[31728] <=  8'h74;        memory[31729] <=  8'h61;        memory[31730] <=  8'h72;        memory[31731] <=  8'h62;        memory[31732] <=  8'h61;        memory[31733] <=  8'h72;        memory[31734] <=  8'h74;        memory[31735] <=  8'h74;        memory[31736] <=  8'h62;        memory[31737] <=  8'h61;        memory[31738] <=  8'h72;        memory[31739] <=  8'h74;        memory[31740] <=  8'h78;        memory[31741] <=  8'h61;        memory[31742] <=  8'h74;        memory[31743] <=  8'h6b;        memory[31744] <=  8'h73;        memory[31745] <=  8'h68;        memory[31746] <=  8'h63;        memory[31747] <=  8'h66;        memory[31748] <=  8'h69;        memory[31749] <=  8'h77;        memory[31750] <=  8'h68;        memory[31751] <=  8'h61;        memory[31752] <=  8'h74;        memory[31753] <=  8'h61;        memory[31754] <=  8'h6e;        memory[31755] <=  8'h61;        memory[31756] <=  8'h62;        memory[31757] <=  8'h61;        memory[31758] <=  8'h63;        memory[31759] <=  8'h61;        memory[31760] <=  8'h74;        memory[31761] <=  8'h61;        memory[31762] <=  8'h62;        memory[31763] <=  8'h61;        memory[31764] <=  8'h72;        memory[31765] <=  8'h63;        memory[31766] <=  8'h61;        memory[31767] <=  8'h68;        memory[31768] <=  8'h64;        memory[31769] <=  8'h75;        memory[31770] <=  8'h63;        memory[31771] <=  8'h74;        memory[31772] <=  8'h61;        memory[31773] <=  8'h64;        memory[31774] <=  8'h61;        memory[31775] <=  8'h61;        memory[31776] <=  8'h63;        memory[31777] <=  8'h61;        memory[31778] <=  8'h72;        memory[31779] <=  8'h63;        memory[31780] <=  8'h74;        memory[31781] <=  8'h72;        memory[31782] <=  8'h63;        memory[31783] <=  8'h61;        memory[31784] <=  8'h74;        memory[31785] <=  8'h72;        memory[31786] <=  8'h63;        memory[31787] <=  8'h61;        memory[31788] <=  8'h74;        memory[31789] <=  8'h63;        memory[31790] <=  8'h62;        memory[31791] <=  8'h61;        memory[31792] <=  8'h74;        memory[31793] <=  8'h62;        memory[31794] <=  8'h72;        memory[31795] <=  8'h63;        memory[31796] <=  8'h61;        memory[31797] <=  8'h74;        memory[31798] <=  8'h72;        memory[31799] <=  8'h6e;        memory[31800] <=  8'h62;        memory[31801] <=  8'h61;        memory[31802] <=  8'h63;        memory[31803] <=  8'h61;        memory[31804] <=  8'h74;        memory[31805] <=  8'h79;        memory[31806] <=  8'h73;        memory[31807] <=  8'h6e;        memory[31808] <=  8'h63;        memory[31809] <=  8'h74;        memory[31810] <=  8'h61;        memory[31811] <=  8'h6e;        memory[31812] <=  8'h62;        memory[31813] <=  8'h61;        memory[31814] <=  8'h63;        memory[31815] <=  8'h72;        memory[31816] <=  8'h6e;        memory[31817] <=  8'h74;        memory[31818] <=  8'h61;        memory[31819] <=  8'h62;        memory[31820] <=  8'h74;        memory[31821] <=  8'h6e;        memory[31822] <=  8'h61;        memory[31823] <=  8'h72;        memory[31824] <=  8'h62;        memory[31825] <=  8'h78;        memory[31826] <=  8'h74;        memory[31827] <=  8'h61;        memory[31828] <=  8'h72;        memory[31829] <=  8'h5d;        memory[31830] <=  8'h5d;        memory[31831] <=  8'h65;        memory[31832] <=  8'h66;        memory[31833] <=  8'h77;        memory[31834] <=  8'h65;        memory[31835] <=  8'h5d;        memory[31836] <=  8'h65;        memory[31837] <=  8'h67;        memory[31838] <=  8'h73;        memory[31839] <=  8'h67;        memory[31840] <=  8'h66;        memory[31841] <=  8'h62;        memory[31842] <=  8'h61;        memory[31843] <=  8'h72;        memory[31844] <=  8'h74;        memory[31845] <=  8'h74;        memory[31846] <=  8'h62;        memory[31847] <=  8'h61;        memory[31848] <=  8'h72;        memory[31849] <=  8'h74;        memory[31850] <=  8'h78;        memory[31851] <=  8'h61;        memory[31852] <=  8'h74;        memory[31853] <=  8'h6b;        memory[31854] <=  8'h73;        memory[31855] <=  8'h68;        memory[31856] <=  8'h63;        memory[31857] <=  8'h66;        memory[31858] <=  8'h69;        memory[31859] <=  8'h77;        memory[31860] <=  8'h68;        memory[31861] <=  8'h61;        memory[31862] <=  8'h74;        memory[31863] <=  8'h61;        memory[31864] <=  8'h6e;        memory[31865] <=  8'h61;        memory[31866] <=  8'h62;        memory[31867] <=  8'h61;        memory[31868] <=  8'h63;        memory[31869] <=  8'h61;        memory[31870] <=  8'h74;        memory[31871] <=  8'h61;        memory[31872] <=  8'h62;        memory[31873] <=  8'h61;        memory[31874] <=  8'h72;        memory[31875] <=  8'h63;        memory[31876] <=  8'h61;        memory[31877] <=  8'h68;        memory[31878] <=  8'h64;        memory[31879] <=  8'h75;        memory[31880] <=  8'h63;        memory[31881] <=  8'h74;        memory[31882] <=  8'h61;        memory[31883] <=  8'h64;        memory[31884] <=  8'h61;        memory[31885] <=  8'h61;        memory[31886] <=  8'h63;        memory[31887] <=  8'h61;        memory[31888] <=  8'h72;        memory[31889] <=  8'h63;        memory[31890] <=  8'h74;        memory[31891] <=  8'h72;        memory[31892] <=  8'h63;        memory[31893] <=  8'h61;        memory[31894] <=  8'h74;        memory[31895] <=  8'h72;        memory[31896] <=  8'h63;        memory[31897] <=  8'h61;        memory[31898] <=  8'h74;        memory[31899] <=  8'h63;        memory[31900] <=  8'h62;        memory[31901] <=  8'h61;        memory[31902] <=  8'h74;        memory[31903] <=  8'h62;        memory[31904] <=  8'h72;        memory[31905] <=  8'h63;        memory[31906] <=  8'h61;        memory[31907] <=  8'h74;        memory[31908] <=  8'h72;        memory[31909] <=  8'h6e;        memory[31910] <=  8'h62;        memory[31911] <=  8'h61;        memory[31912] <=  8'h63;        memory[31913] <=  8'h61;        memory[31914] <=  8'h74;        memory[31915] <=  8'h79;        memory[31916] <=  8'h73;        memory[31917] <=  8'h6e;        memory[31918] <=  8'h63;        memory[31919] <=  8'h74;        memory[31920] <=  8'h61;        memory[31921] <=  8'h6e;        memory[31922] <=  8'h62;        memory[31923] <=  8'h61;        memory[31924] <=  8'h63;        memory[31925] <=  8'h72;        memory[31926] <=  8'h6e;        memory[31927] <=  8'h74;        memory[31928] <=  8'h61;        memory[31929] <=  8'h62;        memory[31930] <=  8'h74;        memory[31931] <=  8'h6e;        memory[31932] <=  8'h61;        memory[31933] <=  8'h72;        memory[31934] <=  8'h62;        memory[31935] <=  8'h78;        memory[31936] <=  8'h74;        memory[31937] <=  8'h61;        memory[31938] <=  8'h72;        memory[31939] <=  8'h62;        memory[31940] <=  8'h61;        memory[31941] <=  8'h72;        memory[31942] <=  8'h74;        memory[31943] <=  8'h74;        memory[31944] <=  8'h62;        memory[31945] <=  8'h61;        memory[31946] <=  8'h72;        memory[31947] <=  8'h74;        memory[31948] <=  8'h78;        memory[31949] <=  8'h61;        memory[31950] <=  8'h74;        memory[31951] <=  8'h6b;        memory[31952] <=  8'h73;        memory[31953] <=  8'h68;        memory[31954] <=  8'h63;        memory[31955] <=  8'h66;        memory[31956] <=  8'h69;        memory[31957] <=  8'h77;        memory[31958] <=  8'h68;        memory[31959] <=  8'h61;        memory[31960] <=  8'h74;        memory[31961] <=  8'h61;        memory[31962] <=  8'h6e;        memory[31963] <=  8'h61;        memory[31964] <=  8'h62;        memory[31965] <=  8'h61;        memory[31966] <=  8'h63;        memory[31967] <=  8'h61;        memory[31968] <=  8'h74;        memory[31969] <=  8'h61;        memory[31970] <=  8'h62;        memory[31971] <=  8'h61;        memory[31972] <=  8'h72;        memory[31973] <=  8'h63;        memory[31974] <=  8'h61;        memory[31975] <=  8'h68;        memory[31976] <=  8'h64;        memory[31977] <=  8'h75;        memory[31978] <=  8'h63;        memory[31979] <=  8'h74;        memory[31980] <=  8'h61;        memory[31981] <=  8'h64;        memory[31982] <=  8'h61;        memory[31983] <=  8'h61;        memory[31984] <=  8'h63;        memory[31985] <=  8'h61;        memory[31986] <=  8'h72;        memory[31987] <=  8'h63;        memory[31988] <=  8'h74;        memory[31989] <=  8'h72;        memory[31990] <=  8'h63;        memory[31991] <=  8'h61;        memory[31992] <=  8'h74;        memory[31993] <=  8'h72;        memory[31994] <=  8'h63;        memory[31995] <=  8'h61;        memory[31996] <=  8'h74;        memory[31997] <=  8'h63;        memory[31998] <=  8'h62;        memory[31999] <=  8'h61;        memory[32000] <=  8'h74;        memory[32001] <=  8'h62;        memory[32002] <=  8'h72;        memory[32003] <=  8'h63;        memory[32004] <=  8'h61;        memory[32005] <=  8'h74;        memory[32006] <=  8'h72;        memory[32007] <=  8'h6e;        memory[32008] <=  8'h62;        memory[32009] <=  8'h61;        memory[32010] <=  8'h63;        memory[32011] <=  8'h61;        memory[32012] <=  8'h74;        memory[32013] <=  8'h79;        memory[32014] <=  8'h73;        memory[32015] <=  8'h6e;        memory[32016] <=  8'h63;        memory[32017] <=  8'h74;        memory[32018] <=  8'h61;        memory[32019] <=  8'h6e;        memory[32020] <=  8'h62;        memory[32021] <=  8'h61;        memory[32022] <=  8'h63;        memory[32023] <=  8'h72;        memory[32024] <=  8'h6e;        memory[32025] <=  8'h74;        memory[32026] <=  8'h61;        memory[32027] <=  8'h62;        memory[32028] <=  8'h74;        memory[32029] <=  8'h6e;        memory[32030] <=  8'h61;        memory[32031] <=  8'h72;        memory[32032] <=  8'h62;        memory[32033] <=  8'h78;        memory[32034] <=  8'h74;        memory[32035] <=  8'h61;        memory[32036] <=  8'h72;        memory[32037] <=  8'h64;        memory[32038] <=  8'h66;        memory[32039] <=  8'h73;        memory[32040] <=  8'h67;        memory[32041] <=  8'h76;        memory[32042] <=  8'h68;        memory[32043] <=  8'h62;        memory[32044] <=  8'h6b;        memory[32045] <=  8'h6a;        memory[32046] <=  8'h6e;        memory[32047] <=  8'h6d;        memory[32048] <=  8'h62;        memory[32049] <=  8'h76;        memory[32050] <=  8'h78;        memory[32051] <=  8'h63;        memory[32052] <=  8'h73;        memory[32053] <=  8'h66;        memory[32054] <=  8'h72;        memory[32055] <=  8'h74;        memory[32056] <=  8'h79;        memory[32057] <=  8'h75;        memory[32058] <=  8'h6a;        memory[32059] <=  8'h6e;        memory[32060] <=  8'h62;        memory[32061] <=  8'h76;        memory[32062] <=  8'h63;        memory[32063] <=  8'h64;        memory[32064] <=  8'h74;        memory[32065] <=  8'h79;        memory[32066] <=  8'h75;        memory[32067] <=  8'h69;        memory[32068] <=  8'h6b;        memory[32069] <=  8'h6d;        memory[32070] <=  8'h6e;        memory[32071] <=  8'h62;        memory[32072] <=  8'h76;        memory[32073] <=  8'h63;        memory[32074] <=  8'h78;        memory[32075] <=  8'h73;        memory[32076] <=  8'h64;        memory[32077] <=  8'h72;        memory[32078] <=  8'h74;        memory[32079] <=  8'h79;        memory[32080] <=  8'h75;        memory[32081] <=  8'h69;        memory[32082] <=  8'h6b;        memory[32083] <=  8'h6d;        memory[32084] <=  8'h6e;        memory[32085] <=  8'h62;        memory[32086] <=  8'h76;        memory[32087] <=  8'h63;        memory[32088] <=  8'h73;        memory[32089] <=  8'h77;        memory[32090] <=  8'h33;        memory[32091] <=  8'h34;        memory[32092] <=  8'h35;        memory[32093] <=  8'h36;        memory[32094] <=  8'h37;        memory[32095] <=  8'h38;        memory[32096] <=  8'h69;        memory[32097] <=  8'h6b;        memory[32098] <=  8'h6d;        memory[32099] <=  8'h6e;        memory[32100] <=  8'h62;        memory[32101] <=  8'h76;        memory[32102] <=  8'h63;        memory[32103] <=  8'h64;        memory[32104] <=  8'h65;        memory[32105] <=  8'h72;        memory[32106] <=  8'h36;        memory[32107] <=  8'h37;        memory[32108] <=  8'h38;        memory[32109] <=  8'h69;        memory[32110] <=  8'h6f;        memory[32111] <=  8'h6b;        memory[32112] <=  8'h6a;        memory[32113] <=  8'h6e;        memory[32114] <=  8'h62;        memory[32115] <=  8'h76;        memory[32116] <=  8'h63;        memory[32117] <=  8'h64;        memory[32118] <=  8'h72;        memory[32119] <=  8'h74;        memory[32120] <=  8'h79;        memory[32121] <=  8'h75;        memory[32122] <=  8'h73;        memory[32123] <=  8'h6a;        memory[32124] <=  8'h63;        memory[32125] <=  8'h6e;        memory[32126] <=  8'h62;        memory[32127] <=  8'h64;        memory[32128] <=  8'h66;        memory[32129] <=  8'h73;        memory[32130] <=  8'h74;        memory[32131] <=  8'h79;        memory[32132] <=  8'h75;        memory[32133] <=  8'h61;        memory[32134] <=  8'h69;        memory[32135] <=  8'h6b;        memory[32136] <=  8'h78;        memory[32137] <=  8'h6d;        memory[32138] <=  8'h6e;        memory[32139] <=  8'h73;        memory[32140] <=  8'h6a;        memory[32141] <=  8'h6f;        memory[32142] <=  8'h64;        memory[32143] <=  8'h6c;        memory[32144] <=  8'h63;        memory[32145] <=  8'h78;        memory[32146] <=  8'h62;        memory[32147] <=  8'h61;        memory[32148] <=  8'h72;        memory[32149] <=  8'h74;        memory[32150] <=  8'h78;        memory[32151] <=  8'h61;        memory[32152] <=  8'h74;        memory[32153] <=  8'h6b;        memory[32154] <=  8'h73;        memory[32155] <=  8'h68;        memory[32156] <=  8'h63;        memory[32157] <=  8'h66;        memory[32158] <=  8'h69;        memory[32159] <=  8'h77;        memory[32160] <=  8'h68;        memory[32161] <=  8'h61;        memory[32162] <=  8'h74;        memory[32163] <=  8'h61;        memory[32164] <=  8'h6e;        memory[32165] <=  8'h61;        memory[32166] <=  8'h62;        memory[32167] <=  8'h61;        memory[32168] <=  8'h63;        memory[32169] <=  8'h61;        memory[32170] <=  8'h74;        memory[32171] <=  8'h61;        memory[32172] <=  8'h62;        memory[32173] <=  8'h61;        memory[32174] <=  8'h72;        memory[32175] <=  8'h63;        memory[32176] <=  8'h61;        memory[32177] <=  8'h68;        memory[32178] <=  8'h64;        memory[32179] <=  8'h75;        memory[32180] <=  8'h63;        memory[32181] <=  8'h74;        memory[32182] <=  8'h61;        memory[32183] <=  8'h64;        memory[32184] <=  8'h61;        memory[32185] <=  8'h61;        memory[32186] <=  8'h63;        memory[32187] <=  8'h61;        memory[32188] <=  8'h72;        memory[32189] <=  8'h62;        memory[32190] <=  8'h61;        memory[32191] <=  8'h72;        memory[32192] <=  8'h74;        memory[32193] <=  8'h78;        memory[32194] <=  8'h61;        memory[32195] <=  8'h74;        memory[32196] <=  8'h6b;        memory[32197] <=  8'h73;        memory[32198] <=  8'h68;        memory[32199] <=  8'h63;        memory[32200] <=  8'h66;        memory[32201] <=  8'h69;        memory[32202] <=  8'h77;        memory[32203] <=  8'h68;        memory[32204] <=  8'h61;        memory[32205] <=  8'h74;        memory[32206] <=  8'h61;        memory[32207] <=  8'h6e;        memory[32208] <=  8'h61;        memory[32209] <=  8'h62;        memory[32210] <=  8'h61;        memory[32211] <=  8'h63;        memory[32212] <=  8'h61;        memory[32213] <=  8'h74;        memory[32214] <=  8'h61;        memory[32215] <=  8'h62;        memory[32216] <=  8'h61;        memory[32217] <=  8'h72;        memory[32218] <=  8'h63;        memory[32219] <=  8'h61;        memory[32220] <=  8'h68;        memory[32221] <=  8'h64;        memory[32222] <=  8'h75;        memory[32223] <=  8'h63;        memory[32224] <=  8'h74;        memory[32225] <=  8'h61;        memory[32226] <=  8'h64;        memory[32227] <=  8'h61;        memory[32228] <=  8'h61;        memory[32229] <=  8'h63;        memory[32230] <=  8'h61;        memory[32231] <=  8'h72;        memory[32232] <=  8'h62;        memory[32233] <=  8'h61;        memory[32234] <=  8'h72;        memory[32235] <=  8'h74;        memory[32236] <=  8'h78;        memory[32237] <=  8'h61;        memory[32238] <=  8'h74;        memory[32239] <=  8'h6b;        memory[32240] <=  8'h73;        memory[32241] <=  8'h68;        memory[32242] <=  8'h63;        memory[32243] <=  8'h66;        memory[32244] <=  8'h69;        memory[32245] <=  8'h77;        memory[32246] <=  8'h68;        memory[32247] <=  8'h61;        memory[32248] <=  8'h74;        memory[32249] <=  8'h61;        memory[32250] <=  8'h6e;        memory[32251] <=  8'h61;        memory[32252] <=  8'h62;        memory[32253] <=  8'h61;        memory[32254] <=  8'h63;        memory[32255] <=  8'h61;        memory[32256] <=  8'h74;        memory[32257] <=  8'h61;        memory[32258] <=  8'h62;        memory[32259] <=  8'h61;        memory[32260] <=  8'h72;        memory[32261] <=  8'h63;        memory[32262] <=  8'h61;        memory[32263] <=  8'h68;        memory[32264] <=  8'h64;        memory[32265] <=  8'h75;        memory[32266] <=  8'h63;        memory[32267] <=  8'h74;        memory[32268] <=  8'h61;        memory[32269] <=  8'h64;        memory[32270] <=  8'h61;        memory[32271] <=  8'h61;        memory[32272] <=  8'h63;        memory[32273] <=  8'h61;        memory[32274] <=  8'h72;        memory[32275] <=  8'h62;        memory[32276] <=  8'h61;        memory[32277] <=  8'h72;        memory[32278] <=  8'h74;        memory[32279] <=  8'h78;        memory[32280] <=  8'h61;        memory[32281] <=  8'h74;        memory[32282] <=  8'h6b;        memory[32283] <=  8'h73;        memory[32284] <=  8'h68;        memory[32285] <=  8'h63;        memory[32286] <=  8'h66;        memory[32287] <=  8'h69;        memory[32288] <=  8'h77;        memory[32289] <=  8'h68;        memory[32290] <=  8'h61;        memory[32291] <=  8'h74;        memory[32292] <=  8'h61;        memory[32293] <=  8'h6e;        memory[32294] <=  8'h61;        memory[32295] <=  8'h62;        memory[32296] <=  8'h61;        memory[32297] <=  8'h63;        memory[32298] <=  8'h61;        memory[32299] <=  8'h74;        memory[32300] <=  8'h61;        memory[32301] <=  8'h62;        memory[32302] <=  8'h61;        memory[32303] <=  8'h72;        memory[32304] <=  8'h63;        memory[32305] <=  8'h61;        memory[32306] <=  8'h68;        memory[32307] <=  8'h64;        memory[32308] <=  8'h75;        memory[32309] <=  8'h63;        memory[32310] <=  8'h74;        memory[32311] <=  8'h61;        memory[32312] <=  8'h64;        memory[32313] <=  8'h61;        memory[32314] <=  8'h61;        memory[32315] <=  8'h63;        memory[32316] <=  8'h61;        memory[32317] <=  8'h72;        memory[32318] <=  8'h62;        memory[32319] <=  8'h61;        memory[32320] <=  8'h72;        memory[32321] <=  8'h74;        memory[32322] <=  8'h78;        memory[32323] <=  8'h61;        memory[32324] <=  8'h74;        memory[32325] <=  8'h6b;        memory[32326] <=  8'h73;        memory[32327] <=  8'h68;        memory[32328] <=  8'h63;        memory[32329] <=  8'h66;        memory[32330] <=  8'h69;        memory[32331] <=  8'h77;        memory[32332] <=  8'h68;        memory[32333] <=  8'h61;        memory[32334] <=  8'h74;        memory[32335] <=  8'h61;        memory[32336] <=  8'h6e;        memory[32337] <=  8'h61;        memory[32338] <=  8'h62;        memory[32339] <=  8'h61;        memory[32340] <=  8'h63;        memory[32341] <=  8'h61;        memory[32342] <=  8'h74;        memory[32343] <=  8'h61;        memory[32344] <=  8'h62;        memory[32345] <=  8'h61;        memory[32346] <=  8'h72;        memory[32347] <=  8'h63;        memory[32348] <=  8'h61;        memory[32349] <=  8'h68;        memory[32350] <=  8'h64;        memory[32351] <=  8'h75;        memory[32352] <=  8'h63;        memory[32353] <=  8'h74;        memory[32354] <=  8'h61;        memory[32355] <=  8'h64;        memory[32356] <=  8'h61;        memory[32357] <=  8'h61;        memory[32358] <=  8'h63;        memory[32359] <=  8'h61;        memory[32360] <=  8'h72;        memory[32361] <=  8'h62;        memory[32362] <=  8'h61;        memory[32363] <=  8'h72;        memory[32364] <=  8'h74;        memory[32365] <=  8'h78;        memory[32366] <=  8'h61;        memory[32367] <=  8'h74;        memory[32368] <=  8'h6b;        memory[32369] <=  8'h73;        memory[32370] <=  8'h68;        memory[32371] <=  8'h63;        memory[32372] <=  8'h66;        memory[32373] <=  8'h69;        memory[32374] <=  8'h77;        memory[32375] <=  8'h68;        memory[32376] <=  8'h61;        memory[32377] <=  8'h74;        memory[32378] <=  8'h61;        memory[32379] <=  8'h6e;        memory[32380] <=  8'h61;        memory[32381] <=  8'h62;        memory[32382] <=  8'h61;        memory[32383] <=  8'h63;        memory[32384] <=  8'h61;        memory[32385] <=  8'h74;        memory[32386] <=  8'h61;        memory[32387] <=  8'h62;        memory[32388] <=  8'h61;        memory[32389] <=  8'h72;        memory[32390] <=  8'h63;        memory[32391] <=  8'h61;        memory[32392] <=  8'h68;        memory[32393] <=  8'h64;        memory[32394] <=  8'h75;        memory[32395] <=  8'h63;        memory[32396] <=  8'h74;        memory[32397] <=  8'h61;        memory[32398] <=  8'h64;        memory[32399] <=  8'h61;        memory[32400] <=  8'h61;        memory[32401] <=  8'h63;        memory[32402] <=  8'h61;        memory[32403] <=  8'h72;        memory[32404] <=  8'h62;        memory[32405] <=  8'h61;        memory[32406] <=  8'h72;        memory[32407] <=  8'h74;        memory[32408] <=  8'h78;        memory[32409] <=  8'h61;        memory[32410] <=  8'h74;        memory[32411] <=  8'h6b;        memory[32412] <=  8'h73;        memory[32413] <=  8'h68;        memory[32414] <=  8'h63;        memory[32415] <=  8'h66;        memory[32416] <=  8'h69;        memory[32417] <=  8'h77;        memory[32418] <=  8'h68;        memory[32419] <=  8'h61;        memory[32420] <=  8'h74;        memory[32421] <=  8'h61;        memory[32422] <=  8'h6e;        memory[32423] <=  8'h61;        memory[32424] <=  8'h62;        memory[32425] <=  8'h61;        memory[32426] <=  8'h63;        memory[32427] <=  8'h61;        memory[32428] <=  8'h74;        memory[32429] <=  8'h61;        memory[32430] <=  8'h62;        memory[32431] <=  8'h61;        memory[32432] <=  8'h72;        memory[32433] <=  8'h63;        memory[32434] <=  8'h61;        memory[32435] <=  8'h68;        memory[32436] <=  8'h64;        memory[32437] <=  8'h75;        memory[32438] <=  8'h63;        memory[32439] <=  8'h74;        memory[32440] <=  8'h61;        memory[32441] <=  8'h64;        memory[32442] <=  8'h61;        memory[32443] <=  8'h61;        memory[32444] <=  8'h63;        memory[32445] <=  8'h61;        memory[32446] <=  8'h72;        memory[32447] <=  8'h62;        memory[32448] <=  8'h61;        memory[32449] <=  8'h72;        memory[32450] <=  8'h74;        memory[32451] <=  8'h78;        memory[32452] <=  8'h61;        memory[32453] <=  8'h74;        memory[32454] <=  8'h6b;        memory[32455] <=  8'h73;        memory[32456] <=  8'h68;        memory[32457] <=  8'h63;        memory[32458] <=  8'h66;        memory[32459] <=  8'h69;        memory[32460] <=  8'h77;        memory[32461] <=  8'h68;        memory[32462] <=  8'h61;        memory[32463] <=  8'h74;        memory[32464] <=  8'h61;        memory[32465] <=  8'h6e;        memory[32466] <=  8'h61;        memory[32467] <=  8'h62;        memory[32468] <=  8'h61;        memory[32469] <=  8'h63;        memory[32470] <=  8'h61;        memory[32471] <=  8'h74;        memory[32472] <=  8'h61;        memory[32473] <=  8'h62;        memory[32474] <=  8'h61;        memory[32475] <=  8'h72;        memory[32476] <=  8'h63;        memory[32477] <=  8'h61;        memory[32478] <=  8'h68;        memory[32479] <=  8'h64;        memory[32480] <=  8'h75;        memory[32481] <=  8'h63;        memory[32482] <=  8'h74;        memory[32483] <=  8'h61;        memory[32484] <=  8'h64;        memory[32485] <=  8'h61;        memory[32486] <=  8'h61;        memory[32487] <=  8'h63;        memory[32488] <=  8'h61;        memory[32489] <=  8'h72;        memory[32490] <=  8'h62;        memory[32491] <=  8'h61;        memory[32492] <=  8'h72;        memory[32493] <=  8'h74;        memory[32494] <=  8'h78;        memory[32495] <=  8'h61;        memory[32496] <=  8'h74;        memory[32497] <=  8'h6b;        memory[32498] <=  8'h73;        memory[32499] <=  8'h68;        memory[32500] <=  8'h63;        memory[32501] <=  8'h66;        memory[32502] <=  8'h69;        memory[32503] <=  8'h77;        memory[32504] <=  8'h68;        memory[32505] <=  8'h61;        memory[32506] <=  8'h74;        memory[32507] <=  8'h61;        memory[32508] <=  8'h6e;        memory[32509] <=  8'h61;        memory[32510] <=  8'h62;        memory[32511] <=  8'h61;        memory[32512] <=  8'h63;        memory[32513] <=  8'h61;        memory[32514] <=  8'h74;        memory[32515] <=  8'h61;        memory[32516] <=  8'h62;        memory[32517] <=  8'h61;        memory[32518] <=  8'h72;        memory[32519] <=  8'h63;        memory[32520] <=  8'h61;        memory[32521] <=  8'h68;        memory[32522] <=  8'h64;        memory[32523] <=  8'h75;        memory[32524] <=  8'h63;        memory[32525] <=  8'h74;        memory[32526] <=  8'h61;        memory[32527] <=  8'h64;        memory[32528] <=  8'h61;        memory[32529] <=  8'h61;        memory[32530] <=  8'h63;        memory[32531] <=  8'h61;        memory[32532] <=  8'h72;        memory[32533] <=  8'h62;        memory[32534] <=  8'h61;        memory[32535] <=  8'h72;        memory[32536] <=  8'h74;        memory[32537] <=  8'h74;        memory[32538] <=  8'h62;        memory[32539] <=  8'h61;        memory[32540] <=  8'h72;        memory[32541] <=  8'h74;        memory[32542] <=  8'h78;        memory[32543] <=  8'h61;        memory[32544] <=  8'h74;        memory[32545] <=  8'h6b;        memory[32546] <=  8'h73;        memory[32547] <=  8'h68;        memory[32548] <=  8'h63;        memory[32549] <=  8'h66;        memory[32550] <=  8'h69;        memory[32551] <=  8'h77;        memory[32552] <=  8'h68;        memory[32553] <=  8'h61;        memory[32554] <=  8'h74;        memory[32555] <=  8'h61;        memory[32556] <=  8'h6e;        memory[32557] <=  8'h61;        memory[32558] <=  8'h62;        memory[32559] <=  8'h61;        memory[32560] <=  8'h63;        memory[32561] <=  8'h61;        memory[32562] <=  8'h74;        memory[32563] <=  8'h61;        memory[32564] <=  8'h62;        memory[32565] <=  8'h61;        memory[32566] <=  8'h72;        memory[32567] <=  8'h63;        memory[32568] <=  8'h61;        memory[32569] <=  8'h68;        memory[32570] <=  8'h64;        memory[32571] <=  8'h75;        memory[32572] <=  8'h63;        memory[32573] <=  8'h74;        memory[32574] <=  8'h61;        memory[32575] <=  8'h64;        memory[32576] <=  8'h61;        memory[32577] <=  8'h61;        memory[32578] <=  8'h63;        memory[32579] <=  8'h61;        memory[32580] <=  8'h72;        memory[32581] <=  8'h63;        memory[32582] <=  8'h74;        memory[32583] <=  8'h72;        memory[32584] <=  8'h63;        memory[32585] <=  8'h61;        memory[32586] <=  8'h74;        memory[32587] <=  8'h72;        memory[32588] <=  8'h63;        memory[32589] <=  8'h61;        memory[32590] <=  8'h74;        memory[32591] <=  8'h63;        memory[32592] <=  8'h62;        memory[32593] <=  8'h61;        memory[32594] <=  8'h74;        memory[32595] <=  8'h62;        memory[32596] <=  8'h72;        memory[32597] <=  8'h63;        memory[32598] <=  8'h61;        memory[32599] <=  8'h72;        memory[32600] <=  8'h62;        memory[32601] <=  8'h78;        memory[32602] <=  8'h74;        memory[32603] <=  8'h61;        memory[32604] <=  8'h72;        memory[32605] <=  8'h64;        memory[32606] <=  8'h66;        memory[32607] <=  8'h73;        memory[32608] <=  8'h67;        memory[32609] <=  8'h76;        memory[32610] <=  8'h68;        memory[32611] <=  8'h62;        memory[32612] <=  8'h6b;        memory[32613] <=  8'h6a;        memory[32614] <=  8'h6e;        memory[32615] <=  8'h6d;        memory[32616] <=  8'h62;        memory[32617] <=  8'h76;        memory[32618] <=  8'h78;        memory[32619] <=  8'h63;        memory[32620] <=  8'h73;        memory[32621] <=  8'h66;        memory[32622] <=  8'h72;        memory[32623] <=  8'h74;        memory[32624] <=  8'h79;        memory[32625] <=  8'h75;        memory[32626] <=  8'h6a;        memory[32627] <=  8'h6e;        memory[32628] <=  8'h62;        memory[32629] <=  8'h76;        memory[32630] <=  8'h63;        memory[32631] <=  8'h64;        memory[32632] <=  8'h74;        memory[32633] <=  8'h79;        memory[32634] <=  8'h75;        memory[32635] <=  8'h69;        memory[32636] <=  8'h6b;        memory[32637] <=  8'h6d;        memory[32638] <=  8'h6e;        memory[32639] <=  8'h62;        memory[32640] <=  8'h76;        memory[32641] <=  8'h63;        memory[32642] <=  8'h78;        memory[32643] <=  8'h73;        memory[32644] <=  8'h64;        memory[32645] <=  8'h72;        memory[32646] <=  8'h74;        memory[32647] <=  8'h79;        memory[32648] <=  8'h75;        memory[32649] <=  8'h69;        memory[32650] <=  8'h6b;        memory[32651] <=  8'h6d;        memory[32652] <=  8'h6e;        memory[32653] <=  8'h62;        memory[32654] <=  8'h76;        memory[32655] <=  8'h63;        memory[32656] <=  8'h73;        memory[32657] <=  8'h77;        memory[32658] <=  8'h33;        memory[32659] <=  8'h34;        memory[32660] <=  8'h35;        memory[32661] <=  8'h36;        memory[32662] <=  8'h37;        memory[32663] <=  8'h38;        memory[32664] <=  8'h69;        memory[32665] <=  8'h6b;        memory[32666] <=  8'h6d;        memory[32667] <=  8'h6e;        memory[32668] <=  8'h62;        memory[32669] <=  8'h76;        memory[32670] <=  8'h63;        memory[32671] <=  8'h64;        memory[32672] <=  8'h65;        memory[32673] <=  8'h72;        memory[32674] <=  8'h36;        memory[32675] <=  8'h37;        memory[32676] <=  8'h38;        memory[32677] <=  8'h69;        memory[32678] <=  8'h6f;        memory[32679] <=  8'h6b;        memory[32680] <=  8'h6a;        memory[32681] <=  8'h6e;        memory[32682] <=  8'h62;        memory[32683] <=  8'h76;        memory[32684] <=  8'h63;        memory[32685] <=  8'h64;        memory[32686] <=  8'h72;        memory[32687] <=  8'h74;        memory[32688] <=  8'h79;        memory[32689] <=  8'h75;        memory[32690] <=  8'h73;        memory[32691] <=  8'h6a;        memory[32692] <=  8'h63;        memory[32693] <=  8'h6e;        memory[32694] <=  8'h62;        memory[32695] <=  8'h64;        memory[32696] <=  8'h66;        memory[32697] <=  8'h73;        memory[32698] <=  8'h74;        memory[32699] <=  8'h79;        memory[32700] <=  8'h75;        memory[32701] <=  8'h61;        memory[32702] <=  8'h69;        memory[32703] <=  8'h6b;        memory[32704] <=  8'h78;        memory[32705] <=  8'h6d;        memory[32706] <=  8'h6e;        memory[32707] <=  8'h73;        memory[32708] <=  8'h6a;        memory[32709] <=  8'h6f;        memory[32710] <=  8'h64;        memory[32711] <=  8'h6c;        memory[32712] <=  8'h63;        memory[32713] <=  8'h78;        memory[32714] <=  8'h2c;        memory[32715] <=  8'h6d;        memory[32716] <=  8'h73;        memory[32717] <=  8'h6b;        memory[32718] <=  8'h64;        memory[32719] <=  8'h6c;        memory[32720] <=  8'h70;        memory[32721] <=  8'h5b;        memory[32722] <=  8'h3b;        memory[32723] <=  8'h73;        memory[32724] <=  8'h6c;        memory[32725] <=  8'h64;        memory[32726] <=  8'h70;        memory[32727] <=  8'h76;        memory[32728] <=  8'h63;        memory[32729] <=  8'h5b;        memory[32730] <=  8'h78;        memory[32731] <=  8'h76;        memory[32732] <=  8'h63;        memory[32733] <=  8'h5b;        memory[32734] <=  8'h78;        memory[32735] <=  8'h70;        memory[32736] <=  8'h6f;        memory[32737] <=  8'h20;        memory[32738] <=  8'h62;        memory[32739] <=  8'h61;        memory[32740] <=  8'h72;        memory[32741] <=  8'h74;        memory[32742] <=  8'h74;        memory[32743] <=  8'h62;        memory[32744] <=  8'h61;        memory[32745] <=  8'h72;        memory[32746] <=  8'h74;        memory[32747] <=  8'h78;        memory[32748] <=  8'h61;        memory[32749] <=  8'h74;        memory[32750] <=  8'h6b;        memory[32751] <=  8'h73;        memory[32752] <=  8'h68;        memory[32753] <=  8'h63;        memory[32754] <=  8'h66;        memory[32755] <=  8'h69;        memory[32756] <=  8'h77;        memory[32757] <=  8'h68;        memory[32758] <=  8'h61;        memory[32759] <=  8'h69;        memory[32760] <=  8'h6a;        memory[32761] <=  8'h78;        memory[32762] <=  8'h5d;        memory[32763] <=  8'h65;        memory[32764] <=  8'h6b;        memory[32765] <=  8'h6f;        memory[32766] <=  8'h39;        memory[32767] <=  8'h64;        memory[32768] <=  8'h75;        memory[32769] <=  8'h38;        memory[32770] <=  8'h79;        memory[32771] <=  8'h20;        memory[32772] <=  8'h37;        memory[32773] <=  8'h63;        memory[32774] <=  8'h67;        memory[32775] <=  8'h78;        memory[32776] <=  8'h63;        memory[32777] <=  8'h75;        memory[32778] <=  8'h68;        memory[32779] <=  8'h69;        memory[32780] <=  8'h6a;        memory[32781] <=  8'h77;        memory[32782] <=  8'h69;        memory[32783] <=  8'h64;        memory[32784] <=  8'h66;        memory[32785] <=  8'h68;        memory[32786] <=  8'h75;        memory[32787] <=  8'h76;        memory[32788] <=  8'h64;        memory[32789] <=  8'h62;        memory[32790] <=  8'h66;        memory[32791] <=  8'h6a;        memory[32792] <=  8'h6e;        memory[32793] <=  8'h6b;        memory[32794] <=  8'h6a;        memory[32795] <=  8'h65;        memory[32796] <=  8'h38;        memory[32797] <=  8'h66;        memory[32798] <=  8'h37;        memory[32799] <=  8'h67;        memory[32800] <=  8'h79;        memory[32801] <=  8'h76;        memory[32802] <=  8'h63;        memory[32803] <=  8'h68;        memory[32804] <=  8'h69;        memory[32805] <=  8'h6a;        memory[32806] <=  8'h33;        memory[32807] <=  8'h65;        memory[32808] <=  8'h67;        memory[32809] <=  8'h79;        memory[32810] <=  8'h72;        memory[32811] <=  8'h64;        memory[32812] <=  8'h62;        memory[32813] <=  8'h6e;        memory[32814] <=  8'h63;        memory[32815] <=  8'h7a;        memory[32816] <=  8'h6a;        memory[32817] <=  8'h6f;        memory[32818] <=  8'h66;        memory[32819] <=  8'h78;        memory[32820] <=  8'h6a;        memory[32821] <=  8'h69;        memory[32822] <=  8'h63;        memory[32823] <=  8'h68;        memory[32824] <=  8'h62;        memory[32825] <=  8'h6e;        memory[32826] <=  8'h6d;        memory[32827] <=  8'h63;        memory[32828] <=  8'h73;        memory[32829] <=  8'h6c;        memory[32830] <=  8'h6b;        memory[32831] <=  8'h6a;        memory[32832] <=  8'h69;        memory[32833] <=  8'h68;        memory[32834] <=  8'h76;        memory[32835] <=  8'h75;        memory[32836] <=  8'h69;        memory[32837] <=  8'h64;        memory[32838] <=  8'h68;        memory[32839] <=  8'h75;        memory[32840] <=  8'h67;        memory[32841] <=  8'h79;        memory[32842] <=  8'h62;        memory[32843] <=  8'h68;        memory[32844] <=  8'h65;        memory[32845] <=  8'h6a;        memory[32846] <=  8'h72;        memory[32847] <=  8'h6b;        memory[32848] <=  8'h6a;        memory[32849] <=  8'h6f;        memory[32850] <=  8'h64;        memory[32851] <=  8'h67;        memory[32852] <=  8'h69;        memory[32853] <=  8'h75;        memory[32854] <=  8'h69;        memory[32855] <=  8'h67;        memory[32856] <=  8'h76;        memory[32857] <=  8'h79;        memory[32858] <=  8'h75;        memory[32859] <=  8'h67;        memory[32860] <=  8'h78;        memory[32861] <=  8'h68;        memory[32862] <=  8'h63;        memory[32863] <=  8'h20;        memory[32864] <=  8'h20;        memory[32865] <=  8'h20;        memory[32866] <=  8'h78;        memory[32867] <=  8'h76;        memory[32868] <=  8'h20;        memory[32869] <=  8'h63;        memory[32870] <=  8'h78;        memory[32871] <=  8'h67;        memory[32872] <=  8'h79;        memory[32873] <=  8'h63;        memory[32874] <=  8'h75;        memory[32875] <=  8'h68;        memory[32876] <=  8'h6a;        memory[32877] <=  8'h6b;        memory[32878] <=  8'h61;        memory[32879] <=  8'h6c;        memory[32880] <=  8'h78;        memory[32881] <=  8'h76;        memory[32882] <=  8'h70;        memory[32883] <=  8'h6f;        memory[32884] <=  8'h69;        memory[32885] <=  8'h6a;        memory[32886] <=  8'h69;        memory[32887] <=  8'h68;        memory[32888] <=  8'h6a;        memory[32889] <=  8'h62;        memory[32890] <=  8'h77;        memory[32891] <=  8'h65;        memory[32892] <=  8'h6e;        memory[32893] <=  8'h61;        memory[32894] <=  8'h66;        memory[32895] <=  8'h6d;        memory[32896] <=  8'h64;        memory[32897] <=  8'h6b;        memory[32898] <=  8'h6d;        memory[32899] <=  8'h76;        memory[32900] <=  8'h6c;        memory[32901] <=  8'h63;        memory[32902] <=  8'h6f;        memory[32903] <=  8'h64;        memory[32904] <=  8'h69;        memory[32905] <=  8'h75;        memory[32906] <=  8'h68;        memory[32907] <=  8'h73;        memory[32908] <=  8'h66;        memory[32909] <=  8'h65;        memory[32910] <=  8'h62;        memory[32911] <=  8'h6e;        memory[32912] <=  8'h64;        memory[32913] <=  8'h73;        memory[32914] <=  8'h63;        memory[32915] <=  8'h6b;        memory[32916] <=  8'h20;        memory[32917] <=  8'h78;        memory[32918] <=  8'h6a;        memory[32919] <=  8'h78;        memory[32920] <=  8'h63;        memory[32921] <=  8'h73;        memory[32922] <=  8'h64;        memory[32923] <=  8'h66;        memory[32924] <=  8'h6b;        memory[32925] <=  8'h64;        memory[32926] <=  8'h6e;        memory[32927] <=  8'h6d;        memory[32928] <=  8'h64;        memory[32929] <=  8'h73;        memory[32930] <=  8'h63;        memory[32931] <=  8'h6b;        memory[32932] <=  8'h78;        memory[32933] <=  8'h6c;        memory[32934] <=  8'h6f;        memory[32935] <=  8'h66;        memory[32936] <=  8'h6a;        memory[32937] <=  8'h69;        memory[32938] <=  8'h61;        memory[32939] <=  8'h62;        memory[32940] <=  8'h6e;        memory[32941] <=  8'h20;        memory[32942] <=  8'h78;        memory[32943] <=  8'h6b;        memory[32944] <=  8'h6d;        memory[32945] <=  8'h20;        memory[32946] <=  8'h6f;        memory[32947] <=  8'h63;        memory[32948] <=  8'h76;        memory[32949] <=  8'h73;        memory[32950] <=  8'h64;        memory[32951] <=  8'h69;        memory[32952] <=  8'h66;        memory[32953] <=  8'h68;        memory[32954] <=  8'h65;        memory[32955] <=  8'h71;        memory[32956] <=  8'h6a;        memory[32957] <=  8'h77;        memory[32958] <=  8'h62;        memory[32959] <=  8'h65;        memory[32960] <=  8'h6e;        memory[32961] <=  8'h20;        memory[32962] <=  8'h6d;        memory[32963] <=  8'h64;        memory[32964] <=  8'h73;        memory[32965] <=  8'h6c;        memory[32966] <=  8'h76;        memory[32967] <=  8'h6b;        memory[32968] <=  8'h63;        memory[32969] <=  8'h78;        memory[32970] <=  8'h20;        memory[32971] <=  8'h6f;        memory[32972] <=  8'h78;        memory[32973] <=  8'h69;        memory[32974] <=  8'h63;        memory[32975] <=  8'h6a;        memory[32976] <=  8'h76;        memory[32977] <=  8'h64;        memory[32978] <=  8'h66;        memory[32979] <=  8'h65;        memory[32980] <=  8'h71;        memory[32981] <=  8'h6e;        memory[32982] <=  8'h20;        memory[32983] <=  8'h64;        memory[32984] <=  8'h6d;        memory[32985] <=  8'h73;        memory[32986] <=  8'h6c;        memory[32987] <=  8'h63;        memory[32988] <=  8'h78;        memory[32989] <=  8'h6b;        memory[32990] <=  8'h20;        memory[32991] <=  8'h6f;        memory[32992] <=  8'h78;        memory[32993] <=  8'h63;        memory[32994] <=  8'h76;        memory[32995] <=  8'h6a;        memory[32996] <=  8'h64;        memory[32997] <=  8'h62;        memory[32998] <=  8'h71;        memory[32999] <=  8'h77;        memory[33000] <=  8'h65;        memory[33001] <=  8'h6e;        memory[33002] <=  8'h6d;        memory[33003] <=  8'h64;        memory[33004] <=  8'h6c;        memory[33005] <=  8'h73;        memory[33006] <=  8'h2c;        memory[33007] <=  8'h76;        memory[33008] <=  8'h63;        memory[33009] <=  8'h78;        memory[33010] <=  8'h20;        memory[33011] <=  8'h63;        memory[33012] <=  8'h6f;        memory[33013] <=  8'h69;        memory[33014] <=  8'h76;        memory[33015] <=  8'h68;        memory[33016] <=  8'h73;        memory[33017] <=  8'h64;        memory[33018] <=  8'h62;        memory[33019] <=  8'h71;        memory[33020] <=  8'h77;        memory[33021] <=  8'h65;        memory[33022] <=  8'h6e;        memory[33023] <=  8'h64;        memory[33024] <=  8'h6b;        memory[33025] <=  8'h73;        memory[33026] <=  8'h76;        memory[33027] <=  8'h6f;        memory[33028] <=  8'h63;        memory[33029] <=  8'h20;        memory[33030] <=  8'h76;        memory[33031] <=  8'h69;        memory[33032] <=  8'h75;        memory[33033] <=  8'h69;        memory[33034] <=  8'h68;        memory[33035] <=  8'h63;        memory[33036] <=  8'h78;        memory[33037] <=  8'h69;        memory[33038] <=  8'h6f;        memory[33039] <=  8'h76;        memory[33040] <=  8'h73;        memory[33041] <=  8'h64;        memory[33042] <=  8'h61;        memory[33043] <=  8'h64;        memory[33044] <=  8'h6e;        memory[33045] <=  8'h77;        memory[33046] <=  8'h71;        memory[33047] <=  8'h6b;        memory[33048] <=  8'h6c;        memory[33049] <=  8'h73;        memory[33050] <=  8'h76;        memory[33051] <=  8'h6e;        memory[33052] <=  8'h62;        memory[33053] <=  8'h20;        memory[33054] <=  8'h64;        memory[33055] <=  8'h66;        memory[33056] <=  8'h6a;        memory[33057] <=  8'h6b;        memory[33058] <=  8'h71;        memory[33059] <=  8'h64;        memory[33060] <=  8'h77;        memory[33061] <=  8'h65;        memory[33062] <=  8'h6e;        memory[33063] <=  8'h62;        memory[33064] <=  8'h20;        memory[33065] <=  8'h64;        memory[33066] <=  8'h73;        memory[33067] <=  8'h76;        memory[33068] <=  8'h68;        memory[33069] <=  8'h64;        memory[33070] <=  8'h61;        memory[33071] <=  8'h71;        memory[33072] <=  8'h77;        memory[33073] <=  8'h6a;        memory[33074] <=  8'h65;        memory[33075] <=  8'h6e;        memory[33076] <=  8'h64;        memory[33077] <=  8'h20;        memory[33078] <=  8'h61;        memory[33079] <=  8'h63;        memory[33080] <=  8'h62;        memory[33081] <=  8'h68;        memory[33082] <=  8'h64;        memory[33083] <=  8'h61;        memory[33084] <=  8'h77;        memory[33085] <=  8'h71;        memory[33086] <=  8'h6e;        memory[33087] <=  8'h20;        memory[33088] <=  8'h62;        memory[33089] <=  8'h73;        memory[33090] <=  8'h76;        memory[33091] <=  8'h61;        memory[33092] <=  8'h67;        memory[33093] <=  8'h76;        memory[33094] <=  8'h68;        memory[33095] <=  8'h67;        memory[33096] <=  8'h61;        memory[33097] <=  8'h73;        memory[33098] <=  8'h6a;        memory[33099] <=  8'h6b;        memory[33100] <=  8'h63;        memory[33101] <=  8'h78;        memory[33102] <=  8'h76;        memory[33103] <=  8'h6e;        memory[33104] <=  8'h73;        memory[33105] <=  8'h64;        memory[33106] <=  8'h20;        memory[33107] <=  8'h66;        memory[33108] <=  8'h62;        memory[33109] <=  8'h64;        memory[33110] <=  8'h61;        memory[33111] <=  8'h73;        memory[33112] <=  8'h76;        memory[33113] <=  8'h67;        memory[33114] <=  8'h63;        memory[33115] <=  8'h79;        memory[33116] <=  8'h7a;        memory[33117] <=  8'h78;        memory[33118] <=  8'h79;        memory[33119] <=  8'h75;        memory[33120] <=  8'h20;        memory[33121] <=  8'h69;        memory[33122] <=  8'h6a;        memory[33123] <=  8'h64;        memory[33124] <=  8'h66;        memory[33125] <=  8'h6b;        memory[33126] <=  8'h61;        memory[33127] <=  8'h64;        memory[33128] <=  8'h63;        memory[33129] <=  8'h78;        memory[33130] <=  8'h68;        memory[33131] <=  8'h20;        memory[33132] <=  8'h67;        memory[33133] <=  8'h61;        memory[33134] <=  8'h68;        memory[33135] <=  8'h75;        memory[33136] <=  8'h64;        memory[33137] <=  8'h73;        memory[33138] <=  8'h69;        memory[33139] <=  8'h6a;        memory[33140] <=  8'h61;        memory[33141] <=  8'h6b;        memory[33142] <=  8'h63;        memory[33143] <=  8'h62;        memory[33144] <=  8'h61;        memory[33145] <=  8'h72;        memory[33146] <=  8'h73;        memory[33147] <=  8'h68;        memory[33148] <=  8'h64;        memory[33149] <=  8'h66;        memory[33150] <=  8'h67;        memory[33151] <=  8'h73;        memory[33152] <=  8'h68;        memory[33153] <=  8'h64;        memory[33154] <=  8'h66;        memory[33155] <=  8'h68;        memory[33156] <=  8'h64;        memory[33157] <=  8'h6a;        memory[33158] <=  8'h68;        memory[33159] <=  8'h62;        memory[33160] <=  8'h67;        memory[33161] <=  8'h63;        memory[33162] <=  8'h61;        memory[33163] <=  8'h66;        memory[33164] <=  8'h73;        memory[33165] <=  8'h79;        memory[33166] <=  8'h67;        memory[33167] <=  8'h6b;        memory[33168] <=  8'h75;        memory[33169] <=  8'h64;        memory[33170] <=  8'h68;        memory[33171] <=  8'h62;        memory[33172] <=  8'h77;        memory[33173] <=  8'h76;        memory[33174] <=  8'h67;        memory[33175] <=  8'h61;        memory[33176] <=  8'h66;        memory[33177] <=  8'h64;        memory[33178] <=  8'h74;        memory[33179] <=  8'h75;        memory[33180] <=  8'h66;        memory[33181] <=  8'h79;        memory[33182] <=  8'h67;        memory[33183] <=  8'h69;        memory[33184] <=  8'h75;        memory[33185] <=  8'h68;        memory[33186] <=  8'h6c;        memory[33187] <=  8'h6a;        memory[33188] <=  8'h62;        memory[33189] <=  8'h6b;        memory[33190] <=  8'h68;        memory[33191] <=  8'h76;        memory[33192] <=  8'h67;        memory[33193] <=  8'h63;        memory[33194] <=  8'h66;        memory[33195] <=  8'h78;        memory[33196] <=  8'h64;        memory[33197] <=  8'h74;        memory[33198] <=  8'h75;        memory[33199] <=  8'h79;        memory[33200] <=  8'h69;        memory[33201] <=  8'h75;        memory[33202] <=  8'h68;        memory[33203] <=  8'h6c;        memory[33204] <=  8'h6a;        memory[33205] <=  8'h6b;        memory[33206] <=  8'h67;        memory[33207] <=  8'h6a;        memory[33208] <=  8'h63;        memory[33209] <=  8'h66;        memory[33210] <=  8'h68;        memory[33211] <=  8'h64;        memory[33212] <=  8'h67;        memory[33213] <=  8'h72;        memory[33214] <=  8'h79;        memory[33215] <=  8'h74;        memory[33216] <=  8'h66;        memory[33217] <=  8'h75;        memory[33218] <=  8'h79;        memory[33219] <=  8'h69;        memory[33220] <=  8'h68;        memory[33221] <=  8'h6c;        memory[33222] <=  8'h62;        memory[33223] <=  8'h6d;        memory[33224] <=  8'h76;        memory[33225] <=  8'h6e;        memory[33226] <=  8'h63;        memory[33227] <=  8'h66;        memory[33228] <=  8'h68;        memory[33229] <=  8'h64;        memory[33230] <=  8'h74;        memory[33231] <=  8'h75;        memory[33232] <=  8'h67;        memory[33233] <=  8'h79;        memory[33234] <=  8'h69;        memory[33235] <=  8'h68;        memory[33236] <=  8'h75;        memory[33237] <=  8'h6a;        memory[33238] <=  8'h6c;        memory[33239] <=  8'h62;        memory[33240] <=  8'h6d;        memory[33241] <=  8'h76;        memory[33242] <=  8'h6e;        memory[33243] <=  8'h63;        memory[33244] <=  8'h66;        memory[33245] <=  8'h68;        memory[33246] <=  8'h67;        memory[33247] <=  8'h79;        memory[33248] <=  8'h68;        memory[33249] <=  8'h75;        memory[33250] <=  8'h6a;        memory[33251] <=  8'h6e;        memory[33252] <=  8'h2c;        memory[33253] <=  8'h62;        memory[33254] <=  8'h6e;        memory[33255] <=  8'h6d;        memory[33256] <=  8'h76;        memory[33257] <=  8'h6e;        memory[33258] <=  8'h63;        memory[33259] <=  8'h66;        memory[33260] <=  8'h68;        memory[33261] <=  8'h74;        memory[33262] <=  8'h79;        memory[33263] <=  8'h69;        memory[33264] <=  8'h75;        memory[33265] <=  8'h6c;        memory[33266] <=  8'h6a;        memory[33267] <=  8'h62;        memory[33268] <=  8'h6d;        memory[33269] <=  8'h76;        memory[33270] <=  8'h6e;        memory[33271] <=  8'h63;        memory[33272] <=  8'h66;        memory[33273] <=  8'h74;        memory[33274] <=  8'h75;        memory[33275] <=  8'h79;        memory[33276] <=  8'h69;        memory[33277] <=  8'h68;        memory[33278] <=  8'h6b;        memory[33279] <=  8'h62;        memory[33280] <=  8'h76;        memory[33281] <=  8'h63;        memory[33282] <=  8'h66;        memory[33283] <=  8'h67;        memory[33284] <=  8'h74;        memory[33285] <=  8'h75;        memory[33286] <=  8'h79;        memory[33287] <=  8'h69;        memory[33288] <=  8'h75;        memory[33289] <=  8'h68;        memory[33290] <=  8'h6a;        memory[33291] <=  8'h6b;        memory[33292] <=  8'h62;        memory[33293] <=  8'h76;        memory[33294] <=  8'h63;        memory[33295] <=  8'h66;        memory[33296] <=  8'h74;        memory[33297] <=  8'h75;        memory[33298] <=  8'h79;        memory[33299] <=  8'h69;        memory[33300] <=  8'h75;        memory[33301] <=  8'h6a;        memory[33302] <=  8'h6b;        memory[33303] <=  8'h6e;        memory[33304] <=  8'h62;        memory[33305] <=  8'h76;        memory[33306] <=  8'h67;        memory[33307] <=  8'h66;        memory[33308] <=  8'h74;        memory[33309] <=  8'h79;        memory[33310] <=  8'h75;        memory[33311] <=  8'h75;        memory[33312] <=  8'h69;        memory[33313] <=  8'h6a;        memory[33314] <=  8'h6b;        memory[33315] <=  8'h68;        memory[33316] <=  8'h62;        memory[33317] <=  8'h6a;        memory[33318] <=  8'h67;        memory[33319] <=  8'h68;        memory[33320] <=  8'h66;        memory[33321] <=  8'h79;        memory[33322] <=  8'h74;        memory[33323] <=  8'h79;        memory[33324] <=  8'h69;        memory[33325] <=  8'h75;        memory[33326] <=  8'h64;        memory[33327] <=  8'h6a;        memory[33328] <=  8'h6b;        memory[33329] <=  8'h68;        memory[33330] <=  8'h63;        memory[33331] <=  8'h7a;        memory[33332] <=  8'h67;        memory[33333] <=  8'h68;        memory[33334] <=  8'h74;        memory[33335] <=  8'h75;        memory[33336] <=  8'h79;        memory[33337] <=  8'h69;        memory[33338] <=  8'h61;        memory[33339] <=  8'h73;        memory[33340] <=  8'h75;        memory[33341] <=  8'h6a;        memory[33342] <=  8'h6b;        memory[33343] <=  8'h62;        memory[33344] <=  8'h6e;        memory[33345] <=  8'h61;        memory[33346] <=  8'h76;        memory[33347] <=  8'h63;        memory[33348] <=  8'h66;        memory[33349] <=  8'h68;        memory[33350] <=  8'h75;        memory[33351] <=  8'h61;        memory[33352] <=  8'h73;        memory[33353] <=  8'h79;        memory[33354] <=  8'h64;        memory[33355] <=  8'h75;        memory[33356] <=  8'h69;        memory[33357] <=  8'h6a;        memory[33358] <=  8'h61;        memory[33359] <=  8'h6b;        memory[33360] <=  8'h62;        memory[33361] <=  8'h63;        memory[33362] <=  8'h78;        memory[33363] <=  8'h68;        memory[33364] <=  8'h67;        memory[33365] <=  8'h79;        memory[33366] <=  8'h75;        memory[33367] <=  8'h7a;        memory[33368] <=  8'h63;        memory[33369] <=  8'h61;        memory[33370] <=  8'h73;        memory[33371] <=  8'h69;        memory[33372] <=  8'h75;        memory[33373] <=  8'h6f;        memory[33374] <=  8'h69;        memory[33375] <=  8'h6a;        memory[33376] <=  8'h61;        memory[33377] <=  8'h6c;        memory[33378] <=  8'h63;        memory[33379] <=  8'h78;        memory[33380] <=  8'h62;        memory[33381] <=  8'h63;        memory[33382] <=  8'h20;        memory[33383] <=  8'h6e;        memory[33384] <=  8'h76;        memory[33385] <=  8'h63;        memory[33386] <=  8'h61;        memory[33387] <=  8'h64;        memory[33388] <=  8'h73;        memory[33389] <=  8'h67;        memory[33390] <=  8'h79;        memory[33391] <=  8'h68;        memory[33392] <=  8'h75;        memory[33393] <=  8'h61;        memory[33394] <=  8'h6a;        memory[33395] <=  8'h6b;        memory[33396] <=  8'h78;        memory[33397] <=  8'h62;        memory[33398] <=  8'h20;        memory[33399] <=  8'h6e;        memory[33400] <=  8'h76;        memory[33401] <=  8'h63;        memory[33402] <=  8'h61;        memory[33403] <=  8'h73;        memory[33404] <=  8'h67;        memory[33405] <=  8'h68;        memory[33406] <=  8'h75;        memory[33407] <=  8'h6a;        memory[33408] <=  8'h6c;        memory[33409] <=  8'h6b;        memory[33410] <=  8'h63;        memory[33411] <=  8'h78;        memory[33412] <=  8'h20;        memory[33413] <=  8'h6a;        memory[33414] <=  8'h6b;        memory[33415] <=  8'h68;        memory[33416] <=  8'h61;        memory[33417] <=  8'h73;        memory[33418] <=  8'h76;        memory[33419] <=  8'h64;        memory[33420] <=  8'h6e;        memory[33421] <=  8'h20;        memory[33422] <=  8'h62;        memory[33423] <=  8'h6e;        memory[33424] <=  8'h6d;        memory[33425] <=  8'h6b;        memory[33426] <=  8'h77;        memory[33427] <=  8'h64;        memory[33428] <=  8'h6f;        memory[33429] <=  8'h77;        memory[33430] <=  8'h69;        memory[33431] <=  8'h6f;        memory[33432] <=  8'h75;        memory[33433] <=  8'h69;        memory[33434] <=  8'h68;        memory[33435] <=  8'h62;        memory[33436] <=  8'h6e;        memory[33437] <=  8'h6b;        memory[33438] <=  8'h77;        memory[33439] <=  8'h69;        memory[33440] <=  8'h6f;        memory[33441] <=  8'h75;        memory[33442] <=  8'h71;        memory[33443] <=  8'h69;        memory[33444] <=  8'h79;        memory[33445] <=  8'h67;        memory[33446] <=  8'h6a;        memory[33447] <=  8'h64;        memory[33448] <=  8'h61;        memory[33449] <=  8'h76;        memory[33450] <=  8'h62;        memory[33451] <=  8'h6e;        memory[33452] <=  8'h6b;        memory[33453] <=  8'h6f;        memory[33454] <=  8'h70;        memory[33455] <=  8'h64;        memory[33456] <=  8'h76;        memory[33457] <=  8'h69;        memory[33458] <=  8'h6f;        memory[33459] <=  8'h75;        memory[33460] <=  8'h69;        memory[33461] <=  8'h48;        memory[33462] <=  8'h42;        memory[33463] <=  8'h6b;        memory[33464] <=  8'h64;        memory[33465] <=  8'h6e;        memory[33466] <=  8'h6c;        memory[33467] <=  8'h71;        memory[33468] <=  8'h6b;        memory[33469] <=  8'h6d;        memory[33470] <=  8'h6a;        memory[33471] <=  8'h70;        memory[33472] <=  8'h69;        memory[33473] <=  8'h6f;        memory[33474] <=  8'h68;        memory[33475] <=  8'h65;        memory[33476] <=  8'h66;        memory[33477] <=  8'h75;        memory[33478] <=  8'h67;        memory[33479] <=  8'h69;        memory[33480] <=  8'h73;        memory[33481] <=  8'h61;        memory[33482] <=  8'h62;        memory[33483] <=  8'h64;        memory[33484] <=  8'h6b;        memory[33485] <=  8'h6a;        memory[33486] <=  8'h6b;        memory[33487] <=  8'h6c;        memory[33488] <=  8'h6a;        memory[33489] <=  8'h69;        memory[33490] <=  8'h73;        memory[33491] <=  8'h6f;        memory[33492] <=  8'h71;        memory[33493] <=  8'h68;        memory[33494] <=  8'h77;        memory[33495] <=  8'h67;        memory[33496] <=  8'h69;        memory[33497] <=  8'h79;        memory[33498] <=  8'h6a;        memory[33499] <=  8'h64;        memory[33500] <=  8'h76;        memory[33501] <=  8'h62;        memory[33502] <=  8'h6e;        memory[33503] <=  8'h61;        memory[33504] <=  8'h73;        memory[33505] <=  8'h66;        memory[33506] <=  8'h6c;        memory[33507] <=  8'h6b;        memory[33508] <=  8'h64;        memory[33509] <=  8'h6a;        memory[33510] <=  8'h68;        memory[33511] <=  8'h63;        memory[33512] <=  8'h67;        memory[33513] <=  8'h6a;        memory[33514] <=  8'h76;        memory[33515] <=  8'h73;        memory[33516] <=  8'h64;        memory[33517] <=  8'h62;        memory[33518] <=  8'h62;        memory[33519] <=  8'h61;        memory[33520] <=  8'h72;        memory[33521] <=  8'h62;        memory[33522] <=  8'h62;        memory[33523] <=  8'h73;        memory[33524] <=  8'h62;        memory[33525] <=  8'h67;        memory[33526] <=  8'h73;        memory[33527] <=  8'h66;        memory[33528] <=  8'h67;        memory[33529] <=  8'h61;        memory[33530] <=  8'h68;        memory[33531] <=  8'h66;        memory[33532] <=  8'h73;        memory[33533] <=  8'h68;        memory[33534] <=  8'h61;        memory[33535] <=  8'h66;        memory[33536] <=  8'h73;        memory[33537] <=  8'h66;        memory[33538] <=  8'h68;        memory[33539] <=  8'h61;        memory[33540] <=  8'h69;        memory[33541] <=  8'h64;        memory[33542] <=  8'h75;        memory[33543] <=  8'h67;        memory[33544] <=  8'h64;        memory[33545] <=  8'h77;        memory[33546] <=  8'h62;        memory[33547] <=  8'h61;        memory[33548] <=  8'h62;        memory[33549] <=  8'h72;        memory[33550] <=  8'h62;        memory[33551] <=  8'h61;        memory[33552] <=  8'h62;        memory[33553] <=  8'h62;        memory[33554] <=  8'h74;        memory[33555] <=  8'h62;        memory[33556] <=  8'h62;        memory[33557] <=  8'h62;        memory[33558] <=  8'h62;        memory[33559] <=  8'h62;        memory[33560] <=  8'h62;        memory[33561] <=  8'h62;        memory[33562] <=  8'h62;        memory[33563] <=  8'h61;        memory[33564] <=  8'h62;        memory[33565] <=  8'h62;        memory[33566] <=  8'h72;        memory[33567] <=  8'h74;        memory[33568] <=  8'h62;        memory[33569] <=  8'h62;        memory[33570] <=  8'h61;        memory[33571] <=  8'h62;        memory[33572] <=  8'h72;        memory[33573] <=  8'h62;        memory[33574] <=  8'h74;        memory[33575] <=  8'h62;        memory[33576] <=  8'h62;        memory[33577] <=  8'h62;        memory[33578] <=  8'h63;        memory[33579] <=  8'h61;        memory[33580] <=  8'h72;        memory[33581] <=  8'h74;        memory[33582] <=  8'h73;        memory[33583] <=  8'h62;        memory[33584] <=  8'h61;        memory[33585] <=  8'h72;        memory[33586] <=  8'h74;        memory[33587] <=  8'h74;        memory[33588] <=  8'h62;        memory[33589] <=  8'h61;        memory[33590] <=  8'h72;        memory[33591] <=  8'h74;        memory[33592] <=  8'h78;        memory[33593] <=  8'h61;        memory[33594] <=  8'h74;        memory[33595] <=  8'h6b;        memory[33596] <=  8'h73;        memory[33597] <=  8'h68;        memory[33598] <=  8'h63;        memory[33599] <=  8'h66;        memory[33600] <=  8'h69;        memory[33601] <=  8'h77;        memory[33602] <=  8'h68;        memory[33603] <=  8'h61;        memory[33604] <=  8'h74;        memory[33605] <=  8'h61;        memory[33606] <=  8'h6e;        memory[33607] <=  8'h61;        memory[33608] <=  8'h62;        memory[33609] <=  8'h61;        memory[33610] <=  8'h63;        memory[33611] <=  8'h61;        memory[33612] <=  8'h74;        memory[33613] <=  8'h61;        memory[33614] <=  8'h62;        memory[33615] <=  8'h61;        memory[33616] <=  8'h72;        memory[33617] <=  8'h63;        memory[33618] <=  8'h61;        memory[33619] <=  8'h68;        memory[33620] <=  8'h64;        memory[33621] <=  8'h75;        memory[33622] <=  8'h63;        memory[33623] <=  8'h74;        memory[33624] <=  8'h61;        memory[33625] <=  8'h64;        memory[33626] <=  8'h61;        memory[33627] <=  8'h61;        memory[33628] <=  8'h63;        memory[33629] <=  8'h61;        memory[33630] <=  8'h72;        memory[33631] <=  8'h63;        memory[33632] <=  8'h74;        memory[33633] <=  8'h72;        memory[33634] <=  8'h63;        memory[33635] <=  8'h61;        memory[33636] <=  8'h74;        memory[33637] <=  8'h72;        memory[33638] <=  8'h63;        memory[33639] <=  8'h61;        memory[33640] <=  8'h74;        memory[33641] <=  8'h63;        memory[33642] <=  8'h62;        memory[33643] <=  8'h61;        memory[33644] <=  8'h74;        memory[33645] <=  8'h62;        memory[33646] <=  8'h72;        memory[33647] <=  8'h63;        memory[33648] <=  8'h61;        memory[33649] <=  8'h74;        memory[33650] <=  8'h72;        memory[33651] <=  8'h6e;        memory[33652] <=  8'h62;        memory[33653] <=  8'h61;        memory[33654] <=  8'h63;        memory[33655] <=  8'h61;        memory[33656] <=  8'h74;        memory[33657] <=  8'h79;        memory[33658] <=  8'h73;        memory[33659] <=  8'h6e;        memory[33660] <=  8'h63;        memory[33661] <=  8'h74;        memory[33662] <=  8'h61;        memory[33663] <=  8'h6e;        memory[33664] <=  8'h62;        memory[33665] <=  8'h61;        memory[33666] <=  8'h63;        memory[33667] <=  8'h72;        memory[33668] <=  8'h6e;        memory[33669] <=  8'h74;        memory[33670] <=  8'h61;        memory[33671] <=  8'h62;        memory[33672] <=  8'h74;        memory[33673] <=  8'h6e;        memory[33674] <=  8'h61;        memory[33675] <=  8'h72;        memory[33676] <=  8'h62;        memory[33677] <=  8'h78;        memory[33678] <=  8'h74;        memory[33679] <=  8'h61;        memory[33680] <=  8'h72;        memory[33681] <=  8'h62;        memory[33682] <=  8'h61;        memory[33683] <=  8'h72;        memory[33684] <=  8'h74;        memory[33685] <=  8'h74;        memory[33686] <=  8'h62;        memory[33687] <=  8'h61;        memory[33688] <=  8'h72;        memory[33689] <=  8'h74;        memory[33690] <=  8'h78;        memory[33691] <=  8'h61;        memory[33692] <=  8'h74;        memory[33693] <=  8'h6b;        memory[33694] <=  8'h73;        memory[33695] <=  8'h68;        memory[33696] <=  8'h63;        memory[33697] <=  8'h66;        memory[33698] <=  8'h69;        memory[33699] <=  8'h77;        memory[33700] <=  8'h68;        memory[33701] <=  8'h61;        memory[33702] <=  8'h74;        memory[33703] <=  8'h61;        memory[33704] <=  8'h6e;        memory[33705] <=  8'h61;        memory[33706] <=  8'h62;        memory[33707] <=  8'h61;        memory[33708] <=  8'h63;        memory[33709] <=  8'h61;        memory[33710] <=  8'h74;        memory[33711] <=  8'h61;        memory[33712] <=  8'h62;        memory[33713] <=  8'h61;        memory[33714] <=  8'h72;        memory[33715] <=  8'h63;        memory[33716] <=  8'h61;        memory[33717] <=  8'h68;        memory[33718] <=  8'h64;        memory[33719] <=  8'h75;        memory[33720] <=  8'h63;        memory[33721] <=  8'h74;        memory[33722] <=  8'h61;        memory[33723] <=  8'h64;        memory[33724] <=  8'h61;        memory[33725] <=  8'h61;        memory[33726] <=  8'h63;        memory[33727] <=  8'h61;        memory[33728] <=  8'h72;        memory[33729] <=  8'h63;        memory[33730] <=  8'h74;        memory[33731] <=  8'h72;        memory[33732] <=  8'h63;        memory[33733] <=  8'h61;        memory[33734] <=  8'h74;        memory[33735] <=  8'h72;        memory[33736] <=  8'h63;        memory[33737] <=  8'h61;        memory[33738] <=  8'h74;        memory[33739] <=  8'h63;        memory[33740] <=  8'h62;        memory[33741] <=  8'h61;        memory[33742] <=  8'h74;        memory[33743] <=  8'h62;        memory[33744] <=  8'h72;        memory[33745] <=  8'h63;        memory[33746] <=  8'h61;        memory[33747] <=  8'h74;        memory[33748] <=  8'h72;        memory[33749] <=  8'h6e;        memory[33750] <=  8'h62;        memory[33751] <=  8'h61;        memory[33752] <=  8'h63;        memory[33753] <=  8'h61;        memory[33754] <=  8'h74;        memory[33755] <=  8'h79;        memory[33756] <=  8'h73;        memory[33757] <=  8'h6e;        memory[33758] <=  8'h63;        memory[33759] <=  8'h74;        memory[33760] <=  8'h61;        memory[33761] <=  8'h6e;        memory[33762] <=  8'h62;        memory[33763] <=  8'h61;        memory[33764] <=  8'h63;        memory[33765] <=  8'h72;        memory[33766] <=  8'h6e;        memory[33767] <=  8'h74;        memory[33768] <=  8'h61;        memory[33769] <=  8'h62;        memory[33770] <=  8'h74;        memory[33771] <=  8'h6e;        memory[33772] <=  8'h61;        memory[33773] <=  8'h72;        memory[33774] <=  8'h62;        memory[33775] <=  8'h78;        memory[33776] <=  8'h74;        memory[33777] <=  8'h61;        memory[33778] <=  8'h72;        memory[33779] <=  8'h62;        memory[33780] <=  8'h61;        memory[33781] <=  8'h72;        memory[33782] <=  8'h74;        memory[33783] <=  8'h74;        memory[33784] <=  8'h62;        memory[33785] <=  8'h61;        memory[33786] <=  8'h72;        memory[33787] <=  8'h74;        memory[33788] <=  8'h78;        memory[33789] <=  8'h61;        memory[33790] <=  8'h74;        memory[33791] <=  8'h6b;        memory[33792] <=  8'h73;        memory[33793] <=  8'h68;        memory[33794] <=  8'h63;        memory[33795] <=  8'h66;        memory[33796] <=  8'h69;        memory[33797] <=  8'h77;        memory[33798] <=  8'h68;        memory[33799] <=  8'h61;        memory[33800] <=  8'h74;        memory[33801] <=  8'h61;        memory[33802] <=  8'h6e;        memory[33803] <=  8'h61;        memory[33804] <=  8'h62;        memory[33805] <=  8'h61;        memory[33806] <=  8'h63;        memory[33807] <=  8'h61;        memory[33808] <=  8'h74;        memory[33809] <=  8'h61;        memory[33810] <=  8'h62;        memory[33811] <=  8'h61;        memory[33812] <=  8'h72;        memory[33813] <=  8'h63;        memory[33814] <=  8'h61;        memory[33815] <=  8'h68;        memory[33816] <=  8'h64;        memory[33817] <=  8'h75;        memory[33818] <=  8'h63;        memory[33819] <=  8'h74;        memory[33820] <=  8'h61;        memory[33821] <=  8'h64;        memory[33822] <=  8'h61;        memory[33823] <=  8'h61;        memory[33824] <=  8'h63;        memory[33825] <=  8'h61;        memory[33826] <=  8'h72;        memory[33827] <=  8'h63;        memory[33828] <=  8'h74;        memory[33829] <=  8'h72;        memory[33830] <=  8'h63;        memory[33831] <=  8'h61;        memory[33832] <=  8'h74;        memory[33833] <=  8'h72;        memory[33834] <=  8'h63;        memory[33835] <=  8'h61;        memory[33836] <=  8'h74;        memory[33837] <=  8'h63;        memory[33838] <=  8'h62;        memory[33839] <=  8'h61;        memory[33840] <=  8'h74;        memory[33841] <=  8'h62;        memory[33842] <=  8'h72;        memory[33843] <=  8'h63;        memory[33844] <=  8'h61;        memory[33845] <=  8'h74;        memory[33846] <=  8'h72;        memory[33847] <=  8'h6e;        memory[33848] <=  8'h62;        memory[33849] <=  8'h61;        memory[33850] <=  8'h63;        memory[33851] <=  8'h61;        memory[33852] <=  8'h74;        memory[33853] <=  8'h79;        memory[33854] <=  8'h73;        memory[33855] <=  8'h6e;        memory[33856] <=  8'h63;        memory[33857] <=  8'h74;        memory[33858] <=  8'h61;        memory[33859] <=  8'h6e;        memory[33860] <=  8'h62;        memory[33861] <=  8'h61;        memory[33862] <=  8'h63;        memory[33863] <=  8'h72;        memory[33864] <=  8'h6e;        memory[33865] <=  8'h74;        memory[33866] <=  8'h61;        memory[33867] <=  8'h62;        memory[33868] <=  8'h74;        memory[33869] <=  8'h6e;        memory[33870] <=  8'h61;        memory[33871] <=  8'h72;        memory[33872] <=  8'h62;        memory[33873] <=  8'h78;        memory[33874] <=  8'h74;        memory[33875] <=  8'h61;        memory[33876] <=  8'h72;        memory[33877] <=  8'h5d;        memory[33878] <=  8'h5d;        memory[33879] <=  8'h65;        memory[33880] <=  8'h66;        memory[33881] <=  8'h77;        memory[33882] <=  8'h65;        memory[33883] <=  8'h5d;        memory[33884] <=  8'h65;        memory[33885] <=  8'h67;        memory[33886] <=  8'h73;        memory[33887] <=  8'h67;        memory[33888] <=  8'h66;        memory[33889] <=  8'h62;        memory[33890] <=  8'h61;        memory[33891] <=  8'h72;        memory[33892] <=  8'h74;        memory[33893] <=  8'h74;        memory[33894] <=  8'h62;        memory[33895] <=  8'h61;        memory[33896] <=  8'h72;        memory[33897] <=  8'h74;        memory[33898] <=  8'h78;        memory[33899] <=  8'h61;        memory[33900] <=  8'h74;        memory[33901] <=  8'h6b;        memory[33902] <=  8'h73;        memory[33903] <=  8'h68;        memory[33904] <=  8'h63;        memory[33905] <=  8'h66;        memory[33906] <=  8'h69;        memory[33907] <=  8'h77;        memory[33908] <=  8'h68;        memory[33909] <=  8'h61;        memory[33910] <=  8'h74;        memory[33911] <=  8'h61;        memory[33912] <=  8'h6e;        memory[33913] <=  8'h61;        memory[33914] <=  8'h62;        memory[33915] <=  8'h61;        memory[33916] <=  8'h63;        memory[33917] <=  8'h61;        memory[33918] <=  8'h74;        memory[33919] <=  8'h61;        memory[33920] <=  8'h62;        memory[33921] <=  8'h61;        memory[33922] <=  8'h72;        memory[33923] <=  8'h63;        memory[33924] <=  8'h61;        memory[33925] <=  8'h68;        memory[33926] <=  8'h64;        memory[33927] <=  8'h75;        memory[33928] <=  8'h63;        memory[33929] <=  8'h74;        memory[33930] <=  8'h61;        memory[33931] <=  8'h64;        memory[33932] <=  8'h61;        memory[33933] <=  8'h61;        memory[33934] <=  8'h63;        memory[33935] <=  8'h61;        memory[33936] <=  8'h72;        memory[33937] <=  8'h63;        memory[33938] <=  8'h74;        memory[33939] <=  8'h72;        memory[33940] <=  8'h63;        memory[33941] <=  8'h61;        memory[33942] <=  8'h74;        memory[33943] <=  8'h72;        memory[33944] <=  8'h63;        memory[33945] <=  8'h61;        memory[33946] <=  8'h74;        memory[33947] <=  8'h63;        memory[33948] <=  8'h62;        memory[33949] <=  8'h61;        memory[33950] <=  8'h74;        memory[33951] <=  8'h62;        memory[33952] <=  8'h72;        memory[33953] <=  8'h63;        memory[33954] <=  8'h61;        memory[33955] <=  8'h74;        memory[33956] <=  8'h72;        memory[33957] <=  8'h6e;        memory[33958] <=  8'h62;        memory[33959] <=  8'h61;        memory[33960] <=  8'h63;        memory[33961] <=  8'h61;        memory[33962] <=  8'h74;        memory[33963] <=  8'h79;        memory[33964] <=  8'h73;        memory[33965] <=  8'h6e;        memory[33966] <=  8'h63;        memory[33967] <=  8'h74;        memory[33968] <=  8'h61;        memory[33969] <=  8'h6e;        memory[33970] <=  8'h62;        memory[33971] <=  8'h61;        memory[33972] <=  8'h63;        memory[33973] <=  8'h72;        memory[33974] <=  8'h6e;        memory[33975] <=  8'h74;        memory[33976] <=  8'h61;        memory[33977] <=  8'h62;        memory[33978] <=  8'h74;        memory[33979] <=  8'h6e;        memory[33980] <=  8'h61;        memory[33981] <=  8'h72;        memory[33982] <=  8'h62;        memory[33983] <=  8'h78;        memory[33984] <=  8'h74;        memory[33985] <=  8'h61;        memory[33986] <=  8'h72;        memory[33987] <=  8'h62;        memory[33988] <=  8'h61;        memory[33989] <=  8'h72;        memory[33990] <=  8'h74;        memory[33991] <=  8'h74;        memory[33992] <=  8'h62;        memory[33993] <=  8'h61;        memory[33994] <=  8'h72;        memory[33995] <=  8'h74;        memory[33996] <=  8'h78;        memory[33997] <=  8'h61;        memory[33998] <=  8'h74;        memory[33999] <=  8'h6b;        memory[34000] <=  8'h73;        memory[34001] <=  8'h68;        memory[34002] <=  8'h63;        memory[34003] <=  8'h66;        memory[34004] <=  8'h69;        memory[34005] <=  8'h77;        memory[34006] <=  8'h68;        memory[34007] <=  8'h61;        memory[34008] <=  8'h74;        memory[34009] <=  8'h61;        memory[34010] <=  8'h6e;        memory[34011] <=  8'h61;        memory[34012] <=  8'h62;        memory[34013] <=  8'h61;        memory[34014] <=  8'h63;        memory[34015] <=  8'h61;        memory[34016] <=  8'h74;        memory[34017] <=  8'h61;        memory[34018] <=  8'h62;        memory[34019] <=  8'h61;        memory[34020] <=  8'h72;        memory[34021] <=  8'h63;        memory[34022] <=  8'h61;        memory[34023] <=  8'h68;        memory[34024] <=  8'h64;        memory[34025] <=  8'h75;        memory[34026] <=  8'h63;        memory[34027] <=  8'h74;        memory[34028] <=  8'h61;        memory[34029] <=  8'h64;        memory[34030] <=  8'h61;        memory[34031] <=  8'h61;        memory[34032] <=  8'h63;        memory[34033] <=  8'h61;        memory[34034] <=  8'h72;        memory[34035] <=  8'h63;        memory[34036] <=  8'h74;        memory[34037] <=  8'h72;        memory[34038] <=  8'h63;        memory[34039] <=  8'h61;        memory[34040] <=  8'h74;        memory[34041] <=  8'h72;        memory[34042] <=  8'h63;        memory[34043] <=  8'h61;        memory[34044] <=  8'h74;        memory[34045] <=  8'h63;        memory[34046] <=  8'h62;        memory[34047] <=  8'h61;        memory[34048] <=  8'h74;        memory[34049] <=  8'h62;        memory[34050] <=  8'h72;        memory[34051] <=  8'h63;        memory[34052] <=  8'h61;        memory[34053] <=  8'h74;        memory[34054] <=  8'h72;        memory[34055] <=  8'h6e;        memory[34056] <=  8'h62;        memory[34057] <=  8'h61;        memory[34058] <=  8'h63;        memory[34059] <=  8'h61;        memory[34060] <=  8'h74;        memory[34061] <=  8'h79;        memory[34062] <=  8'h73;        memory[34063] <=  8'h6e;        memory[34064] <=  8'h63;        memory[34065] <=  8'h74;        memory[34066] <=  8'h61;        memory[34067] <=  8'h6e;        memory[34068] <=  8'h62;        memory[34069] <=  8'h61;        memory[34070] <=  8'h63;        memory[34071] <=  8'h72;        memory[34072] <=  8'h6e;        memory[34073] <=  8'h74;        memory[34074] <=  8'h61;        memory[34075] <=  8'h62;        memory[34076] <=  8'h74;        memory[34077] <=  8'h6e;        memory[34078] <=  8'h61;        memory[34079] <=  8'h72;        memory[34080] <=  8'h62;        memory[34081] <=  8'h78;        memory[34082] <=  8'h74;        memory[34083] <=  8'h61;        memory[34084] <=  8'h72;        memory[34085] <=  8'h64;        memory[34086] <=  8'h66;        memory[34087] <=  8'h73;        memory[34088] <=  8'h67;        memory[34089] <=  8'h76;        memory[34090] <=  8'h68;        memory[34091] <=  8'h62;        memory[34092] <=  8'h6b;        memory[34093] <=  8'h6a;        memory[34094] <=  8'h6e;        memory[34095] <=  8'h6d;        memory[34096] <=  8'h62;        memory[34097] <=  8'h76;        memory[34098] <=  8'h78;        memory[34099] <=  8'h63;        memory[34100] <=  8'h73;        memory[34101] <=  8'h66;        memory[34102] <=  8'h72;        memory[34103] <=  8'h74;        memory[34104] <=  8'h79;        memory[34105] <=  8'h75;        memory[34106] <=  8'h6a;        memory[34107] <=  8'h6e;        memory[34108] <=  8'h62;        memory[34109] <=  8'h76;        memory[34110] <=  8'h63;        memory[34111] <=  8'h64;        memory[34112] <=  8'h74;        memory[34113] <=  8'h79;        memory[34114] <=  8'h75;        memory[34115] <=  8'h69;        memory[34116] <=  8'h6b;        memory[34117] <=  8'h6d;        memory[34118] <=  8'h6e;        memory[34119] <=  8'h62;        memory[34120] <=  8'h76;        memory[34121] <=  8'h63;        memory[34122] <=  8'h78;        memory[34123] <=  8'h73;        memory[34124] <=  8'h64;        memory[34125] <=  8'h72;        memory[34126] <=  8'h74;        memory[34127] <=  8'h79;        memory[34128] <=  8'h75;        memory[34129] <=  8'h69;        memory[34130] <=  8'h6b;        memory[34131] <=  8'h6d;        memory[34132] <=  8'h6e;        memory[34133] <=  8'h62;        memory[34134] <=  8'h76;        memory[34135] <=  8'h63;        memory[34136] <=  8'h73;        memory[34137] <=  8'h77;        memory[34138] <=  8'h33;        memory[34139] <=  8'h34;        memory[34140] <=  8'h35;        memory[34141] <=  8'h36;        memory[34142] <=  8'h37;        memory[34143] <=  8'h38;        memory[34144] <=  8'h69;        memory[34145] <=  8'h6b;        memory[34146] <=  8'h6d;        memory[34147] <=  8'h6e;        memory[34148] <=  8'h62;        memory[34149] <=  8'h76;        memory[34150] <=  8'h63;        memory[34151] <=  8'h64;        memory[34152] <=  8'h65;        memory[34153] <=  8'h72;        memory[34154] <=  8'h36;        memory[34155] <=  8'h37;        memory[34156] <=  8'h38;        memory[34157] <=  8'h69;        memory[34158] <=  8'h6f;        memory[34159] <=  8'h6b;        memory[34160] <=  8'h6a;        memory[34161] <=  8'h6e;        memory[34162] <=  8'h62;        memory[34163] <=  8'h76;        memory[34164] <=  8'h63;        memory[34165] <=  8'h64;        memory[34166] <=  8'h72;        memory[34167] <=  8'h74;        memory[34168] <=  8'h79;        memory[34169] <=  8'h75;        memory[34170] <=  8'h73;        memory[34171] <=  8'h6a;        memory[34172] <=  8'h63;        memory[34173] <=  8'h6e;        memory[34174] <=  8'h62;        memory[34175] <=  8'h64;        memory[34176] <=  8'h66;        memory[34177] <=  8'h73;        memory[34178] <=  8'h74;        memory[34179] <=  8'h79;        memory[34180] <=  8'h75;        memory[34181] <=  8'h61;        memory[34182] <=  8'h69;        memory[34183] <=  8'h6b;        memory[34184] <=  8'h78;        memory[34185] <=  8'h6d;        memory[34186] <=  8'h6e;        memory[34187] <=  8'h73;        memory[34188] <=  8'h6a;        memory[34189] <=  8'h6f;        memory[34190] <=  8'h64;        memory[34191] <=  8'h6c;        memory[34192] <=  8'h63;        memory[34193] <=  8'h78;        memory[34194] <=  8'h62;        memory[34195] <=  8'h61;        memory[34196] <=  8'h72;        memory[34197] <=  8'h74;        memory[34198] <=  8'h78;        memory[34199] <=  8'h61;        memory[34200] <=  8'h74;        memory[34201] <=  8'h6b;        memory[34202] <=  8'h73;        memory[34203] <=  8'h68;        memory[34204] <=  8'h63;        memory[34205] <=  8'h66;        memory[34206] <=  8'h69;        memory[34207] <=  8'h77;        memory[34208] <=  8'h68;        memory[34209] <=  8'h61;        memory[34210] <=  8'h74;        memory[34211] <=  8'h61;        memory[34212] <=  8'h6e;        memory[34213] <=  8'h61;        memory[34214] <=  8'h62;        memory[34215] <=  8'h61;        memory[34216] <=  8'h63;        memory[34217] <=  8'h61;        memory[34218] <=  8'h74;        memory[34219] <=  8'h61;        memory[34220] <=  8'h62;        memory[34221] <=  8'h61;        memory[34222] <=  8'h72;        memory[34223] <=  8'h63;        memory[34224] <=  8'h61;        memory[34225] <=  8'h68;        memory[34226] <=  8'h64;        memory[34227] <=  8'h75;        memory[34228] <=  8'h63;        memory[34229] <=  8'h74;        memory[34230] <=  8'h61;        memory[34231] <=  8'h64;        memory[34232] <=  8'h61;        memory[34233] <=  8'h61;        memory[34234] <=  8'h63;        memory[34235] <=  8'h61;        memory[34236] <=  8'h72;        memory[34237] <=  8'h62;        memory[34238] <=  8'h61;        memory[34239] <=  8'h72;        memory[34240] <=  8'h74;        memory[34241] <=  8'h78;        memory[34242] <=  8'h61;        memory[34243] <=  8'h74;        memory[34244] <=  8'h6b;        memory[34245] <=  8'h73;        memory[34246] <=  8'h68;        memory[34247] <=  8'h63;        memory[34248] <=  8'h66;        memory[34249] <=  8'h69;        memory[34250] <=  8'h77;        memory[34251] <=  8'h68;        memory[34252] <=  8'h61;        memory[34253] <=  8'h74;        memory[34254] <=  8'h61;        memory[34255] <=  8'h6e;        memory[34256] <=  8'h61;        memory[34257] <=  8'h62;        memory[34258] <=  8'h61;        memory[34259] <=  8'h63;        memory[34260] <=  8'h61;        memory[34261] <=  8'h74;        memory[34262] <=  8'h61;        memory[34263] <=  8'h62;        memory[34264] <=  8'h61;        memory[34265] <=  8'h72;        memory[34266] <=  8'h63;        memory[34267] <=  8'h61;        memory[34268] <=  8'h68;        memory[34269] <=  8'h64;        memory[34270] <=  8'h75;        memory[34271] <=  8'h63;        memory[34272] <=  8'h74;        memory[34273] <=  8'h61;        memory[34274] <=  8'h64;        memory[34275] <=  8'h61;        memory[34276] <=  8'h61;        memory[34277] <=  8'h63;        memory[34278] <=  8'h61;        memory[34279] <=  8'h72;        memory[34280] <=  8'h62;        memory[34281] <=  8'h61;        memory[34282] <=  8'h72;        memory[34283] <=  8'h74;        memory[34284] <=  8'h78;        memory[34285] <=  8'h61;        memory[34286] <=  8'h74;        memory[34287] <=  8'h6b;        memory[34288] <=  8'h73;        memory[34289] <=  8'h68;        memory[34290] <=  8'h63;        memory[34291] <=  8'h66;        memory[34292] <=  8'h69;        memory[34293] <=  8'h77;        memory[34294] <=  8'h68;        memory[34295] <=  8'h61;        memory[34296] <=  8'h74;        memory[34297] <=  8'h61;        memory[34298] <=  8'h6e;        memory[34299] <=  8'h61;        memory[34300] <=  8'h62;        memory[34301] <=  8'h61;        memory[34302] <=  8'h63;        memory[34303] <=  8'h61;        memory[34304] <=  8'h74;        memory[34305] <=  8'h61;        memory[34306] <=  8'h62;        memory[34307] <=  8'h61;        memory[34308] <=  8'h72;        memory[34309] <=  8'h63;        memory[34310] <=  8'h61;        memory[34311] <=  8'h68;        memory[34312] <=  8'h64;        memory[34313] <=  8'h75;        memory[34314] <=  8'h63;        memory[34315] <=  8'h74;        memory[34316] <=  8'h61;        memory[34317] <=  8'h64;        memory[34318] <=  8'h61;        memory[34319] <=  8'h61;        memory[34320] <=  8'h63;        memory[34321] <=  8'h61;        memory[34322] <=  8'h72;        memory[34323] <=  8'h62;        memory[34324] <=  8'h61;        memory[34325] <=  8'h72;        memory[34326] <=  8'h74;        memory[34327] <=  8'h78;        memory[34328] <=  8'h61;        memory[34329] <=  8'h74;        memory[34330] <=  8'h6b;        memory[34331] <=  8'h73;        memory[34332] <=  8'h68;        memory[34333] <=  8'h63;        memory[34334] <=  8'h66;        memory[34335] <=  8'h69;        memory[34336] <=  8'h77;        memory[34337] <=  8'h68;        memory[34338] <=  8'h61;        memory[34339] <=  8'h74;        memory[34340] <=  8'h61;        memory[34341] <=  8'h6e;        memory[34342] <=  8'h61;        memory[34343] <=  8'h62;        memory[34344] <=  8'h61;        memory[34345] <=  8'h63;        memory[34346] <=  8'h61;        memory[34347] <=  8'h74;        memory[34348] <=  8'h61;        memory[34349] <=  8'h62;        memory[34350] <=  8'h61;        memory[34351] <=  8'h72;        memory[34352] <=  8'h63;        memory[34353] <=  8'h61;        memory[34354] <=  8'h68;        memory[34355] <=  8'h64;        memory[34356] <=  8'h75;        memory[34357] <=  8'h63;        memory[34358] <=  8'h74;        memory[34359] <=  8'h61;        memory[34360] <=  8'h64;        memory[34361] <=  8'h61;        memory[34362] <=  8'h61;        memory[34363] <=  8'h63;        memory[34364] <=  8'h61;        memory[34365] <=  8'h72;        memory[34366] <=  8'h62;        memory[34367] <=  8'h61;        memory[34368] <=  8'h72;        memory[34369] <=  8'h74;        memory[34370] <=  8'h78;        memory[34371] <=  8'h61;        memory[34372] <=  8'h74;        memory[34373] <=  8'h6b;        memory[34374] <=  8'h73;        memory[34375] <=  8'h68;        memory[34376] <=  8'h63;        memory[34377] <=  8'h66;        memory[34378] <=  8'h69;        memory[34379] <=  8'h77;        memory[34380] <=  8'h68;        memory[34381] <=  8'h61;        memory[34382] <=  8'h74;        memory[34383] <=  8'h61;        memory[34384] <=  8'h6e;        memory[34385] <=  8'h61;        memory[34386] <=  8'h62;        memory[34387] <=  8'h61;        memory[34388] <=  8'h63;        memory[34389] <=  8'h61;        memory[34390] <=  8'h74;        memory[34391] <=  8'h61;        memory[34392] <=  8'h62;        memory[34393] <=  8'h61;        memory[34394] <=  8'h72;        memory[34395] <=  8'h63;        memory[34396] <=  8'h61;        memory[34397] <=  8'h68;        memory[34398] <=  8'h64;        memory[34399] <=  8'h75;        memory[34400] <=  8'h63;        memory[34401] <=  8'h74;        memory[34402] <=  8'h61;        memory[34403] <=  8'h64;        memory[34404] <=  8'h61;        memory[34405] <=  8'h61;        memory[34406] <=  8'h63;        memory[34407] <=  8'h61;        memory[34408] <=  8'h72;        memory[34409] <=  8'h62;        memory[34410] <=  8'h61;        memory[34411] <=  8'h72;        memory[34412] <=  8'h74;        memory[34413] <=  8'h78;        memory[34414] <=  8'h61;        memory[34415] <=  8'h74;        memory[34416] <=  8'h6b;        memory[34417] <=  8'h73;        memory[34418] <=  8'h68;        memory[34419] <=  8'h63;        memory[34420] <=  8'h66;        memory[34421] <=  8'h69;        memory[34422] <=  8'h77;        memory[34423] <=  8'h68;        memory[34424] <=  8'h61;        memory[34425] <=  8'h74;        memory[34426] <=  8'h61;        memory[34427] <=  8'h6e;        memory[34428] <=  8'h61;        memory[34429] <=  8'h62;        memory[34430] <=  8'h61;        memory[34431] <=  8'h63;        memory[34432] <=  8'h61;        memory[34433] <=  8'h74;        memory[34434] <=  8'h61;        memory[34435] <=  8'h62;        memory[34436] <=  8'h61;        memory[34437] <=  8'h72;        memory[34438] <=  8'h63;        memory[34439] <=  8'h61;        memory[34440] <=  8'h68;        memory[34441] <=  8'h64;        memory[34442] <=  8'h75;        memory[34443] <=  8'h63;        memory[34444] <=  8'h74;        memory[34445] <=  8'h61;        memory[34446] <=  8'h64;        memory[34447] <=  8'h61;        memory[34448] <=  8'h61;        memory[34449] <=  8'h63;        memory[34450] <=  8'h61;        memory[34451] <=  8'h72;        memory[34452] <=  8'h62;        memory[34453] <=  8'h61;        memory[34454] <=  8'h72;        memory[34455] <=  8'h74;        memory[34456] <=  8'h78;        memory[34457] <=  8'h61;        memory[34458] <=  8'h74;        memory[34459] <=  8'h6b;        memory[34460] <=  8'h73;        memory[34461] <=  8'h68;        memory[34462] <=  8'h63;        memory[34463] <=  8'h66;        memory[34464] <=  8'h69;        memory[34465] <=  8'h77;        memory[34466] <=  8'h68;        memory[34467] <=  8'h61;        memory[34468] <=  8'h74;        memory[34469] <=  8'h61;        memory[34470] <=  8'h6e;        memory[34471] <=  8'h61;        memory[34472] <=  8'h62;        memory[34473] <=  8'h61;        memory[34474] <=  8'h63;        memory[34475] <=  8'h61;        memory[34476] <=  8'h74;        memory[34477] <=  8'h61;        memory[34478] <=  8'h62;        memory[34479] <=  8'h61;        memory[34480] <=  8'h72;        memory[34481] <=  8'h63;        memory[34482] <=  8'h61;        memory[34483] <=  8'h68;        memory[34484] <=  8'h64;        memory[34485] <=  8'h75;        memory[34486] <=  8'h63;        memory[34487] <=  8'h74;        memory[34488] <=  8'h61;        memory[34489] <=  8'h64;        memory[34490] <=  8'h61;        memory[34491] <=  8'h61;        memory[34492] <=  8'h63;        memory[34493] <=  8'h61;        memory[34494] <=  8'h72;        memory[34495] <=  8'h62;        memory[34496] <=  8'h61;        memory[34497] <=  8'h72;        memory[34498] <=  8'h74;        memory[34499] <=  8'h78;        memory[34500] <=  8'h61;        memory[34501] <=  8'h74;        memory[34502] <=  8'h6b;        memory[34503] <=  8'h73;        memory[34504] <=  8'h68;        memory[34505] <=  8'h63;        memory[34506] <=  8'h66;        memory[34507] <=  8'h69;        memory[34508] <=  8'h77;        memory[34509] <=  8'h68;        memory[34510] <=  8'h61;        memory[34511] <=  8'h74;        memory[34512] <=  8'h61;        memory[34513] <=  8'h6e;        memory[34514] <=  8'h61;        memory[34515] <=  8'h62;        memory[34516] <=  8'h61;        memory[34517] <=  8'h63;        memory[34518] <=  8'h61;        memory[34519] <=  8'h74;        memory[34520] <=  8'h61;        memory[34521] <=  8'h62;        memory[34522] <=  8'h61;        memory[34523] <=  8'h72;        memory[34524] <=  8'h63;        memory[34525] <=  8'h61;        memory[34526] <=  8'h68;        memory[34527] <=  8'h64;        memory[34528] <=  8'h75;        memory[34529] <=  8'h63;        memory[34530] <=  8'h74;        memory[34531] <=  8'h61;        memory[34532] <=  8'h64;        memory[34533] <=  8'h61;        memory[34534] <=  8'h61;        memory[34535] <=  8'h63;        memory[34536] <=  8'h61;        memory[34537] <=  8'h72;        memory[34538] <=  8'h62;        memory[34539] <=  8'h61;        memory[34540] <=  8'h72;        memory[34541] <=  8'h74;        memory[34542] <=  8'h78;        memory[34543] <=  8'h61;        memory[34544] <=  8'h74;        memory[34545] <=  8'h6b;        memory[34546] <=  8'h73;        memory[34547] <=  8'h68;        memory[34548] <=  8'h63;        memory[34549] <=  8'h66;        memory[34550] <=  8'h69;        memory[34551] <=  8'h77;        memory[34552] <=  8'h68;        memory[34553] <=  8'h61;        memory[34554] <=  8'h74;        memory[34555] <=  8'h61;        memory[34556] <=  8'h6e;        memory[34557] <=  8'h61;        memory[34558] <=  8'h62;        memory[34559] <=  8'h61;        memory[34560] <=  8'h63;        memory[34561] <=  8'h61;        memory[34562] <=  8'h74;        memory[34563] <=  8'h61;        memory[34564] <=  8'h62;        memory[34565] <=  8'h61;        memory[34566] <=  8'h72;        memory[34567] <=  8'h63;        memory[34568] <=  8'h61;        memory[34569] <=  8'h68;        memory[34570] <=  8'h64;        memory[34571] <=  8'h75;        memory[34572] <=  8'h63;        memory[34573] <=  8'h74;        memory[34574] <=  8'h61;        memory[34575] <=  8'h64;        memory[34576] <=  8'h61;        memory[34577] <=  8'h61;        memory[34578] <=  8'h63;        memory[34579] <=  8'h61;        memory[34580] <=  8'h72;        memory[34581] <=  8'h62;        memory[34582] <=  8'h61;        memory[34583] <=  8'h72;        memory[34584] <=  8'h74;        memory[34585] <=  8'h74;        memory[34586] <=  8'h62;        memory[34587] <=  8'h61;        memory[34588] <=  8'h72;        memory[34589] <=  8'h74;        memory[34590] <=  8'h78;        memory[34591] <=  8'h61;        memory[34592] <=  8'h74;        memory[34593] <=  8'h6b;        memory[34594] <=  8'h73;        memory[34595] <=  8'h68;        memory[34596] <=  8'h63;        memory[34597] <=  8'h66;        memory[34598] <=  8'h69;        memory[34599] <=  8'h77;        memory[34600] <=  8'h68;        memory[34601] <=  8'h61;        memory[34602] <=  8'h74;        memory[34603] <=  8'h61;        memory[34604] <=  8'h6e;        memory[34605] <=  8'h61;        memory[34606] <=  8'h62;        memory[34607] <=  8'h61;        memory[34608] <=  8'h63;        memory[34609] <=  8'h61;        memory[34610] <=  8'h74;        memory[34611] <=  8'h61;        memory[34612] <=  8'h62;        memory[34613] <=  8'h61;        memory[34614] <=  8'h72;        memory[34615] <=  8'h63;        memory[34616] <=  8'h61;        memory[34617] <=  8'h68;        memory[34618] <=  8'h64;        memory[34619] <=  8'h75;        memory[34620] <=  8'h63;        memory[34621] <=  8'h74;        memory[34622] <=  8'h61;        memory[34623] <=  8'h64;        memory[34624] <=  8'h61;        memory[34625] <=  8'h61;        memory[34626] <=  8'h63;        memory[34627] <=  8'h61;        memory[34628] <=  8'h72;        memory[34629] <=  8'h63;        memory[34630] <=  8'h74;        memory[34631] <=  8'h72;        memory[34632] <=  8'h63;        memory[34633] <=  8'h61;        memory[34634] <=  8'h74;        memory[34635] <=  8'h72;        memory[34636] <=  8'h63;        memory[34637] <=  8'h61;        memory[34638] <=  8'h74;        memory[34639] <=  8'h63;        memory[34640] <=  8'h62;        memory[34641] <=  8'h61;        memory[34642] <=  8'h74;        memory[34643] <=  8'h62;        memory[34644] <=  8'h72;        memory[34645] <=  8'h63;        memory[34646] <=  8'h61;        memory[34647] <=  8'h72;        memory[34648] <=  8'h62;        memory[34649] <=  8'h78;        memory[34650] <=  8'h74;        memory[34651] <=  8'h61;        memory[34652] <=  8'h72;        memory[34653] <=  8'h64;        memory[34654] <=  8'h66;        memory[34655] <=  8'h73;        memory[34656] <=  8'h67;        memory[34657] <=  8'h76;        memory[34658] <=  8'h68;        memory[34659] <=  8'h62;        memory[34660] <=  8'h6b;        memory[34661] <=  8'h6a;        memory[34662] <=  8'h6e;        memory[34663] <=  8'h6d;        memory[34664] <=  8'h62;        memory[34665] <=  8'h76;        memory[34666] <=  8'h78;        memory[34667] <=  8'h63;        memory[34668] <=  8'h73;        memory[34669] <=  8'h66;        memory[34670] <=  8'h72;        memory[34671] <=  8'h74;        memory[34672] <=  8'h79;        memory[34673] <=  8'h75;        memory[34674] <=  8'h6a;        memory[34675] <=  8'h6e;        memory[34676] <=  8'h62;        memory[34677] <=  8'h76;        memory[34678] <=  8'h63;        memory[34679] <=  8'h64;        memory[34680] <=  8'h74;        memory[34681] <=  8'h79;        memory[34682] <=  8'h75;        memory[34683] <=  8'h69;        memory[34684] <=  8'h6b;        memory[34685] <=  8'h6d;        memory[34686] <=  8'h6e;        memory[34687] <=  8'h62;        memory[34688] <=  8'h76;        memory[34689] <=  8'h63;        memory[34690] <=  8'h78;        memory[34691] <=  8'h73;        memory[34692] <=  8'h64;        memory[34693] <=  8'h72;        memory[34694] <=  8'h74;        memory[34695] <=  8'h79;        memory[34696] <=  8'h75;        memory[34697] <=  8'h69;        memory[34698] <=  8'h6b;        memory[34699] <=  8'h6d;        memory[34700] <=  8'h6e;        memory[34701] <=  8'h62;        memory[34702] <=  8'h76;        memory[34703] <=  8'h63;        memory[34704] <=  8'h73;        memory[34705] <=  8'h77;        memory[34706] <=  8'h33;        memory[34707] <=  8'h34;        memory[34708] <=  8'h35;        memory[34709] <=  8'h36;        memory[34710] <=  8'h37;        memory[34711] <=  8'h38;        memory[34712] <=  8'h69;        memory[34713] <=  8'h6b;        memory[34714] <=  8'h6d;        memory[34715] <=  8'h6e;        memory[34716] <=  8'h62;        memory[34717] <=  8'h76;        memory[34718] <=  8'h63;        memory[34719] <=  8'h64;        memory[34720] <=  8'h65;        memory[34721] <=  8'h72;        memory[34722] <=  8'h36;        memory[34723] <=  8'h37;        memory[34724] <=  8'h38;        memory[34725] <=  8'h69;        memory[34726] <=  8'h6f;        memory[34727] <=  8'h6b;        memory[34728] <=  8'h6a;        memory[34729] <=  8'h6e;        memory[34730] <=  8'h62;        memory[34731] <=  8'h76;        memory[34732] <=  8'h63;        memory[34733] <=  8'h64;        memory[34734] <=  8'h72;        memory[34735] <=  8'h74;        memory[34736] <=  8'h79;        memory[34737] <=  8'h75;        memory[34738] <=  8'h73;        memory[34739] <=  8'h6a;        memory[34740] <=  8'h63;        memory[34741] <=  8'h6e;        memory[34742] <=  8'h62;        memory[34743] <=  8'h64;        memory[34744] <=  8'h66;        memory[34745] <=  8'h73;        memory[34746] <=  8'h74;        memory[34747] <=  8'h79;        memory[34748] <=  8'h75;        memory[34749] <=  8'h61;        memory[34750] <=  8'h69;        memory[34751] <=  8'h6b;        memory[34752] <=  8'h78;        memory[34753] <=  8'h6d;        memory[34754] <=  8'h6e;        memory[34755] <=  8'h73;        memory[34756] <=  8'h6a;        memory[34757] <=  8'h6f;        memory[34758] <=  8'h64;        memory[34759] <=  8'h6c;        memory[34760] <=  8'h63;        memory[34761] <=  8'h78;        memory[34762] <=  8'h2c;        memory[34763] <=  8'h6d;        memory[34764] <=  8'h73;        memory[34765] <=  8'h6b;        memory[34766] <=  8'h64;        memory[34767] <=  8'h6c;        memory[34768] <=  8'h70;        memory[34769] <=  8'h5b;        memory[34770] <=  8'h3b;        memory[34771] <=  8'h73;        memory[34772] <=  8'h6c;        memory[34773] <=  8'h64;        memory[34774] <=  8'h70;        memory[34775] <=  8'h76;        memory[34776] <=  8'h63;        memory[34777] <=  8'h5b;        memory[34778] <=  8'h78;        memory[34779] <=  8'h76;        memory[34780] <=  8'h63;        memory[34781] <=  8'h5b;        memory[34782] <=  8'h78;        memory[34783] <=  8'h70;        memory[34784] <=  8'h6f;        memory[34785] <=  8'h20;        memory[34786] <=  8'h62;        memory[34787] <=  8'h61;        memory[34788] <=  8'h72;        memory[34789] <=  8'h74;        memory[34790] <=  8'h74;        memory[34791] <=  8'h62;        memory[34792] <=  8'h61;        memory[34793] <=  8'h72;        memory[34794] <=  8'h74;        memory[34795] <=  8'h78;        memory[34796] <=  8'h61;        memory[34797] <=  8'h74;        memory[34798] <=  8'h6b;        memory[34799] <=  8'h73;        memory[34800] <=  8'h68;        memory[34801] <=  8'h63;        memory[34802] <=  8'h66;        memory[34803] <=  8'h69;        memory[34804] <=  8'h77;        memory[34805] <=  8'h68;        memory[34806] <=  8'h61;        memory[34807] <=  8'h69;        memory[34808] <=  8'h6a;        memory[34809] <=  8'h78;        memory[34810] <=  8'h5d;        memory[34811] <=  8'h65;        memory[34812] <=  8'h6b;        memory[34813] <=  8'h6f;        memory[34814] <=  8'h39;        memory[34815] <=  8'h64;        memory[34816] <=  8'h75;        memory[34817] <=  8'h38;        memory[34818] <=  8'h79;        memory[34819] <=  8'h20;        memory[34820] <=  8'h37;        memory[34821] <=  8'h63;        memory[34822] <=  8'h67;        memory[34823] <=  8'h78;        memory[34824] <=  8'h63;        memory[34825] <=  8'h75;        memory[34826] <=  8'h68;        memory[34827] <=  8'h69;        memory[34828] <=  8'h6a;        memory[34829] <=  8'h77;        memory[34830] <=  8'h69;        memory[34831] <=  8'h64;        memory[34832] <=  8'h66;        memory[34833] <=  8'h68;        memory[34834] <=  8'h75;        memory[34835] <=  8'h76;        memory[34836] <=  8'h64;        memory[34837] <=  8'h62;        memory[34838] <=  8'h66;        memory[34839] <=  8'h6a;        memory[34840] <=  8'h6e;        memory[34841] <=  8'h6b;        memory[34842] <=  8'h6a;        memory[34843] <=  8'h65;        memory[34844] <=  8'h38;        memory[34845] <=  8'h66;        memory[34846] <=  8'h37;        memory[34847] <=  8'h67;        memory[34848] <=  8'h79;        memory[34849] <=  8'h76;        memory[34850] <=  8'h63;        memory[34851] <=  8'h68;        memory[34852] <=  8'h69;        memory[34853] <=  8'h6a;        memory[34854] <=  8'h33;        memory[34855] <=  8'h65;        memory[34856] <=  8'h67;        memory[34857] <=  8'h79;        memory[34858] <=  8'h72;        memory[34859] <=  8'h64;        memory[34860] <=  8'h62;        memory[34861] <=  8'h6e;        memory[34862] <=  8'h63;        memory[34863] <=  8'h7a;        memory[34864] <=  8'h6a;        memory[34865] <=  8'h6f;        memory[34866] <=  8'h66;        memory[34867] <=  8'h78;        memory[34868] <=  8'h6a;        memory[34869] <=  8'h69;        memory[34870] <=  8'h63;        memory[34871] <=  8'h68;        memory[34872] <=  8'h62;        memory[34873] <=  8'h6e;        memory[34874] <=  8'h6d;        memory[34875] <=  8'h63;        memory[34876] <=  8'h73;        memory[34877] <=  8'h6c;        memory[34878] <=  8'h6b;        memory[34879] <=  8'h6a;        memory[34880] <=  8'h69;        memory[34881] <=  8'h68;        memory[34882] <=  8'h76;        memory[34883] <=  8'h75;        memory[34884] <=  8'h69;        memory[34885] <=  8'h64;        memory[34886] <=  8'h68;        memory[34887] <=  8'h75;        memory[34888] <=  8'h67;        memory[34889] <=  8'h79;        memory[34890] <=  8'h62;        memory[34891] <=  8'h68;        memory[34892] <=  8'h65;        memory[34893] <=  8'h6a;        memory[34894] <=  8'h72;        memory[34895] <=  8'h6b;        memory[34896] <=  8'h6a;        memory[34897] <=  8'h6f;        memory[34898] <=  8'h64;        memory[34899] <=  8'h67;        memory[34900] <=  8'h69;        memory[34901] <=  8'h75;        memory[34902] <=  8'h69;        memory[34903] <=  8'h67;        memory[34904] <=  8'h76;        memory[34905] <=  8'h79;        memory[34906] <=  8'h75;        memory[34907] <=  8'h67;        memory[34908] <=  8'h78;        memory[34909] <=  8'h68;        memory[34910] <=  8'h63;        memory[34911] <=  8'h20;        memory[34912] <=  8'h20;        memory[34913] <=  8'h20;        memory[34914] <=  8'h78;        memory[34915] <=  8'h76;        memory[34916] <=  8'h20;        memory[34917] <=  8'h63;        memory[34918] <=  8'h78;        memory[34919] <=  8'h67;        memory[34920] <=  8'h79;        memory[34921] <=  8'h63;        memory[34922] <=  8'h75;        memory[34923] <=  8'h68;        memory[34924] <=  8'h6a;        memory[34925] <=  8'h6b;        memory[34926] <=  8'h61;        memory[34927] <=  8'h6c;        memory[34928] <=  8'h78;        memory[34929] <=  8'h76;        memory[34930] <=  8'h70;        memory[34931] <=  8'h6f;        memory[34932] <=  8'h69;        memory[34933] <=  8'h6a;        memory[34934] <=  8'h69;        memory[34935] <=  8'h68;        memory[34936] <=  8'h6a;        memory[34937] <=  8'h62;        memory[34938] <=  8'h77;        memory[34939] <=  8'h65;        memory[34940] <=  8'h6e;        memory[34941] <=  8'h61;        memory[34942] <=  8'h66;        memory[34943] <=  8'h6d;        memory[34944] <=  8'h64;        memory[34945] <=  8'h6b;        memory[34946] <=  8'h6d;        memory[34947] <=  8'h76;        memory[34948] <=  8'h6c;        memory[34949] <=  8'h63;        memory[34950] <=  8'h6f;        memory[34951] <=  8'h64;        memory[34952] <=  8'h69;        memory[34953] <=  8'h75;        memory[34954] <=  8'h68;        memory[34955] <=  8'h73;        memory[34956] <=  8'h66;        memory[34957] <=  8'h65;        memory[34958] <=  8'h62;        memory[34959] <=  8'h6e;        memory[34960] <=  8'h64;        memory[34961] <=  8'h73;        memory[34962] <=  8'h63;        memory[34963] <=  8'h6b;        memory[34964] <=  8'h20;        memory[34965] <=  8'h78;        memory[34966] <=  8'h6a;        memory[34967] <=  8'h78;        memory[34968] <=  8'h63;        memory[34969] <=  8'h73;        memory[34970] <=  8'h64;        memory[34971] <=  8'h66;        memory[34972] <=  8'h6b;        memory[34973] <=  8'h64;        memory[34974] <=  8'h6e;        memory[34975] <=  8'h6d;        memory[34976] <=  8'h64;        memory[34977] <=  8'h73;        memory[34978] <=  8'h63;        memory[34979] <=  8'h6b;        memory[34980] <=  8'h78;        memory[34981] <=  8'h6c;        memory[34982] <=  8'h6f;        memory[34983] <=  8'h66;        memory[34984] <=  8'h6a;        memory[34985] <=  8'h69;        memory[34986] <=  8'h61;        memory[34987] <=  8'h62;        memory[34988] <=  8'h6e;        memory[34989] <=  8'h20;        memory[34990] <=  8'h78;        memory[34991] <=  8'h6b;        memory[34992] <=  8'h6d;        memory[34993] <=  8'h20;        memory[34994] <=  8'h6f;        memory[34995] <=  8'h63;        memory[34996] <=  8'h76;        memory[34997] <=  8'h73;        memory[34998] <=  8'h64;        memory[34999] <=  8'h69;        memory[35000] <=  8'h66;        memory[35001] <=  8'h68;        memory[35002] <=  8'h65;        memory[35003] <=  8'h71;        memory[35004] <=  8'h6a;        memory[35005] <=  8'h77;        memory[35006] <=  8'h62;        memory[35007] <=  8'h65;        memory[35008] <=  8'h6e;        memory[35009] <=  8'h20;        memory[35010] <=  8'h6d;        memory[35011] <=  8'h64;        memory[35012] <=  8'h73;        memory[35013] <=  8'h6c;        memory[35014] <=  8'h76;        memory[35015] <=  8'h6b;        memory[35016] <=  8'h63;        memory[35017] <=  8'h78;        memory[35018] <=  8'h20;        memory[35019] <=  8'h6f;        memory[35020] <=  8'h78;        memory[35021] <=  8'h69;        memory[35022] <=  8'h63;        memory[35023] <=  8'h6a;        memory[35024] <=  8'h76;        memory[35025] <=  8'h64;        memory[35026] <=  8'h66;        memory[35027] <=  8'h65;        memory[35028] <=  8'h71;        memory[35029] <=  8'h6e;        memory[35030] <=  8'h20;        memory[35031] <=  8'h64;        memory[35032] <=  8'h6d;        memory[35033] <=  8'h73;        memory[35034] <=  8'h6c;        memory[35035] <=  8'h63;        memory[35036] <=  8'h78;        memory[35037] <=  8'h6b;        memory[35038] <=  8'h20;        memory[35039] <=  8'h6f;        memory[35040] <=  8'h78;        memory[35041] <=  8'h63;        memory[35042] <=  8'h76;        memory[35043] <=  8'h6a;        memory[35044] <=  8'h64;        memory[35045] <=  8'h62;        memory[35046] <=  8'h71;        memory[35047] <=  8'h77;        memory[35048] <=  8'h65;        memory[35049] <=  8'h6e;        memory[35050] <=  8'h6d;        memory[35051] <=  8'h64;        memory[35052] <=  8'h6c;        memory[35053] <=  8'h73;        memory[35054] <=  8'h2c;        memory[35055] <=  8'h76;        memory[35056] <=  8'h63;        memory[35057] <=  8'h78;        memory[35058] <=  8'h20;        memory[35059] <=  8'h63;        memory[35060] <=  8'h6f;        memory[35061] <=  8'h69;        memory[35062] <=  8'h76;        memory[35063] <=  8'h68;        memory[35064] <=  8'h73;        memory[35065] <=  8'h64;        memory[35066] <=  8'h62;        memory[35067] <=  8'h71;        memory[35068] <=  8'h77;        memory[35069] <=  8'h65;        memory[35070] <=  8'h6e;        memory[35071] <=  8'h64;        memory[35072] <=  8'h6b;        memory[35073] <=  8'h73;        memory[35074] <=  8'h76;        memory[35075] <=  8'h6f;        memory[35076] <=  8'h63;        memory[35077] <=  8'h20;        memory[35078] <=  8'h76;        memory[35079] <=  8'h69;        memory[35080] <=  8'h75;        memory[35081] <=  8'h69;        memory[35082] <=  8'h68;        memory[35083] <=  8'h63;        memory[35084] <=  8'h78;        memory[35085] <=  8'h69;        memory[35086] <=  8'h6f;        memory[35087] <=  8'h76;        memory[35088] <=  8'h73;        memory[35089] <=  8'h64;        memory[35090] <=  8'h61;        memory[35091] <=  8'h64;        memory[35092] <=  8'h6e;        memory[35093] <=  8'h77;        memory[35094] <=  8'h71;        memory[35095] <=  8'h6b;        memory[35096] <=  8'h6c;        memory[35097] <=  8'h73;        memory[35098] <=  8'h76;        memory[35099] <=  8'h6e;        memory[35100] <=  8'h62;        memory[35101] <=  8'h20;        memory[35102] <=  8'h64;        memory[35103] <=  8'h66;        memory[35104] <=  8'h6a;        memory[35105] <=  8'h6b;        memory[35106] <=  8'h71;        memory[35107] <=  8'h64;        memory[35108] <=  8'h77;        memory[35109] <=  8'h65;        memory[35110] <=  8'h6e;        memory[35111] <=  8'h62;        memory[35112] <=  8'h20;        memory[35113] <=  8'h64;        memory[35114] <=  8'h73;        memory[35115] <=  8'h76;        memory[35116] <=  8'h68;        memory[35117] <=  8'h64;        memory[35118] <=  8'h61;        memory[35119] <=  8'h71;        memory[35120] <=  8'h77;        memory[35121] <=  8'h6a;        memory[35122] <=  8'h65;        memory[35123] <=  8'h6e;        memory[35124] <=  8'h64;        memory[35125] <=  8'h20;        memory[35126] <=  8'h61;        memory[35127] <=  8'h63;        memory[35128] <=  8'h62;        memory[35129] <=  8'h68;        memory[35130] <=  8'h64;        memory[35131] <=  8'h61;        memory[35132] <=  8'h77;        memory[35133] <=  8'h71;        memory[35134] <=  8'h6e;        memory[35135] <=  8'h20;        memory[35136] <=  8'h62;        memory[35137] <=  8'h73;        memory[35138] <=  8'h76;        memory[35139] <=  8'h61;        memory[35140] <=  8'h67;        memory[35141] <=  8'h76;        memory[35142] <=  8'h68;        memory[35143] <=  8'h67;        memory[35144] <=  8'h61;        memory[35145] <=  8'h73;        memory[35146] <=  8'h6a;        memory[35147] <=  8'h6b;        memory[35148] <=  8'h63;        memory[35149] <=  8'h78;        memory[35150] <=  8'h76;        memory[35151] <=  8'h6e;        memory[35152] <=  8'h73;        memory[35153] <=  8'h64;        memory[35154] <=  8'h20;        memory[35155] <=  8'h66;        memory[35156] <=  8'h62;        memory[35157] <=  8'h64;        memory[35158] <=  8'h61;        memory[35159] <=  8'h73;        memory[35160] <=  8'h76;        memory[35161] <=  8'h67;        memory[35162] <=  8'h63;        memory[35163] <=  8'h79;        memory[35164] <=  8'h7a;        memory[35165] <=  8'h78;        memory[35166] <=  8'h79;        memory[35167] <=  8'h75;        memory[35168] <=  8'h20;        memory[35169] <=  8'h69;        memory[35170] <=  8'h6a;        memory[35171] <=  8'h64;        memory[35172] <=  8'h66;        memory[35173] <=  8'h6b;        memory[35174] <=  8'h61;        memory[35175] <=  8'h64;        memory[35176] <=  8'h63;        memory[35177] <=  8'h78;        memory[35178] <=  8'h68;        memory[35179] <=  8'h20;        memory[35180] <=  8'h67;        memory[35181] <=  8'h61;        memory[35182] <=  8'h68;        memory[35183] <=  8'h75;        memory[35184] <=  8'h64;        memory[35185] <=  8'h73;        memory[35186] <=  8'h69;        memory[35187] <=  8'h6a;        memory[35188] <=  8'h61;        memory[35189] <=  8'h6b;        memory[35190] <=  8'h63;        memory[35191] <=  8'h62;        memory[35192] <=  8'h61;        memory[35193] <=  8'h72;        memory[35194] <=  8'h73;        memory[35195] <=  8'h68;        memory[35196] <=  8'h64;        memory[35197] <=  8'h66;        memory[35198] <=  8'h67;        memory[35199] <=  8'h73;        memory[35200] <=  8'h68;        memory[35201] <=  8'h64;        memory[35202] <=  8'h66;        memory[35203] <=  8'h68;        memory[35204] <=  8'h64;        memory[35205] <=  8'h6a;        memory[35206] <=  8'h68;        memory[35207] <=  8'h62;        memory[35208] <=  8'h67;        memory[35209] <=  8'h63;        memory[35210] <=  8'h61;        memory[35211] <=  8'h66;        memory[35212] <=  8'h73;        memory[35213] <=  8'h79;        memory[35214] <=  8'h67;        memory[35215] <=  8'h6b;        memory[35216] <=  8'h75;        memory[35217] <=  8'h64;        memory[35218] <=  8'h68;        memory[35219] <=  8'h62;        memory[35220] <=  8'h77;        memory[35221] <=  8'h76;        memory[35222] <=  8'h67;        memory[35223] <=  8'h61;        memory[35224] <=  8'h66;        memory[35225] <=  8'h64;        memory[35226] <=  8'h74;        memory[35227] <=  8'h75;        memory[35228] <=  8'h66;        memory[35229] <=  8'h79;        memory[35230] <=  8'h67;        memory[35231] <=  8'h69;        memory[35232] <=  8'h75;        memory[35233] <=  8'h68;        memory[35234] <=  8'h6c;        memory[35235] <=  8'h6a;        memory[35236] <=  8'h62;        memory[35237] <=  8'h6b;        memory[35238] <=  8'h68;        memory[35239] <=  8'h76;        memory[35240] <=  8'h67;        memory[35241] <=  8'h63;        memory[35242] <=  8'h66;        memory[35243] <=  8'h78;        memory[35244] <=  8'h64;        memory[35245] <=  8'h74;        memory[35246] <=  8'h75;        memory[35247] <=  8'h79;        memory[35248] <=  8'h69;        memory[35249] <=  8'h75;        memory[35250] <=  8'h68;        memory[35251] <=  8'h6c;        memory[35252] <=  8'h6a;        memory[35253] <=  8'h6b;        memory[35254] <=  8'h67;        memory[35255] <=  8'h6a;        memory[35256] <=  8'h63;        memory[35257] <=  8'h66;        memory[35258] <=  8'h68;        memory[35259] <=  8'h64;        memory[35260] <=  8'h67;        memory[35261] <=  8'h72;        memory[35262] <=  8'h79;        memory[35263] <=  8'h74;        memory[35264] <=  8'h66;        memory[35265] <=  8'h75;        memory[35266] <=  8'h79;        memory[35267] <=  8'h69;        memory[35268] <=  8'h68;        memory[35269] <=  8'h6c;        memory[35270] <=  8'h62;        memory[35271] <=  8'h6d;        memory[35272] <=  8'h76;        memory[35273] <=  8'h6e;        memory[35274] <=  8'h63;        memory[35275] <=  8'h66;        memory[35276] <=  8'h68;        memory[35277] <=  8'h64;        memory[35278] <=  8'h74;        memory[35279] <=  8'h75;        memory[35280] <=  8'h67;        memory[35281] <=  8'h79;        memory[35282] <=  8'h69;        memory[35283] <=  8'h68;        memory[35284] <=  8'h75;        memory[35285] <=  8'h6a;        memory[35286] <=  8'h6c;        memory[35287] <=  8'h62;        memory[35288] <=  8'h6d;        memory[35289] <=  8'h76;        memory[35290] <=  8'h6e;        memory[35291] <=  8'h63;        memory[35292] <=  8'h66;        memory[35293] <=  8'h68;        memory[35294] <=  8'h67;        memory[35295] <=  8'h79;        memory[35296] <=  8'h68;        memory[35297] <=  8'h75;        memory[35298] <=  8'h6a;        memory[35299] <=  8'h6e;        memory[35300] <=  8'h2c;        memory[35301] <=  8'h62;        memory[35302] <=  8'h6e;        memory[35303] <=  8'h6d;        memory[35304] <=  8'h76;        memory[35305] <=  8'h6e;        memory[35306] <=  8'h63;        memory[35307] <=  8'h66;        memory[35308] <=  8'h68;        memory[35309] <=  8'h74;        memory[35310] <=  8'h79;        memory[35311] <=  8'h69;        memory[35312] <=  8'h75;        memory[35313] <=  8'h6c;        memory[35314] <=  8'h6a;        memory[35315] <=  8'h62;        memory[35316] <=  8'h6d;        memory[35317] <=  8'h76;        memory[35318] <=  8'h6e;        memory[35319] <=  8'h63;        memory[35320] <=  8'h66;        memory[35321] <=  8'h74;        memory[35322] <=  8'h75;        memory[35323] <=  8'h79;        memory[35324] <=  8'h69;        memory[35325] <=  8'h68;        memory[35326] <=  8'h6b;        memory[35327] <=  8'h62;        memory[35328] <=  8'h76;        memory[35329] <=  8'h63;        memory[35330] <=  8'h66;        memory[35331] <=  8'h67;        memory[35332] <=  8'h74;        memory[35333] <=  8'h75;        memory[35334] <=  8'h79;        memory[35335] <=  8'h69;        memory[35336] <=  8'h75;        memory[35337] <=  8'h68;        memory[35338] <=  8'h6a;        memory[35339] <=  8'h6b;        memory[35340] <=  8'h62;        memory[35341] <=  8'h76;        memory[35342] <=  8'h63;        memory[35343] <=  8'h66;        memory[35344] <=  8'h74;        memory[35345] <=  8'h75;        memory[35346] <=  8'h79;        memory[35347] <=  8'h69;        memory[35348] <=  8'h75;        memory[35349] <=  8'h6a;        memory[35350] <=  8'h6b;        memory[35351] <=  8'h6e;        memory[35352] <=  8'h62;        memory[35353] <=  8'h76;        memory[35354] <=  8'h67;        memory[35355] <=  8'h66;        memory[35356] <=  8'h74;        memory[35357] <=  8'h79;        memory[35358] <=  8'h75;        memory[35359] <=  8'h75;        memory[35360] <=  8'h69;        memory[35361] <=  8'h6a;        memory[35362] <=  8'h6b;        memory[35363] <=  8'h68;        memory[35364] <=  8'h62;        memory[35365] <=  8'h6a;        memory[35366] <=  8'h67;        memory[35367] <=  8'h68;        memory[35368] <=  8'h66;        memory[35369] <=  8'h79;        memory[35370] <=  8'h74;        memory[35371] <=  8'h79;        memory[35372] <=  8'h69;        memory[35373] <=  8'h75;        memory[35374] <=  8'h64;        memory[35375] <=  8'h6a;        memory[35376] <=  8'h6b;        memory[35377] <=  8'h68;        memory[35378] <=  8'h63;        memory[35379] <=  8'h7a;        memory[35380] <=  8'h67;        memory[35381] <=  8'h68;        memory[35382] <=  8'h74;        memory[35383] <=  8'h75;        memory[35384] <=  8'h79;        memory[35385] <=  8'h69;        memory[35386] <=  8'h61;        memory[35387] <=  8'h73;        memory[35388] <=  8'h75;        memory[35389] <=  8'h6a;        memory[35390] <=  8'h6b;        memory[35391] <=  8'h62;        memory[35392] <=  8'h6e;        memory[35393] <=  8'h61;        memory[35394] <=  8'h76;        memory[35395] <=  8'h63;        memory[35396] <=  8'h66;        memory[35397] <=  8'h68;        memory[35398] <=  8'h75;        memory[35399] <=  8'h61;        memory[35400] <=  8'h73;        memory[35401] <=  8'h79;        memory[35402] <=  8'h64;        memory[35403] <=  8'h75;        memory[35404] <=  8'h69;        memory[35405] <=  8'h6a;        memory[35406] <=  8'h61;        memory[35407] <=  8'h6b;        memory[35408] <=  8'h62;        memory[35409] <=  8'h63;        memory[35410] <=  8'h78;        memory[35411] <=  8'h68;        memory[35412] <=  8'h67;        memory[35413] <=  8'h79;        memory[35414] <=  8'h75;        memory[35415] <=  8'h7a;        memory[35416] <=  8'h63;        memory[35417] <=  8'h61;        memory[35418] <=  8'h73;        memory[35419] <=  8'h69;        memory[35420] <=  8'h75;        memory[35421] <=  8'h6f;        memory[35422] <=  8'h69;        memory[35423] <=  8'h6a;        memory[35424] <=  8'h61;        memory[35425] <=  8'h6c;        memory[35426] <=  8'h63;        memory[35427] <=  8'h78;        memory[35428] <=  8'h62;        memory[35429] <=  8'h63;        memory[35430] <=  8'h20;        memory[35431] <=  8'h6e;        memory[35432] <=  8'h76;        memory[35433] <=  8'h63;        memory[35434] <=  8'h61;        memory[35435] <=  8'h64;        memory[35436] <=  8'h73;        memory[35437] <=  8'h67;        memory[35438] <=  8'h79;        memory[35439] <=  8'h68;        memory[35440] <=  8'h75;        memory[35441] <=  8'h61;        memory[35442] <=  8'h6a;        memory[35443] <=  8'h6b;        memory[35444] <=  8'h78;        memory[35445] <=  8'h62;        memory[35446] <=  8'h20;        memory[35447] <=  8'h6e;        memory[35448] <=  8'h76;        memory[35449] <=  8'h63;        memory[35450] <=  8'h61;        memory[35451] <=  8'h73;        memory[35452] <=  8'h67;        memory[35453] <=  8'h68;        memory[35454] <=  8'h75;        memory[35455] <=  8'h6a;        memory[35456] <=  8'h6c;        memory[35457] <=  8'h6b;        memory[35458] <=  8'h63;        memory[35459] <=  8'h78;        memory[35460] <=  8'h20;        memory[35461] <=  8'h6a;        memory[35462] <=  8'h6b;        memory[35463] <=  8'h68;        memory[35464] <=  8'h61;        memory[35465] <=  8'h73;        memory[35466] <=  8'h76;        memory[35467] <=  8'h64;        memory[35468] <=  8'h6e;        memory[35469] <=  8'h20;        memory[35470] <=  8'h62;        memory[35471] <=  8'h6e;        memory[35472] <=  8'h6d;        memory[35473] <=  8'h6b;        memory[35474] <=  8'h77;        memory[35475] <=  8'h64;        memory[35476] <=  8'h6f;        memory[35477] <=  8'h77;        memory[35478] <=  8'h69;        memory[35479] <=  8'h6f;        memory[35480] <=  8'h75;        memory[35481] <=  8'h69;        memory[35482] <=  8'h68;        memory[35483] <=  8'h62;        memory[35484] <=  8'h6e;        memory[35485] <=  8'h6b;        memory[35486] <=  8'h77;        memory[35487] <=  8'h69;        memory[35488] <=  8'h6f;        memory[35489] <=  8'h75;        memory[35490] <=  8'h71;        memory[35491] <=  8'h69;        memory[35492] <=  8'h79;        memory[35493] <=  8'h67;        memory[35494] <=  8'h6a;        memory[35495] <=  8'h64;        memory[35496] <=  8'h61;        memory[35497] <=  8'h76;        memory[35498] <=  8'h62;        memory[35499] <=  8'h6e;        memory[35500] <=  8'h6b;        memory[35501] <=  8'h6f;        memory[35502] <=  8'h70;        memory[35503] <=  8'h64;        memory[35504] <=  8'h76;        memory[35505] <=  8'h69;        memory[35506] <=  8'h6f;        memory[35507] <=  8'h75;        memory[35508] <=  8'h69;        memory[35509] <=  8'h48;        memory[35510] <=  8'h42;        memory[35511] <=  8'h6b;        memory[35512] <=  8'h64;        memory[35513] <=  8'h6e;        memory[35514] <=  8'h6c;        memory[35515] <=  8'h71;        memory[35516] <=  8'h6b;        memory[35517] <=  8'h6d;        memory[35518] <=  8'h6a;        memory[35519] <=  8'h70;        memory[35520] <=  8'h69;        memory[35521] <=  8'h6f;        memory[35522] <=  8'h68;        memory[35523] <=  8'h65;        memory[35524] <=  8'h66;        memory[35525] <=  8'h75;        memory[35526] <=  8'h67;        memory[35527] <=  8'h69;        memory[35528] <=  8'h73;        memory[35529] <=  8'h61;        memory[35530] <=  8'h62;        memory[35531] <=  8'h64;        memory[35532] <=  8'h6b;        memory[35533] <=  8'h6a;        memory[35534] <=  8'h6b;        memory[35535] <=  8'h6c;        memory[35536] <=  8'h6a;        memory[35537] <=  8'h69;        memory[35538] <=  8'h73;        memory[35539] <=  8'h6f;        memory[35540] <=  8'h71;        memory[35541] <=  8'h68;        memory[35542] <=  8'h77;        memory[35543] <=  8'h67;        memory[35544] <=  8'h69;        memory[35545] <=  8'h79;        memory[35546] <=  8'h6a;        memory[35547] <=  8'h64;        memory[35548] <=  8'h76;        memory[35549] <=  8'h62;        memory[35550] <=  8'h6e;        memory[35551] <=  8'h61;        memory[35552] <=  8'h73;        memory[35553] <=  8'h66;        memory[35554] <=  8'h6c;        memory[35555] <=  8'h6b;        memory[35556] <=  8'h64;        memory[35557] <=  8'h6a;        memory[35558] <=  8'h68;        memory[35559] <=  8'h63;        memory[35560] <=  8'h67;        memory[35561] <=  8'h6a;        memory[35562] <=  8'h76;        memory[35563] <=  8'h73;        memory[35564] <=  8'h64;        memory[35565] <=  8'h62;        memory[35566] <=  8'h62;        memory[35567] <=  8'h61;        memory[35568] <=  8'h72;        memory[35569] <=  8'h62;        memory[35570] <=  8'h62;        memory[35571] <=  8'h73;        memory[35572] <=  8'h62;        memory[35573] <=  8'h67;        memory[35574] <=  8'h73;        memory[35575] <=  8'h66;        memory[35576] <=  8'h67;        memory[35577] <=  8'h61;        memory[35578] <=  8'h68;        memory[35579] <=  8'h66;        memory[35580] <=  8'h73;        memory[35581] <=  8'h68;        memory[35582] <=  8'h61;        memory[35583] <=  8'h66;        memory[35584] <=  8'h73;        memory[35585] <=  8'h66;        memory[35586] <=  8'h68;        memory[35587] <=  8'h61;        memory[35588] <=  8'h69;        memory[35589] <=  8'h64;        memory[35590] <=  8'h75;        memory[35591] <=  8'h67;        memory[35592] <=  8'h64;        memory[35593] <=  8'h77;        memory[35594] <=  8'h62;        memory[35595] <=  8'h61;        memory[35596] <=  8'h62;        memory[35597] <=  8'h72;        memory[35598] <=  8'h62;        memory[35599] <=  8'h61;        memory[35600] <=  8'h62;        memory[35601] <=  8'h62;        memory[35602] <=  8'h74;        memory[35603] <=  8'h62;        memory[35604] <=  8'h62;        memory[35605] <=  8'h62;        memory[35606] <=  8'h62;        memory[35607] <=  8'h62;        memory[35608] <=  8'h62;        memory[35609] <=  8'h62;        memory[35610] <=  8'h62;        memory[35611] <=  8'h61;        memory[35612] <=  8'h62;        memory[35613] <=  8'h62;        memory[35614] <=  8'h72;        memory[35615] <=  8'h74;        memory[35616] <=  8'h62;        memory[35617] <=  8'h62;        memory[35618] <=  8'h61;        memory[35619] <=  8'h62;        memory[35620] <=  8'h72;        memory[35621] <=  8'h62;        memory[35622] <=  8'h74;        memory[35623] <=  8'h62;        memory[35624] <=  8'h62;        memory[35625] <=  8'h62;        memory[35626] <=  8'h63;        memory[35627] <=  8'h61;        memory[35628] <=  8'h72;        memory[35629] <=  8'h74;        memory[35630] <=  8'h73;        memory[35631] <=  8'h62;        memory[35632] <=  8'h61;        memory[35633] <=  8'h72;        memory[35634] <=  8'h74;        memory[35635] <=  8'h74;        memory[35636] <=  8'h62;        memory[35637] <=  8'h61;        memory[35638] <=  8'h72;        memory[35639] <=  8'h74;        memory[35640] <=  8'h78;        memory[35641] <=  8'h61;        memory[35642] <=  8'h74;        memory[35643] <=  8'h6b;        memory[35644] <=  8'h73;        memory[35645] <=  8'h68;        memory[35646] <=  8'h63;        memory[35647] <=  8'h66;        memory[35648] <=  8'h69;        memory[35649] <=  8'h77;        memory[35650] <=  8'h68;        memory[35651] <=  8'h61;        memory[35652] <=  8'h74;        memory[35653] <=  8'h61;        memory[35654] <=  8'h6e;        memory[35655] <=  8'h61;        memory[35656] <=  8'h62;        memory[35657] <=  8'h61;        memory[35658] <=  8'h63;        memory[35659] <=  8'h61;        memory[35660] <=  8'h74;        memory[35661] <=  8'h61;        memory[35662] <=  8'h62;        memory[35663] <=  8'h61;        memory[35664] <=  8'h72;        memory[35665] <=  8'h63;        memory[35666] <=  8'h61;        memory[35667] <=  8'h68;        memory[35668] <=  8'h64;        memory[35669] <=  8'h75;        memory[35670] <=  8'h63;        memory[35671] <=  8'h74;        memory[35672] <=  8'h61;        memory[35673] <=  8'h64;        memory[35674] <=  8'h61;        memory[35675] <=  8'h61;        memory[35676] <=  8'h63;        memory[35677] <=  8'h61;        memory[35678] <=  8'h72;        memory[35679] <=  8'h63;        memory[35680] <=  8'h74;        memory[35681] <=  8'h72;        memory[35682] <=  8'h63;        memory[35683] <=  8'h61;        memory[35684] <=  8'h74;        memory[35685] <=  8'h72;        memory[35686] <=  8'h63;        memory[35687] <=  8'h61;        memory[35688] <=  8'h74;        memory[35689] <=  8'h63;        memory[35690] <=  8'h62;        memory[35691] <=  8'h61;        memory[35692] <=  8'h74;        memory[35693] <=  8'h62;        memory[35694] <=  8'h72;        memory[35695] <=  8'h63;        memory[35696] <=  8'h61;        memory[35697] <=  8'h74;        memory[35698] <=  8'h72;        memory[35699] <=  8'h6e;        memory[35700] <=  8'h62;        memory[35701] <=  8'h61;        memory[35702] <=  8'h63;        memory[35703] <=  8'h61;        memory[35704] <=  8'h74;        memory[35705] <=  8'h79;        memory[35706] <=  8'h73;        memory[35707] <=  8'h6e;        memory[35708] <=  8'h63;        memory[35709] <=  8'h74;        memory[35710] <=  8'h61;        memory[35711] <=  8'h6e;        memory[35712] <=  8'h62;        memory[35713] <=  8'h61;        memory[35714] <=  8'h63;        memory[35715] <=  8'h72;        memory[35716] <=  8'h6e;        memory[35717] <=  8'h74;        memory[35718] <=  8'h61;        memory[35719] <=  8'h62;        memory[35720] <=  8'h74;        memory[35721] <=  8'h6e;        memory[35722] <=  8'h61;        memory[35723] <=  8'h72;        memory[35724] <=  8'h62;        memory[35725] <=  8'h78;        memory[35726] <=  8'h74;        memory[35727] <=  8'h61;        memory[35728] <=  8'h72;        memory[35729] <=  8'h62;        memory[35730] <=  8'h61;        memory[35731] <=  8'h72;        memory[35732] <=  8'h74;        memory[35733] <=  8'h74;        memory[35734] <=  8'h62;        memory[35735] <=  8'h61;        memory[35736] <=  8'h72;        memory[35737] <=  8'h74;        memory[35738] <=  8'h78;        memory[35739] <=  8'h61;        memory[35740] <=  8'h74;        memory[35741] <=  8'h6b;        memory[35742] <=  8'h73;        memory[35743] <=  8'h68;        memory[35744] <=  8'h63;        memory[35745] <=  8'h66;        memory[35746] <=  8'h69;        memory[35747] <=  8'h77;        memory[35748] <=  8'h68;        memory[35749] <=  8'h61;        memory[35750] <=  8'h74;        memory[35751] <=  8'h61;        memory[35752] <=  8'h6e;        memory[35753] <=  8'h61;        memory[35754] <=  8'h62;        memory[35755] <=  8'h61;        memory[35756] <=  8'h63;        memory[35757] <=  8'h61;        memory[35758] <=  8'h74;        memory[35759] <=  8'h61;        memory[35760] <=  8'h62;        memory[35761] <=  8'h61;        memory[35762] <=  8'h72;        memory[35763] <=  8'h63;        memory[35764] <=  8'h61;        memory[35765] <=  8'h68;        memory[35766] <=  8'h64;        memory[35767] <=  8'h75;        memory[35768] <=  8'h63;        memory[35769] <=  8'h74;        memory[35770] <=  8'h61;        memory[35771] <=  8'h64;        memory[35772] <=  8'h61;        memory[35773] <=  8'h61;        memory[35774] <=  8'h63;        memory[35775] <=  8'h61;        memory[35776] <=  8'h72;        memory[35777] <=  8'h63;        memory[35778] <=  8'h74;        memory[35779] <=  8'h72;        memory[35780] <=  8'h63;        memory[35781] <=  8'h61;        memory[35782] <=  8'h74;        memory[35783] <=  8'h72;        memory[35784] <=  8'h63;        memory[35785] <=  8'h61;        memory[35786] <=  8'h74;        memory[35787] <=  8'h63;        memory[35788] <=  8'h62;        memory[35789] <=  8'h61;        memory[35790] <=  8'h74;        memory[35791] <=  8'h62;        memory[35792] <=  8'h72;        memory[35793] <=  8'h63;        memory[35794] <=  8'h61;        memory[35795] <=  8'h74;        memory[35796] <=  8'h72;        memory[35797] <=  8'h6e;        memory[35798] <=  8'h62;        memory[35799] <=  8'h61;        memory[35800] <=  8'h63;        memory[35801] <=  8'h61;        memory[35802] <=  8'h74;        memory[35803] <=  8'h79;        memory[35804] <=  8'h73;        memory[35805] <=  8'h6e;        memory[35806] <=  8'h63;        memory[35807] <=  8'h74;        memory[35808] <=  8'h61;        memory[35809] <=  8'h6e;        memory[35810] <=  8'h62;        memory[35811] <=  8'h61;        memory[35812] <=  8'h63;        memory[35813] <=  8'h72;        memory[35814] <=  8'h6e;        memory[35815] <=  8'h74;        memory[35816] <=  8'h61;        memory[35817] <=  8'h62;        memory[35818] <=  8'h74;        memory[35819] <=  8'h6e;        memory[35820] <=  8'h61;        memory[35821] <=  8'h72;        memory[35822] <=  8'h62;        memory[35823] <=  8'h78;        memory[35824] <=  8'h74;        memory[35825] <=  8'h61;        memory[35826] <=  8'h72;        memory[35827] <=  8'h62;        memory[35828] <=  8'h61;        memory[35829] <=  8'h72;        memory[35830] <=  8'h74;        memory[35831] <=  8'h74;        memory[35832] <=  8'h62;        memory[35833] <=  8'h61;        memory[35834] <=  8'h72;        memory[35835] <=  8'h74;        memory[35836] <=  8'h78;        memory[35837] <=  8'h61;        memory[35838] <=  8'h74;        memory[35839] <=  8'h6b;        memory[35840] <=  8'h73;        memory[35841] <=  8'h68;        memory[35842] <=  8'h63;        memory[35843] <=  8'h66;        memory[35844] <=  8'h69;        memory[35845] <=  8'h77;        memory[35846] <=  8'h68;        memory[35847] <=  8'h61;        memory[35848] <=  8'h74;        memory[35849] <=  8'h61;        memory[35850] <=  8'h6e;        memory[35851] <=  8'h61;        memory[35852] <=  8'h62;        memory[35853] <=  8'h61;        memory[35854] <=  8'h63;        memory[35855] <=  8'h61;        memory[35856] <=  8'h74;        memory[35857] <=  8'h61;        memory[35858] <=  8'h62;        memory[35859] <=  8'h61;        memory[35860] <=  8'h72;        memory[35861] <=  8'h63;        memory[35862] <=  8'h61;        memory[35863] <=  8'h68;        memory[35864] <=  8'h64;        memory[35865] <=  8'h75;        memory[35866] <=  8'h63;        memory[35867] <=  8'h74;        memory[35868] <=  8'h61;        memory[35869] <=  8'h64;        memory[35870] <=  8'h61;        memory[35871] <=  8'h61;        memory[35872] <=  8'h63;        memory[35873] <=  8'h61;        memory[35874] <=  8'h72;        memory[35875] <=  8'h63;        memory[35876] <=  8'h74;        memory[35877] <=  8'h72;        memory[35878] <=  8'h63;        memory[35879] <=  8'h61;        memory[35880] <=  8'h74;        memory[35881] <=  8'h72;        memory[35882] <=  8'h63;        memory[35883] <=  8'h61;        memory[35884] <=  8'h74;        memory[35885] <=  8'h63;        memory[35886] <=  8'h62;        memory[35887] <=  8'h61;        memory[35888] <=  8'h74;        memory[35889] <=  8'h62;        memory[35890] <=  8'h72;        memory[35891] <=  8'h63;        memory[35892] <=  8'h61;        memory[35893] <=  8'h74;        memory[35894] <=  8'h72;        memory[35895] <=  8'h6e;        memory[35896] <=  8'h62;        memory[35897] <=  8'h61;        memory[35898] <=  8'h63;        memory[35899] <=  8'h61;        memory[35900] <=  8'h74;        memory[35901] <=  8'h79;        memory[35902] <=  8'h73;        memory[35903] <=  8'h6e;        memory[35904] <=  8'h63;        memory[35905] <=  8'h74;        memory[35906] <=  8'h61;        memory[35907] <=  8'h6e;        memory[35908] <=  8'h62;        memory[35909] <=  8'h61;        memory[35910] <=  8'h63;        memory[35911] <=  8'h72;        memory[35912] <=  8'h6e;        memory[35913] <=  8'h74;        memory[35914] <=  8'h61;        memory[35915] <=  8'h62;        memory[35916] <=  8'h74;        memory[35917] <=  8'h6e;        memory[35918] <=  8'h61;        memory[35919] <=  8'h72;        memory[35920] <=  8'h62;        memory[35921] <=  8'h78;        memory[35922] <=  8'h74;        memory[35923] <=  8'h61;        memory[35924] <=  8'h72;        memory[35925] <=  8'h5d;        memory[35926] <=  8'h5d;        memory[35927] <=  8'h65;        memory[35928] <=  8'h66;        memory[35929] <=  8'h77;        memory[35930] <=  8'h65;        memory[35931] <=  8'h5d;        memory[35932] <=  8'h65;        memory[35933] <=  8'h67;        memory[35934] <=  8'h73;        memory[35935] <=  8'h67;        memory[35936] <=  8'h66;        memory[35937] <=  8'h62;        memory[35938] <=  8'h61;        memory[35939] <=  8'h72;        memory[35940] <=  8'h74;        memory[35941] <=  8'h74;        memory[35942] <=  8'h62;        memory[35943] <=  8'h61;        memory[35944] <=  8'h72;        memory[35945] <=  8'h74;        memory[35946] <=  8'h78;        memory[35947] <=  8'h61;        memory[35948] <=  8'h74;        memory[35949] <=  8'h6b;        memory[35950] <=  8'h73;        memory[35951] <=  8'h68;        memory[35952] <=  8'h63;        memory[35953] <=  8'h66;        memory[35954] <=  8'h69;        memory[35955] <=  8'h77;        memory[35956] <=  8'h68;        memory[35957] <=  8'h61;        memory[35958] <=  8'h74;        memory[35959] <=  8'h61;        memory[35960] <=  8'h6e;        memory[35961] <=  8'h61;        memory[35962] <=  8'h62;        memory[35963] <=  8'h61;        memory[35964] <=  8'h63;        memory[35965] <=  8'h61;        memory[35966] <=  8'h74;        memory[35967] <=  8'h61;        memory[35968] <=  8'h62;        memory[35969] <=  8'h61;        memory[35970] <=  8'h72;        memory[35971] <=  8'h63;        memory[35972] <=  8'h61;        memory[35973] <=  8'h68;        memory[35974] <=  8'h64;        memory[35975] <=  8'h75;        memory[35976] <=  8'h63;        memory[35977] <=  8'h74;        memory[35978] <=  8'h61;        memory[35979] <=  8'h64;        memory[35980] <=  8'h61;        memory[35981] <=  8'h61;        memory[35982] <=  8'h63;        memory[35983] <=  8'h61;        memory[35984] <=  8'h72;        memory[35985] <=  8'h63;        memory[35986] <=  8'h74;        memory[35987] <=  8'h72;        memory[35988] <=  8'h63;        memory[35989] <=  8'h61;        memory[35990] <=  8'h74;        memory[35991] <=  8'h72;        memory[35992] <=  8'h63;        memory[35993] <=  8'h61;        memory[35994] <=  8'h74;        memory[35995] <=  8'h63;        memory[35996] <=  8'h62;        memory[35997] <=  8'h61;        memory[35998] <=  8'h74;        memory[35999] <=  8'h62;        memory[36000] <=  8'h72;        memory[36001] <=  8'h63;        memory[36002] <=  8'h61;        memory[36003] <=  8'h74;        memory[36004] <=  8'h72;        memory[36005] <=  8'h6e;        memory[36006] <=  8'h62;        memory[36007] <=  8'h61;        memory[36008] <=  8'h63;        memory[36009] <=  8'h61;        memory[36010] <=  8'h74;        memory[36011] <=  8'h79;        memory[36012] <=  8'h73;        memory[36013] <=  8'h6e;        memory[36014] <=  8'h63;        memory[36015] <=  8'h74;        memory[36016] <=  8'h61;        memory[36017] <=  8'h6e;        memory[36018] <=  8'h62;        memory[36019] <=  8'h61;        memory[36020] <=  8'h63;        memory[36021] <=  8'h72;        memory[36022] <=  8'h6e;        memory[36023] <=  8'h74;        memory[36024] <=  8'h61;        memory[36025] <=  8'h62;        memory[36026] <=  8'h74;        memory[36027] <=  8'h6e;        memory[36028] <=  8'h61;        memory[36029] <=  8'h72;        memory[36030] <=  8'h62;        memory[36031] <=  8'h78;        memory[36032] <=  8'h74;        memory[36033] <=  8'h61;        memory[36034] <=  8'h72;        memory[36035] <=  8'h62;        memory[36036] <=  8'h61;        memory[36037] <=  8'h72;        memory[36038] <=  8'h74;        memory[36039] <=  8'h74;        memory[36040] <=  8'h62;        memory[36041] <=  8'h61;        memory[36042] <=  8'h72;        memory[36043] <=  8'h74;        memory[36044] <=  8'h78;        memory[36045] <=  8'h61;        memory[36046] <=  8'h74;        memory[36047] <=  8'h6b;        memory[36048] <=  8'h73;        memory[36049] <=  8'h68;        memory[36050] <=  8'h63;        memory[36051] <=  8'h66;        memory[36052] <=  8'h69;        memory[36053] <=  8'h77;        memory[36054] <=  8'h68;        memory[36055] <=  8'h61;        memory[36056] <=  8'h74;        memory[36057] <=  8'h61;        memory[36058] <=  8'h6e;        memory[36059] <=  8'h61;        memory[36060] <=  8'h62;        memory[36061] <=  8'h61;        memory[36062] <=  8'h63;        memory[36063] <=  8'h61;        memory[36064] <=  8'h74;        memory[36065] <=  8'h61;        memory[36066] <=  8'h62;        memory[36067] <=  8'h61;        memory[36068] <=  8'h72;        memory[36069] <=  8'h63;        memory[36070] <=  8'h61;        memory[36071] <=  8'h68;        memory[36072] <=  8'h64;        memory[36073] <=  8'h75;        memory[36074] <=  8'h63;        memory[36075] <=  8'h74;        memory[36076] <=  8'h61;        memory[36077] <=  8'h64;        memory[36078] <=  8'h61;        memory[36079] <=  8'h61;        memory[36080] <=  8'h63;        memory[36081] <=  8'h61;        memory[36082] <=  8'h72;        memory[36083] <=  8'h63;        memory[36084] <=  8'h74;        memory[36085] <=  8'h72;        memory[36086] <=  8'h63;        memory[36087] <=  8'h61;        memory[36088] <=  8'h74;        memory[36089] <=  8'h72;        memory[36090] <=  8'h63;        memory[36091] <=  8'h61;        memory[36092] <=  8'h74;        memory[36093] <=  8'h63;        memory[36094] <=  8'h62;        memory[36095] <=  8'h61;        memory[36096] <=  8'h74;        memory[36097] <=  8'h62;        memory[36098] <=  8'h72;        memory[36099] <=  8'h63;        memory[36100] <=  8'h61;        memory[36101] <=  8'h74;        memory[36102] <=  8'h72;        memory[36103] <=  8'h6e;        memory[36104] <=  8'h62;        memory[36105] <=  8'h61;        memory[36106] <=  8'h63;        memory[36107] <=  8'h61;        memory[36108] <=  8'h74;        memory[36109] <=  8'h79;        memory[36110] <=  8'h73;        memory[36111] <=  8'h6e;        memory[36112] <=  8'h63;        memory[36113] <=  8'h74;        memory[36114] <=  8'h61;        memory[36115] <=  8'h6e;        memory[36116] <=  8'h62;        memory[36117] <=  8'h61;        memory[36118] <=  8'h63;        memory[36119] <=  8'h72;        memory[36120] <=  8'h6e;        memory[36121] <=  8'h74;        memory[36122] <=  8'h61;        memory[36123] <=  8'h62;        memory[36124] <=  8'h74;        memory[36125] <=  8'h6e;        memory[36126] <=  8'h61;        memory[36127] <=  8'h72;        memory[36128] <=  8'h62;        memory[36129] <=  8'h78;        memory[36130] <=  8'h74;        memory[36131] <=  8'h61;        memory[36132] <=  8'h72;        memory[36133] <=  8'h64;        memory[36134] <=  8'h66;        memory[36135] <=  8'h73;        memory[36136] <=  8'h67;        memory[36137] <=  8'h76;        memory[36138] <=  8'h68;        memory[36139] <=  8'h62;        memory[36140] <=  8'h6b;        memory[36141] <=  8'h6a;        memory[36142] <=  8'h6e;        memory[36143] <=  8'h6d;        memory[36144] <=  8'h62;        memory[36145] <=  8'h76;        memory[36146] <=  8'h78;        memory[36147] <=  8'h63;        memory[36148] <=  8'h73;        memory[36149] <=  8'h66;        memory[36150] <=  8'h72;        memory[36151] <=  8'h74;        memory[36152] <=  8'h79;        memory[36153] <=  8'h75;        memory[36154] <=  8'h6a;        memory[36155] <=  8'h6e;        memory[36156] <=  8'h62;        memory[36157] <=  8'h76;        memory[36158] <=  8'h63;        memory[36159] <=  8'h64;        memory[36160] <=  8'h74;        memory[36161] <=  8'h79;        memory[36162] <=  8'h75;        memory[36163] <=  8'h69;        memory[36164] <=  8'h6b;        memory[36165] <=  8'h6d;        memory[36166] <=  8'h6e;        memory[36167] <=  8'h62;        memory[36168] <=  8'h76;        memory[36169] <=  8'h63;        memory[36170] <=  8'h78;        memory[36171] <=  8'h73;        memory[36172] <=  8'h64;        memory[36173] <=  8'h72;        memory[36174] <=  8'h74;        memory[36175] <=  8'h79;        memory[36176] <=  8'h75;        memory[36177] <=  8'h69;        memory[36178] <=  8'h6b;        memory[36179] <=  8'h6d;        memory[36180] <=  8'h6e;        memory[36181] <=  8'h62;        memory[36182] <=  8'h76;        memory[36183] <=  8'h63;        memory[36184] <=  8'h73;        memory[36185] <=  8'h77;        memory[36186] <=  8'h33;        memory[36187] <=  8'h34;        memory[36188] <=  8'h35;        memory[36189] <=  8'h36;        memory[36190] <=  8'h37;        memory[36191] <=  8'h38;        memory[36192] <=  8'h69;        memory[36193] <=  8'h6b;        memory[36194] <=  8'h6d;        memory[36195] <=  8'h6e;        memory[36196] <=  8'h62;        memory[36197] <=  8'h76;        memory[36198] <=  8'h63;        memory[36199] <=  8'h64;        memory[36200] <=  8'h65;        memory[36201] <=  8'h72;        memory[36202] <=  8'h36;        memory[36203] <=  8'h37;        memory[36204] <=  8'h38;        memory[36205] <=  8'h69;        memory[36206] <=  8'h6f;        memory[36207] <=  8'h6b;        memory[36208] <=  8'h6a;        memory[36209] <=  8'h6e;        memory[36210] <=  8'h62;        memory[36211] <=  8'h76;        memory[36212] <=  8'h63;        memory[36213] <=  8'h64;        memory[36214] <=  8'h72;        memory[36215] <=  8'h74;        memory[36216] <=  8'h79;        memory[36217] <=  8'h75;        memory[36218] <=  8'h73;        memory[36219] <=  8'h6a;        memory[36220] <=  8'h63;        memory[36221] <=  8'h6e;        memory[36222] <=  8'h62;        memory[36223] <=  8'h64;        memory[36224] <=  8'h66;        memory[36225] <=  8'h73;        memory[36226] <=  8'h74;        memory[36227] <=  8'h79;        memory[36228] <=  8'h75;        memory[36229] <=  8'h61;        memory[36230] <=  8'h69;        memory[36231] <=  8'h6b;        memory[36232] <=  8'h78;        memory[36233] <=  8'h6d;        memory[36234] <=  8'h6e;        memory[36235] <=  8'h73;        memory[36236] <=  8'h6a;        memory[36237] <=  8'h6f;        memory[36238] <=  8'h64;        memory[36239] <=  8'h6c;        memory[36240] <=  8'h63;        memory[36241] <=  8'h78;        memory[36242] <=  8'h62;        memory[36243] <=  8'h61;        memory[36244] <=  8'h72;        memory[36245] <=  8'h74;        memory[36246] <=  8'h78;        memory[36247] <=  8'h61;        memory[36248] <=  8'h74;        memory[36249] <=  8'h6b;        memory[36250] <=  8'h73;        memory[36251] <=  8'h68;        memory[36252] <=  8'h63;        memory[36253] <=  8'h66;        memory[36254] <=  8'h69;        memory[36255] <=  8'h77;        memory[36256] <=  8'h68;        memory[36257] <=  8'h61;        memory[36258] <=  8'h74;        memory[36259] <=  8'h61;        memory[36260] <=  8'h6e;        memory[36261] <=  8'h61;        memory[36262] <=  8'h62;        memory[36263] <=  8'h61;        memory[36264] <=  8'h63;        memory[36265] <=  8'h61;        memory[36266] <=  8'h74;        memory[36267] <=  8'h61;        memory[36268] <=  8'h62;        memory[36269] <=  8'h61;        memory[36270] <=  8'h72;        memory[36271] <=  8'h63;        memory[36272] <=  8'h61;        memory[36273] <=  8'h68;        memory[36274] <=  8'h64;        memory[36275] <=  8'h75;        memory[36276] <=  8'h63;        memory[36277] <=  8'h74;        memory[36278] <=  8'h61;        memory[36279] <=  8'h64;        memory[36280] <=  8'h61;        memory[36281] <=  8'h61;        memory[36282] <=  8'h63;        memory[36283] <=  8'h61;        memory[36284] <=  8'h72;        memory[36285] <=  8'h62;        memory[36286] <=  8'h61;        memory[36287] <=  8'h72;        memory[36288] <=  8'h74;        memory[36289] <=  8'h78;        memory[36290] <=  8'h61;        memory[36291] <=  8'h74;        memory[36292] <=  8'h6b;        memory[36293] <=  8'h73;        memory[36294] <=  8'h68;        memory[36295] <=  8'h63;        memory[36296] <=  8'h66;        memory[36297] <=  8'h69;        memory[36298] <=  8'h77;        memory[36299] <=  8'h68;        memory[36300] <=  8'h61;        memory[36301] <=  8'h74;        memory[36302] <=  8'h61;        memory[36303] <=  8'h6e;        memory[36304] <=  8'h61;        memory[36305] <=  8'h62;        memory[36306] <=  8'h61;        memory[36307] <=  8'h63;        memory[36308] <=  8'h61;        memory[36309] <=  8'h74;        memory[36310] <=  8'h61;        memory[36311] <=  8'h62;        memory[36312] <=  8'h61;        memory[36313] <=  8'h72;        memory[36314] <=  8'h63;        memory[36315] <=  8'h61;        memory[36316] <=  8'h68;        memory[36317] <=  8'h64;        memory[36318] <=  8'h75;        memory[36319] <=  8'h63;        memory[36320] <=  8'h74;        memory[36321] <=  8'h61;        memory[36322] <=  8'h64;        memory[36323] <=  8'h61;        memory[36324] <=  8'h61;        memory[36325] <=  8'h63;        memory[36326] <=  8'h61;        memory[36327] <=  8'h72;        memory[36328] <=  8'h62;        memory[36329] <=  8'h61;        memory[36330] <=  8'h72;        memory[36331] <=  8'h74;        memory[36332] <=  8'h78;        memory[36333] <=  8'h61;        memory[36334] <=  8'h74;        memory[36335] <=  8'h6b;        memory[36336] <=  8'h73;        memory[36337] <=  8'h68;        memory[36338] <=  8'h63;        memory[36339] <=  8'h66;        memory[36340] <=  8'h69;        memory[36341] <=  8'h77;        memory[36342] <=  8'h68;        memory[36343] <=  8'h61;        memory[36344] <=  8'h74;        memory[36345] <=  8'h61;        memory[36346] <=  8'h6e;        memory[36347] <=  8'h61;        memory[36348] <=  8'h62;        memory[36349] <=  8'h61;        memory[36350] <=  8'h63;        memory[36351] <=  8'h61;        memory[36352] <=  8'h74;        memory[36353] <=  8'h61;        memory[36354] <=  8'h62;        memory[36355] <=  8'h61;        memory[36356] <=  8'h72;        memory[36357] <=  8'h63;        memory[36358] <=  8'h61;        memory[36359] <=  8'h68;        memory[36360] <=  8'h64;        memory[36361] <=  8'h75;        memory[36362] <=  8'h63;        memory[36363] <=  8'h74;        memory[36364] <=  8'h61;        memory[36365] <=  8'h64;        memory[36366] <=  8'h61;        memory[36367] <=  8'h61;        memory[36368] <=  8'h63;        memory[36369] <=  8'h61;        memory[36370] <=  8'h72;        memory[36371] <=  8'h62;        memory[36372] <=  8'h61;        memory[36373] <=  8'h72;        memory[36374] <=  8'h74;        memory[36375] <=  8'h78;        memory[36376] <=  8'h61;        memory[36377] <=  8'h74;        memory[36378] <=  8'h6b;        memory[36379] <=  8'h73;        memory[36380] <=  8'h68;        memory[36381] <=  8'h63;        memory[36382] <=  8'h66;        memory[36383] <=  8'h69;        memory[36384] <=  8'h77;        memory[36385] <=  8'h68;        memory[36386] <=  8'h61;        memory[36387] <=  8'h74;        memory[36388] <=  8'h61;        memory[36389] <=  8'h6e;        memory[36390] <=  8'h61;        memory[36391] <=  8'h62;        memory[36392] <=  8'h61;        memory[36393] <=  8'h63;        memory[36394] <=  8'h61;        memory[36395] <=  8'h74;        memory[36396] <=  8'h61;        memory[36397] <=  8'h62;        memory[36398] <=  8'h61;        memory[36399] <=  8'h72;        memory[36400] <=  8'h63;        memory[36401] <=  8'h61;        memory[36402] <=  8'h68;        memory[36403] <=  8'h64;        memory[36404] <=  8'h75;        memory[36405] <=  8'h63;        memory[36406] <=  8'h74;        memory[36407] <=  8'h61;        memory[36408] <=  8'h64;        memory[36409] <=  8'h61;        memory[36410] <=  8'h61;        memory[36411] <=  8'h63;        memory[36412] <=  8'h61;        memory[36413] <=  8'h72;        memory[36414] <=  8'h62;        memory[36415] <=  8'h61;        memory[36416] <=  8'h72;        memory[36417] <=  8'h74;        memory[36418] <=  8'h78;        memory[36419] <=  8'h61;        memory[36420] <=  8'h74;        memory[36421] <=  8'h6b;        memory[36422] <=  8'h73;        memory[36423] <=  8'h68;        memory[36424] <=  8'h63;        memory[36425] <=  8'h66;        memory[36426] <=  8'h69;        memory[36427] <=  8'h77;        memory[36428] <=  8'h68;        memory[36429] <=  8'h61;        memory[36430] <=  8'h74;        memory[36431] <=  8'h61;        memory[36432] <=  8'h6e;        memory[36433] <=  8'h61;        memory[36434] <=  8'h62;        memory[36435] <=  8'h61;        memory[36436] <=  8'h63;        memory[36437] <=  8'h61;        memory[36438] <=  8'h74;        memory[36439] <=  8'h61;        memory[36440] <=  8'h62;        memory[36441] <=  8'h61;        memory[36442] <=  8'h72;        memory[36443] <=  8'h63;        memory[36444] <=  8'h61;        memory[36445] <=  8'h68;        memory[36446] <=  8'h64;        memory[36447] <=  8'h75;        memory[36448] <=  8'h63;        memory[36449] <=  8'h74;        memory[36450] <=  8'h61;        memory[36451] <=  8'h64;        memory[36452] <=  8'h61;        memory[36453] <=  8'h61;        memory[36454] <=  8'h63;        memory[36455] <=  8'h61;        memory[36456] <=  8'h72;        memory[36457] <=  8'h62;        memory[36458] <=  8'h61;        memory[36459] <=  8'h72;        memory[36460] <=  8'h74;        memory[36461] <=  8'h78;        memory[36462] <=  8'h61;        memory[36463] <=  8'h74;        memory[36464] <=  8'h6b;        memory[36465] <=  8'h73;        memory[36466] <=  8'h68;        memory[36467] <=  8'h63;        memory[36468] <=  8'h66;        memory[36469] <=  8'h69;        memory[36470] <=  8'h77;        memory[36471] <=  8'h68;        memory[36472] <=  8'h61;        memory[36473] <=  8'h74;        memory[36474] <=  8'h61;        memory[36475] <=  8'h6e;        memory[36476] <=  8'h61;        memory[36477] <=  8'h62;        memory[36478] <=  8'h61;        memory[36479] <=  8'h63;        memory[36480] <=  8'h61;        memory[36481] <=  8'h74;        memory[36482] <=  8'h61;        memory[36483] <=  8'h62;        memory[36484] <=  8'h61;        memory[36485] <=  8'h72;        memory[36486] <=  8'h63;        memory[36487] <=  8'h61;        memory[36488] <=  8'h68;        memory[36489] <=  8'h64;        memory[36490] <=  8'h75;        memory[36491] <=  8'h63;        memory[36492] <=  8'h74;        memory[36493] <=  8'h61;        memory[36494] <=  8'h64;        memory[36495] <=  8'h61;        memory[36496] <=  8'h61;        memory[36497] <=  8'h63;        memory[36498] <=  8'h61;        memory[36499] <=  8'h72;        memory[36500] <=  8'h62;        memory[36501] <=  8'h61;        memory[36502] <=  8'h72;        memory[36503] <=  8'h74;        memory[36504] <=  8'h78;        memory[36505] <=  8'h61;        memory[36506] <=  8'h74;        memory[36507] <=  8'h6b;        memory[36508] <=  8'h73;        memory[36509] <=  8'h68;        memory[36510] <=  8'h63;        memory[36511] <=  8'h66;        memory[36512] <=  8'h69;        memory[36513] <=  8'h77;        memory[36514] <=  8'h68;        memory[36515] <=  8'h61;        memory[36516] <=  8'h74;        memory[36517] <=  8'h61;        memory[36518] <=  8'h6e;        memory[36519] <=  8'h61;        memory[36520] <=  8'h62;        memory[36521] <=  8'h61;        memory[36522] <=  8'h63;        memory[36523] <=  8'h61;        memory[36524] <=  8'h74;        memory[36525] <=  8'h61;        memory[36526] <=  8'h62;        memory[36527] <=  8'h61;        memory[36528] <=  8'h72;        memory[36529] <=  8'h63;        memory[36530] <=  8'h61;        memory[36531] <=  8'h68;        memory[36532] <=  8'h64;        memory[36533] <=  8'h75;        memory[36534] <=  8'h63;        memory[36535] <=  8'h74;        memory[36536] <=  8'h61;        memory[36537] <=  8'h64;        memory[36538] <=  8'h61;        memory[36539] <=  8'h61;        memory[36540] <=  8'h63;        memory[36541] <=  8'h61;        memory[36542] <=  8'h72;        memory[36543] <=  8'h62;        memory[36544] <=  8'h61;        memory[36545] <=  8'h72;        memory[36546] <=  8'h74;        memory[36547] <=  8'h78;        memory[36548] <=  8'h61;        memory[36549] <=  8'h74;        memory[36550] <=  8'h6b;        memory[36551] <=  8'h73;        memory[36552] <=  8'h68;        memory[36553] <=  8'h63;        memory[36554] <=  8'h66;        memory[36555] <=  8'h69;        memory[36556] <=  8'h77;        memory[36557] <=  8'h68;        memory[36558] <=  8'h61;        memory[36559] <=  8'h74;        memory[36560] <=  8'h61;        memory[36561] <=  8'h6e;        memory[36562] <=  8'h61;        memory[36563] <=  8'h62;        memory[36564] <=  8'h61;        memory[36565] <=  8'h63;        memory[36566] <=  8'h61;        memory[36567] <=  8'h74;        memory[36568] <=  8'h61;        memory[36569] <=  8'h62;        memory[36570] <=  8'h61;        memory[36571] <=  8'h72;        memory[36572] <=  8'h63;        memory[36573] <=  8'h61;        memory[36574] <=  8'h68;        memory[36575] <=  8'h64;        memory[36576] <=  8'h75;        memory[36577] <=  8'h63;        memory[36578] <=  8'h74;        memory[36579] <=  8'h61;        memory[36580] <=  8'h64;        memory[36581] <=  8'h61;        memory[36582] <=  8'h61;        memory[36583] <=  8'h63;        memory[36584] <=  8'h61;        memory[36585] <=  8'h72;        memory[36586] <=  8'h62;        memory[36587] <=  8'h61;        memory[36588] <=  8'h72;        memory[36589] <=  8'h74;        memory[36590] <=  8'h78;        memory[36591] <=  8'h61;        memory[36592] <=  8'h74;        memory[36593] <=  8'h6b;        memory[36594] <=  8'h73;        memory[36595] <=  8'h68;        memory[36596] <=  8'h63;        memory[36597] <=  8'h66;        memory[36598] <=  8'h69;        memory[36599] <=  8'h77;        memory[36600] <=  8'h68;        memory[36601] <=  8'h61;        memory[36602] <=  8'h74;        memory[36603] <=  8'h61;        memory[36604] <=  8'h6e;        memory[36605] <=  8'h61;        memory[36606] <=  8'h62;        memory[36607] <=  8'h61;        memory[36608] <=  8'h63;        memory[36609] <=  8'h61;        memory[36610] <=  8'h74;        memory[36611] <=  8'h61;        memory[36612] <=  8'h62;        memory[36613] <=  8'h61;        memory[36614] <=  8'h72;        memory[36615] <=  8'h63;        memory[36616] <=  8'h61;        memory[36617] <=  8'h68;        memory[36618] <=  8'h64;        memory[36619] <=  8'h75;        memory[36620] <=  8'h63;        memory[36621] <=  8'h74;        memory[36622] <=  8'h61;        memory[36623] <=  8'h64;        memory[36624] <=  8'h61;        memory[36625] <=  8'h61;        memory[36626] <=  8'h63;        memory[36627] <=  8'h61;        memory[36628] <=  8'h72;        memory[36629] <=  8'h62;        memory[36630] <=  8'h61;        memory[36631] <=  8'h72;        memory[36632] <=  8'h74;        memory[36633] <=  8'h74;        memory[36634] <=  8'h62;        memory[36635] <=  8'h61;        memory[36636] <=  8'h72;        memory[36637] <=  8'h74;        memory[36638] <=  8'h78;        memory[36639] <=  8'h61;        memory[36640] <=  8'h74;        memory[36641] <=  8'h6b;        memory[36642] <=  8'h73;        memory[36643] <=  8'h68;        memory[36644] <=  8'h63;        memory[36645] <=  8'h66;        memory[36646] <=  8'h69;        memory[36647] <=  8'h77;        memory[36648] <=  8'h68;        memory[36649] <=  8'h61;        memory[36650] <=  8'h74;        memory[36651] <=  8'h61;        memory[36652] <=  8'h6e;        memory[36653] <=  8'h61;        memory[36654] <=  8'h62;        memory[36655] <=  8'h61;        memory[36656] <=  8'h63;        memory[36657] <=  8'h61;        memory[36658] <=  8'h74;        memory[36659] <=  8'h61;        memory[36660] <=  8'h62;        memory[36661] <=  8'h61;        memory[36662] <=  8'h72;        memory[36663] <=  8'h63;        memory[36664] <=  8'h61;        memory[36665] <=  8'h68;        memory[36666] <=  8'h64;        memory[36667] <=  8'h75;        memory[36668] <=  8'h63;        memory[36669] <=  8'h74;        memory[36670] <=  8'h61;        memory[36671] <=  8'h64;        memory[36672] <=  8'h61;        memory[36673] <=  8'h61;        memory[36674] <=  8'h63;        memory[36675] <=  8'h61;        memory[36676] <=  8'h72;        memory[36677] <=  8'h63;        memory[36678] <=  8'h74;        memory[36679] <=  8'h72;        memory[36680] <=  8'h63;        memory[36681] <=  8'h61;        memory[36682] <=  8'h74;        memory[36683] <=  8'h72;        memory[36684] <=  8'h63;        memory[36685] <=  8'h61;        memory[36686] <=  8'h74;        memory[36687] <=  8'h63;        memory[36688] <=  8'h62;        memory[36689] <=  8'h61;        memory[36690] <=  8'h74;        memory[36691] <=  8'h62;        memory[36692] <=  8'h72;        memory[36693] <=  8'h63;        memory[36694] <=  8'h61;        memory[36695] <=  8'h72;        memory[36696] <=  8'h62;        memory[36697] <=  8'h78;        memory[36698] <=  8'h74;        memory[36699] <=  8'h61;        memory[36700] <=  8'h72;        memory[36701] <=  8'h64;        memory[36702] <=  8'h66;        memory[36703] <=  8'h73;        memory[36704] <=  8'h67;        memory[36705] <=  8'h76;        memory[36706] <=  8'h68;        memory[36707] <=  8'h62;        memory[36708] <=  8'h6b;        memory[36709] <=  8'h6a;        memory[36710] <=  8'h6e;        memory[36711] <=  8'h6d;        memory[36712] <=  8'h62;        memory[36713] <=  8'h76;        memory[36714] <=  8'h78;        memory[36715] <=  8'h63;        memory[36716] <=  8'h73;        memory[36717] <=  8'h66;        memory[36718] <=  8'h72;        memory[36719] <=  8'h74;        memory[36720] <=  8'h79;        memory[36721] <=  8'h75;        memory[36722] <=  8'h6a;        memory[36723] <=  8'h6e;        memory[36724] <=  8'h62;        memory[36725] <=  8'h76;        memory[36726] <=  8'h63;        memory[36727] <=  8'h64;        memory[36728] <=  8'h74;        memory[36729] <=  8'h79;        memory[36730] <=  8'h75;        memory[36731] <=  8'h69;        memory[36732] <=  8'h6b;        memory[36733] <=  8'h6d;        memory[36734] <=  8'h6e;        memory[36735] <=  8'h62;        memory[36736] <=  8'h76;        memory[36737] <=  8'h63;        memory[36738] <=  8'h78;        memory[36739] <=  8'h73;        memory[36740] <=  8'h64;        memory[36741] <=  8'h72;        memory[36742] <=  8'h74;        memory[36743] <=  8'h79;        memory[36744] <=  8'h75;        memory[36745] <=  8'h69;        memory[36746] <=  8'h6b;        memory[36747] <=  8'h6d;        memory[36748] <=  8'h6e;        memory[36749] <=  8'h62;        memory[36750] <=  8'h76;        memory[36751] <=  8'h63;        memory[36752] <=  8'h73;        memory[36753] <=  8'h77;        memory[36754] <=  8'h33;        memory[36755] <=  8'h34;        memory[36756] <=  8'h35;        memory[36757] <=  8'h36;        memory[36758] <=  8'h37;        memory[36759] <=  8'h38;        memory[36760] <=  8'h69;        memory[36761] <=  8'h6b;        memory[36762] <=  8'h6d;        memory[36763] <=  8'h6e;        memory[36764] <=  8'h62;        memory[36765] <=  8'h76;        memory[36766] <=  8'h63;        memory[36767] <=  8'h64;        memory[36768] <=  8'h65;        memory[36769] <=  8'h72;        memory[36770] <=  8'h36;        memory[36771] <=  8'h37;        memory[36772] <=  8'h38;        memory[36773] <=  8'h69;        memory[36774] <=  8'h6f;        memory[36775] <=  8'h6b;        memory[36776] <=  8'h6a;        memory[36777] <=  8'h6e;        memory[36778] <=  8'h62;        memory[36779] <=  8'h76;        memory[36780] <=  8'h63;        memory[36781] <=  8'h64;        memory[36782] <=  8'h72;        memory[36783] <=  8'h74;        memory[36784] <=  8'h79;        memory[36785] <=  8'h75;        memory[36786] <=  8'h73;        memory[36787] <=  8'h6a;        memory[36788] <=  8'h63;        memory[36789] <=  8'h6e;        memory[36790] <=  8'h62;        memory[36791] <=  8'h64;        memory[36792] <=  8'h66;        memory[36793] <=  8'h73;        memory[36794] <=  8'h74;        memory[36795] <=  8'h79;        memory[36796] <=  8'h75;        memory[36797] <=  8'h61;        memory[36798] <=  8'h69;        memory[36799] <=  8'h6b;        memory[36800] <=  8'h78;        memory[36801] <=  8'h6d;        memory[36802] <=  8'h6e;        memory[36803] <=  8'h73;        memory[36804] <=  8'h6a;        memory[36805] <=  8'h6f;        memory[36806] <=  8'h64;        memory[36807] <=  8'h6c;        memory[36808] <=  8'h63;        memory[36809] <=  8'h78;        memory[36810] <=  8'h2c;        memory[36811] <=  8'h6d;        memory[36812] <=  8'h73;        memory[36813] <=  8'h6b;        memory[36814] <=  8'h64;        memory[36815] <=  8'h6c;        memory[36816] <=  8'h70;        memory[36817] <=  8'h5b;        memory[36818] <=  8'h3b;        memory[36819] <=  8'h73;        memory[36820] <=  8'h6c;        memory[36821] <=  8'h64;        memory[36822] <=  8'h70;        memory[36823] <=  8'h76;        memory[36824] <=  8'h63;        memory[36825] <=  8'h5b;        memory[36826] <=  8'h78;        memory[36827] <=  8'h76;        memory[36828] <=  8'h63;        memory[36829] <=  8'h5b;        memory[36830] <=  8'h78;        memory[36831] <=  8'h70;        memory[36832] <=  8'h6f;        memory[36833] <=  8'h20;        memory[36834] <=  8'h62;        memory[36835] <=  8'h61;        memory[36836] <=  8'h72;        memory[36837] <=  8'h74;        memory[36838] <=  8'h74;        memory[36839] <=  8'h62;        memory[36840] <=  8'h61;        memory[36841] <=  8'h72;        memory[36842] <=  8'h74;        memory[36843] <=  8'h78;        memory[36844] <=  8'h61;        memory[36845] <=  8'h74;        memory[36846] <=  8'h6b;        memory[36847] <=  8'h73;        memory[36848] <=  8'h68;        memory[36849] <=  8'h63;        memory[36850] <=  8'h66;        memory[36851] <=  8'h69;        memory[36852] <=  8'h77;        memory[36853] <=  8'h68;        memory[36854] <=  8'h61;        memory[36855] <=  8'h69;        memory[36856] <=  8'h6a;        memory[36857] <=  8'h78;        memory[36858] <=  8'h5d;        memory[36859] <=  8'h65;        memory[36860] <=  8'h6b;        memory[36861] <=  8'h6f;        memory[36862] <=  8'h39;        memory[36863] <=  8'h64;        memory[36864] <=  8'h75;        memory[36865] <=  8'h38;        memory[36866] <=  8'h79;        memory[36867] <=  8'h20;        memory[36868] <=  8'h37;        memory[36869] <=  8'h63;        memory[36870] <=  8'h67;        memory[36871] <=  8'h78;        memory[36872] <=  8'h63;        memory[36873] <=  8'h75;        memory[36874] <=  8'h68;        memory[36875] <=  8'h69;        memory[36876] <=  8'h6a;        memory[36877] <=  8'h77;        memory[36878] <=  8'h69;        memory[36879] <=  8'h64;        memory[36880] <=  8'h66;        memory[36881] <=  8'h68;        memory[36882] <=  8'h75;        memory[36883] <=  8'h76;        memory[36884] <=  8'h64;        memory[36885] <=  8'h62;        memory[36886] <=  8'h66;        memory[36887] <=  8'h6a;        memory[36888] <=  8'h6e;        memory[36889] <=  8'h6b;        memory[36890] <=  8'h6a;        memory[36891] <=  8'h65;        memory[36892] <=  8'h38;        memory[36893] <=  8'h66;        memory[36894] <=  8'h37;        memory[36895] <=  8'h67;        memory[36896] <=  8'h79;        memory[36897] <=  8'h76;        memory[36898] <=  8'h63;        memory[36899] <=  8'h68;        memory[36900] <=  8'h69;        memory[36901] <=  8'h6a;        memory[36902] <=  8'h33;        memory[36903] <=  8'h65;        memory[36904] <=  8'h67;        memory[36905] <=  8'h79;        memory[36906] <=  8'h72;        memory[36907] <=  8'h64;        memory[36908] <=  8'h62;        memory[36909] <=  8'h6e;        memory[36910] <=  8'h63;        memory[36911] <=  8'h7a;        memory[36912] <=  8'h6a;        memory[36913] <=  8'h6f;        memory[36914] <=  8'h66;        memory[36915] <=  8'h78;        memory[36916] <=  8'h6a;        memory[36917] <=  8'h69;        memory[36918] <=  8'h63;        memory[36919] <=  8'h68;        memory[36920] <=  8'h62;        memory[36921] <=  8'h6e;        memory[36922] <=  8'h6d;        memory[36923] <=  8'h63;        memory[36924] <=  8'h73;        memory[36925] <=  8'h6c;        memory[36926] <=  8'h6b;        memory[36927] <=  8'h6a;        memory[36928] <=  8'h69;        memory[36929] <=  8'h68;        memory[36930] <=  8'h76;        memory[36931] <=  8'h75;        memory[36932] <=  8'h69;        memory[36933] <=  8'h64;        memory[36934] <=  8'h68;        memory[36935] <=  8'h75;        memory[36936] <=  8'h67;        memory[36937] <=  8'h79;        memory[36938] <=  8'h62;        memory[36939] <=  8'h68;        memory[36940] <=  8'h65;        memory[36941] <=  8'h6a;        memory[36942] <=  8'h72;        memory[36943] <=  8'h6b;        memory[36944] <=  8'h6a;        memory[36945] <=  8'h6f;        memory[36946] <=  8'h64;        memory[36947] <=  8'h67;        memory[36948] <=  8'h69;        memory[36949] <=  8'h75;        memory[36950] <=  8'h69;        memory[36951] <=  8'h67;        memory[36952] <=  8'h76;        memory[36953] <=  8'h79;        memory[36954] <=  8'h75;        memory[36955] <=  8'h67;        memory[36956] <=  8'h78;        memory[36957] <=  8'h68;        memory[36958] <=  8'h63;        memory[36959] <=  8'h20;        memory[36960] <=  8'h20;        memory[36961] <=  8'h20;        memory[36962] <=  8'h78;        memory[36963] <=  8'h76;        memory[36964] <=  8'h20;        memory[36965] <=  8'h63;        memory[36966] <=  8'h78;        memory[36967] <=  8'h67;        memory[36968] <=  8'h79;        memory[36969] <=  8'h63;        memory[36970] <=  8'h75;        memory[36971] <=  8'h68;        memory[36972] <=  8'h6a;        memory[36973] <=  8'h6b;        memory[36974] <=  8'h61;        memory[36975] <=  8'h6c;        memory[36976] <=  8'h78;        memory[36977] <=  8'h76;        memory[36978] <=  8'h70;        memory[36979] <=  8'h6f;        memory[36980] <=  8'h69;        memory[36981] <=  8'h6a;        memory[36982] <=  8'h69;        memory[36983] <=  8'h68;        memory[36984] <=  8'h6a;        memory[36985] <=  8'h62;        memory[36986] <=  8'h77;        memory[36987] <=  8'h65;        memory[36988] <=  8'h6e;        memory[36989] <=  8'h61;        memory[36990] <=  8'h66;        memory[36991] <=  8'h6d;        memory[36992] <=  8'h64;        memory[36993] <=  8'h6b;        memory[36994] <=  8'h6d;        memory[36995] <=  8'h76;        memory[36996] <=  8'h6c;        memory[36997] <=  8'h63;        memory[36998] <=  8'h6f;        memory[36999] <=  8'h64;        memory[37000] <=  8'h69;        memory[37001] <=  8'h75;        memory[37002] <=  8'h68;        memory[37003] <=  8'h73;        memory[37004] <=  8'h66;        memory[37005] <=  8'h65;        memory[37006] <=  8'h62;        memory[37007] <=  8'h6e;        memory[37008] <=  8'h64;        memory[37009] <=  8'h73;        memory[37010] <=  8'h63;        memory[37011] <=  8'h6b;        memory[37012] <=  8'h20;        memory[37013] <=  8'h78;        memory[37014] <=  8'h6a;        memory[37015] <=  8'h78;        memory[37016] <=  8'h63;        memory[37017] <=  8'h73;        memory[37018] <=  8'h64;        memory[37019] <=  8'h66;        memory[37020] <=  8'h6b;        memory[37021] <=  8'h64;        memory[37022] <=  8'h6e;        memory[37023] <=  8'h6d;        memory[37024] <=  8'h64;        memory[37025] <=  8'h73;        memory[37026] <=  8'h63;        memory[37027] <=  8'h6b;        memory[37028] <=  8'h78;        memory[37029] <=  8'h6c;        memory[37030] <=  8'h6f;        memory[37031] <=  8'h66;        memory[37032] <=  8'h6a;        memory[37033] <=  8'h69;        memory[37034] <=  8'h61;        memory[37035] <=  8'h62;        memory[37036] <=  8'h6e;        memory[37037] <=  8'h20;        memory[37038] <=  8'h78;        memory[37039] <=  8'h6b;        memory[37040] <=  8'h6d;        memory[37041] <=  8'h20;        memory[37042] <=  8'h6f;        memory[37043] <=  8'h63;        memory[37044] <=  8'h76;        memory[37045] <=  8'h73;        memory[37046] <=  8'h64;        memory[37047] <=  8'h69;        memory[37048] <=  8'h66;        memory[37049] <=  8'h68;        memory[37050] <=  8'h65;        memory[37051] <=  8'h71;        memory[37052] <=  8'h6a;        memory[37053] <=  8'h77;        memory[37054] <=  8'h62;        memory[37055] <=  8'h65;        memory[37056] <=  8'h6e;        memory[37057] <=  8'h20;        memory[37058] <=  8'h6d;        memory[37059] <=  8'h64;        memory[37060] <=  8'h73;        memory[37061] <=  8'h6c;        memory[37062] <=  8'h76;        memory[37063] <=  8'h6b;        memory[37064] <=  8'h63;        memory[37065] <=  8'h78;        memory[37066] <=  8'h20;        memory[37067] <=  8'h6f;        memory[37068] <=  8'h78;        memory[37069] <=  8'h69;        memory[37070] <=  8'h63;        memory[37071] <=  8'h6a;        memory[37072] <=  8'h76;        memory[37073] <=  8'h64;        memory[37074] <=  8'h66;        memory[37075] <=  8'h65;        memory[37076] <=  8'h71;        memory[37077] <=  8'h6e;        memory[37078] <=  8'h20;        memory[37079] <=  8'h64;        memory[37080] <=  8'h6d;        memory[37081] <=  8'h73;        memory[37082] <=  8'h6c;        memory[37083] <=  8'h63;        memory[37084] <=  8'h78;        memory[37085] <=  8'h6b;        memory[37086] <=  8'h20;        memory[37087] <=  8'h6f;        memory[37088] <=  8'h78;        memory[37089] <=  8'h63;        memory[37090] <=  8'h76;        memory[37091] <=  8'h6a;        memory[37092] <=  8'h64;        memory[37093] <=  8'h62;        memory[37094] <=  8'h71;        memory[37095] <=  8'h77;        memory[37096] <=  8'h65;        memory[37097] <=  8'h6e;        memory[37098] <=  8'h6d;        memory[37099] <=  8'h64;        memory[37100] <=  8'h6c;        memory[37101] <=  8'h73;        memory[37102] <=  8'h2c;        memory[37103] <=  8'h76;        memory[37104] <=  8'h63;        memory[37105] <=  8'h78;        memory[37106] <=  8'h20;        memory[37107] <=  8'h63;        memory[37108] <=  8'h6f;        memory[37109] <=  8'h69;        memory[37110] <=  8'h76;        memory[37111] <=  8'h68;        memory[37112] <=  8'h73;        memory[37113] <=  8'h64;        memory[37114] <=  8'h62;        memory[37115] <=  8'h71;        memory[37116] <=  8'h77;        memory[37117] <=  8'h65;        memory[37118] <=  8'h6e;        memory[37119] <=  8'h64;        memory[37120] <=  8'h6b;        memory[37121] <=  8'h73;        memory[37122] <=  8'h76;        memory[37123] <=  8'h6f;        memory[37124] <=  8'h63;        memory[37125] <=  8'h20;        memory[37126] <=  8'h76;        memory[37127] <=  8'h69;        memory[37128] <=  8'h75;        memory[37129] <=  8'h69;        memory[37130] <=  8'h68;        memory[37131] <=  8'h63;        memory[37132] <=  8'h78;        memory[37133] <=  8'h69;        memory[37134] <=  8'h6f;        memory[37135] <=  8'h76;        memory[37136] <=  8'h73;        memory[37137] <=  8'h64;        memory[37138] <=  8'h61;        memory[37139] <=  8'h64;        memory[37140] <=  8'h6e;        memory[37141] <=  8'h77;        memory[37142] <=  8'h71;        memory[37143] <=  8'h6b;        memory[37144] <=  8'h6c;        memory[37145] <=  8'h73;        memory[37146] <=  8'h76;        memory[37147] <=  8'h6e;        memory[37148] <=  8'h62;        memory[37149] <=  8'h20;        memory[37150] <=  8'h64;        memory[37151] <=  8'h66;        memory[37152] <=  8'h6a;        memory[37153] <=  8'h6b;        memory[37154] <=  8'h71;        memory[37155] <=  8'h64;        memory[37156] <=  8'h77;        memory[37157] <=  8'h65;        memory[37158] <=  8'h6e;        memory[37159] <=  8'h62;        memory[37160] <=  8'h20;        memory[37161] <=  8'h64;        memory[37162] <=  8'h73;        memory[37163] <=  8'h76;        memory[37164] <=  8'h68;        memory[37165] <=  8'h64;        memory[37166] <=  8'h61;        memory[37167] <=  8'h71;        memory[37168] <=  8'h77;        memory[37169] <=  8'h6a;        memory[37170] <=  8'h65;        memory[37171] <=  8'h6e;        memory[37172] <=  8'h64;        memory[37173] <=  8'h20;        memory[37174] <=  8'h61;        memory[37175] <=  8'h63;        memory[37176] <=  8'h62;        memory[37177] <=  8'h68;        memory[37178] <=  8'h64;        memory[37179] <=  8'h61;        memory[37180] <=  8'h77;        memory[37181] <=  8'h71;        memory[37182] <=  8'h6e;        memory[37183] <=  8'h20;        memory[37184] <=  8'h62;        memory[37185] <=  8'h73;        memory[37186] <=  8'h76;        memory[37187] <=  8'h61;        memory[37188] <=  8'h67;        memory[37189] <=  8'h76;        memory[37190] <=  8'h68;        memory[37191] <=  8'h67;        memory[37192] <=  8'h61;        memory[37193] <=  8'h73;        memory[37194] <=  8'h6a;        memory[37195] <=  8'h6b;        memory[37196] <=  8'h63;        memory[37197] <=  8'h78;        memory[37198] <=  8'h76;        memory[37199] <=  8'h6e;        memory[37200] <=  8'h73;        memory[37201] <=  8'h64;        memory[37202] <=  8'h20;        memory[37203] <=  8'h66;        memory[37204] <=  8'h62;        memory[37205] <=  8'h64;        memory[37206] <=  8'h61;        memory[37207] <=  8'h73;        memory[37208] <=  8'h76;        memory[37209] <=  8'h67;        memory[37210] <=  8'h63;        memory[37211] <=  8'h79;        memory[37212] <=  8'h7a;        memory[37213] <=  8'h78;        memory[37214] <=  8'h79;        memory[37215] <=  8'h75;        memory[37216] <=  8'h20;        memory[37217] <=  8'h69;        memory[37218] <=  8'h6a;        memory[37219] <=  8'h64;        memory[37220] <=  8'h66;        memory[37221] <=  8'h6b;        memory[37222] <=  8'h61;        memory[37223] <=  8'h64;        memory[37224] <=  8'h63;        memory[37225] <=  8'h78;        memory[37226] <=  8'h68;        memory[37227] <=  8'h20;        memory[37228] <=  8'h67;        memory[37229] <=  8'h61;        memory[37230] <=  8'h68;        memory[37231] <=  8'h75;        memory[37232] <=  8'h64;        memory[37233] <=  8'h73;        memory[37234] <=  8'h69;        memory[37235] <=  8'h6a;        memory[37236] <=  8'h61;        memory[37237] <=  8'h6b;        memory[37238] <=  8'h63;        memory[37239] <=  8'h62;        memory[37240] <=  8'h61;        memory[37241] <=  8'h72;        memory[37242] <=  8'h73;        memory[37243] <=  8'h68;        memory[37244] <=  8'h64;        memory[37245] <=  8'h66;        memory[37246] <=  8'h67;        memory[37247] <=  8'h73;        memory[37248] <=  8'h68;        memory[37249] <=  8'h64;        memory[37250] <=  8'h66;        memory[37251] <=  8'h68;        memory[37252] <=  8'h64;        memory[37253] <=  8'h6a;        memory[37254] <=  8'h68;        memory[37255] <=  8'h62;        memory[37256] <=  8'h67;        memory[37257] <=  8'h63;        memory[37258] <=  8'h61;        memory[37259] <=  8'h66;        memory[37260] <=  8'h73;        memory[37261] <=  8'h79;        memory[37262] <=  8'h67;        memory[37263] <=  8'h6b;        memory[37264] <=  8'h75;        memory[37265] <=  8'h64;        memory[37266] <=  8'h68;        memory[37267] <=  8'h62;        memory[37268] <=  8'h77;        memory[37269] <=  8'h76;        memory[37270] <=  8'h67;        memory[37271] <=  8'h61;        memory[37272] <=  8'h66;        memory[37273] <=  8'h64;        memory[37274] <=  8'h74;        memory[37275] <=  8'h75;        memory[37276] <=  8'h66;        memory[37277] <=  8'h79;        memory[37278] <=  8'h67;        memory[37279] <=  8'h69;        memory[37280] <=  8'h75;        memory[37281] <=  8'h68;        memory[37282] <=  8'h6c;        memory[37283] <=  8'h6a;        memory[37284] <=  8'h62;        memory[37285] <=  8'h6b;        memory[37286] <=  8'h68;        memory[37287] <=  8'h76;        memory[37288] <=  8'h67;        memory[37289] <=  8'h63;        memory[37290] <=  8'h66;        memory[37291] <=  8'h78;        memory[37292] <=  8'h64;        memory[37293] <=  8'h74;        memory[37294] <=  8'h75;        memory[37295] <=  8'h79;        memory[37296] <=  8'h69;        memory[37297] <=  8'h75;        memory[37298] <=  8'h68;        memory[37299] <=  8'h6c;        memory[37300] <=  8'h6a;        memory[37301] <=  8'h6b;        memory[37302] <=  8'h67;        memory[37303] <=  8'h6a;        memory[37304] <=  8'h63;        memory[37305] <=  8'h66;        memory[37306] <=  8'h68;        memory[37307] <=  8'h64;        memory[37308] <=  8'h67;        memory[37309] <=  8'h72;        memory[37310] <=  8'h79;        memory[37311] <=  8'h74;        memory[37312] <=  8'h66;        memory[37313] <=  8'h75;        memory[37314] <=  8'h79;        memory[37315] <=  8'h69;        memory[37316] <=  8'h68;        memory[37317] <=  8'h6c;        memory[37318] <=  8'h62;        memory[37319] <=  8'h6d;        memory[37320] <=  8'h76;        memory[37321] <=  8'h6e;        memory[37322] <=  8'h63;        memory[37323] <=  8'h66;        memory[37324] <=  8'h68;        memory[37325] <=  8'h64;        memory[37326] <=  8'h74;        memory[37327] <=  8'h75;        memory[37328] <=  8'h67;        memory[37329] <=  8'h79;        memory[37330] <=  8'h69;        memory[37331] <=  8'h68;        memory[37332] <=  8'h75;        memory[37333] <=  8'h6a;        memory[37334] <=  8'h6c;        memory[37335] <=  8'h62;        memory[37336] <=  8'h6d;        memory[37337] <=  8'h76;        memory[37338] <=  8'h6e;        memory[37339] <=  8'h63;        memory[37340] <=  8'h66;        memory[37341] <=  8'h68;        memory[37342] <=  8'h67;        memory[37343] <=  8'h79;        memory[37344] <=  8'h68;        memory[37345] <=  8'h75;        memory[37346] <=  8'h6a;        memory[37347] <=  8'h6e;        memory[37348] <=  8'h2c;        memory[37349] <=  8'h62;        memory[37350] <=  8'h6e;        memory[37351] <=  8'h6d;        memory[37352] <=  8'h76;        memory[37353] <=  8'h6e;        memory[37354] <=  8'h63;        memory[37355] <=  8'h66;        memory[37356] <=  8'h68;        memory[37357] <=  8'h74;        memory[37358] <=  8'h79;        memory[37359] <=  8'h69;        memory[37360] <=  8'h75;        memory[37361] <=  8'h6c;        memory[37362] <=  8'h6a;        memory[37363] <=  8'h62;        memory[37364] <=  8'h6d;        memory[37365] <=  8'h76;        memory[37366] <=  8'h6e;        memory[37367] <=  8'h63;        memory[37368] <=  8'h66;        memory[37369] <=  8'h74;        memory[37370] <=  8'h75;        memory[37371] <=  8'h79;        memory[37372] <=  8'h69;        memory[37373] <=  8'h68;        memory[37374] <=  8'h6b;        memory[37375] <=  8'h62;        memory[37376] <=  8'h76;        memory[37377] <=  8'h63;        memory[37378] <=  8'h66;        memory[37379] <=  8'h67;        memory[37380] <=  8'h74;        memory[37381] <=  8'h75;        memory[37382] <=  8'h79;        memory[37383] <=  8'h69;        memory[37384] <=  8'h75;        memory[37385] <=  8'h68;        memory[37386] <=  8'h6a;        memory[37387] <=  8'h6b;        memory[37388] <=  8'h62;        memory[37389] <=  8'h76;        memory[37390] <=  8'h63;        memory[37391] <=  8'h66;        memory[37392] <=  8'h74;        memory[37393] <=  8'h75;        memory[37394] <=  8'h79;        memory[37395] <=  8'h69;        memory[37396] <=  8'h75;        memory[37397] <=  8'h6a;        memory[37398] <=  8'h6b;        memory[37399] <=  8'h6e;        memory[37400] <=  8'h62;        memory[37401] <=  8'h76;        memory[37402] <=  8'h67;        memory[37403] <=  8'h66;        memory[37404] <=  8'h74;        memory[37405] <=  8'h79;        memory[37406] <=  8'h75;        memory[37407] <=  8'h75;        memory[37408] <=  8'h69;        memory[37409] <=  8'h6a;        memory[37410] <=  8'h6b;        memory[37411] <=  8'h68;        memory[37412] <=  8'h62;        memory[37413] <=  8'h6a;        memory[37414] <=  8'h67;        memory[37415] <=  8'h68;        memory[37416] <=  8'h66;        memory[37417] <=  8'h79;        memory[37418] <=  8'h74;        memory[37419] <=  8'h79;        memory[37420] <=  8'h69;        memory[37421] <=  8'h75;        memory[37422] <=  8'h64;        memory[37423] <=  8'h6a;        memory[37424] <=  8'h6b;        memory[37425] <=  8'h68;        memory[37426] <=  8'h63;        memory[37427] <=  8'h7a;        memory[37428] <=  8'h67;        memory[37429] <=  8'h68;        memory[37430] <=  8'h74;        memory[37431] <=  8'h75;        memory[37432] <=  8'h79;        memory[37433] <=  8'h69;        memory[37434] <=  8'h61;        memory[37435] <=  8'h73;        memory[37436] <=  8'h75;        memory[37437] <=  8'h6a;        memory[37438] <=  8'h6b;        memory[37439] <=  8'h62;        memory[37440] <=  8'h6e;        memory[37441] <=  8'h61;        memory[37442] <=  8'h76;        memory[37443] <=  8'h63;        memory[37444] <=  8'h66;        memory[37445] <=  8'h68;        memory[37446] <=  8'h75;        memory[37447] <=  8'h61;        memory[37448] <=  8'h73;        memory[37449] <=  8'h79;        memory[37450] <=  8'h64;        memory[37451] <=  8'h75;        memory[37452] <=  8'h69;        memory[37453] <=  8'h6a;        memory[37454] <=  8'h61;        memory[37455] <=  8'h6b;        memory[37456] <=  8'h62;        memory[37457] <=  8'h63;        memory[37458] <=  8'h78;        memory[37459] <=  8'h68;        memory[37460] <=  8'h67;        memory[37461] <=  8'h79;        memory[37462] <=  8'h75;        memory[37463] <=  8'h7a;        memory[37464] <=  8'h63;        memory[37465] <=  8'h61;        memory[37466] <=  8'h73;        memory[37467] <=  8'h69;        memory[37468] <=  8'h75;        memory[37469] <=  8'h6f;        memory[37470] <=  8'h69;        memory[37471] <=  8'h6a;        memory[37472] <=  8'h61;        memory[37473] <=  8'h6c;        memory[37474] <=  8'h63;        memory[37475] <=  8'h78;        memory[37476] <=  8'h62;        memory[37477] <=  8'h63;        memory[37478] <=  8'h20;        memory[37479] <=  8'h6e;        memory[37480] <=  8'h76;        memory[37481] <=  8'h63;        memory[37482] <=  8'h61;        memory[37483] <=  8'h64;        memory[37484] <=  8'h73;        memory[37485] <=  8'h67;        memory[37486] <=  8'h79;        memory[37487] <=  8'h68;        memory[37488] <=  8'h75;        memory[37489] <=  8'h61;        memory[37490] <=  8'h6a;        memory[37491] <=  8'h6b;        memory[37492] <=  8'h78;        memory[37493] <=  8'h62;        memory[37494] <=  8'h20;        memory[37495] <=  8'h6e;        memory[37496] <=  8'h76;        memory[37497] <=  8'h63;        memory[37498] <=  8'h61;        memory[37499] <=  8'h73;        memory[37500] <=  8'h67;        memory[37501] <=  8'h68;        memory[37502] <=  8'h75;        memory[37503] <=  8'h6a;        memory[37504] <=  8'h6c;        memory[37505] <=  8'h6b;        memory[37506] <=  8'h63;        memory[37507] <=  8'h78;        memory[37508] <=  8'h20;        memory[37509] <=  8'h6a;        memory[37510] <=  8'h6b;        memory[37511] <=  8'h68;        memory[37512] <=  8'h61;        memory[37513] <=  8'h73;        memory[37514] <=  8'h76;        memory[37515] <=  8'h64;        memory[37516] <=  8'h6e;        memory[37517] <=  8'h20;        memory[37518] <=  8'h62;        memory[37519] <=  8'h6e;        memory[37520] <=  8'h6d;        memory[37521] <=  8'h6b;        memory[37522] <=  8'h77;        memory[37523] <=  8'h64;        memory[37524] <=  8'h6f;        memory[37525] <=  8'h77;        memory[37526] <=  8'h69;        memory[37527] <=  8'h6f;        memory[37528] <=  8'h75;        memory[37529] <=  8'h69;        memory[37530] <=  8'h68;        memory[37531] <=  8'h62;        memory[37532] <=  8'h6e;        memory[37533] <=  8'h6b;        memory[37534] <=  8'h77;        memory[37535] <=  8'h69;        memory[37536] <=  8'h6f;        memory[37537] <=  8'h75;        memory[37538] <=  8'h71;        memory[37539] <=  8'h69;        memory[37540] <=  8'h79;        memory[37541] <=  8'h67;        memory[37542] <=  8'h6a;        memory[37543] <=  8'h64;        memory[37544] <=  8'h61;        memory[37545] <=  8'h76;        memory[37546] <=  8'h62;        memory[37547] <=  8'h6e;        memory[37548] <=  8'h6b;        memory[37549] <=  8'h6f;        memory[37550] <=  8'h70;        memory[37551] <=  8'h64;        memory[37552] <=  8'h76;        memory[37553] <=  8'h69;        memory[37554] <=  8'h6f;        memory[37555] <=  8'h75;        memory[37556] <=  8'h69;        memory[37557] <=  8'h48;        memory[37558] <=  8'h42;        memory[37559] <=  8'h6b;        memory[37560] <=  8'h64;        memory[37561] <=  8'h6e;        memory[37562] <=  8'h6c;        memory[37563] <=  8'h71;        memory[37564] <=  8'h6b;        memory[37565] <=  8'h6d;        memory[37566] <=  8'h6a;        memory[37567] <=  8'h70;        memory[37568] <=  8'h69;        memory[37569] <=  8'h6f;        memory[37570] <=  8'h68;        memory[37571] <=  8'h65;        memory[37572] <=  8'h66;        memory[37573] <=  8'h75;        memory[37574] <=  8'h67;        memory[37575] <=  8'h69;        memory[37576] <=  8'h73;        memory[37577] <=  8'h61;        memory[37578] <=  8'h62;        memory[37579] <=  8'h64;        memory[37580] <=  8'h6b;        memory[37581] <=  8'h6a;        memory[37582] <=  8'h6b;        memory[37583] <=  8'h6c;        memory[37584] <=  8'h6a;        memory[37585] <=  8'h69;        memory[37586] <=  8'h73;        memory[37587] <=  8'h6f;        memory[37588] <=  8'h71;        memory[37589] <=  8'h68;        memory[37590] <=  8'h77;        memory[37591] <=  8'h67;        memory[37592] <=  8'h69;        memory[37593] <=  8'h79;        memory[37594] <=  8'h6a;        memory[37595] <=  8'h64;        memory[37596] <=  8'h76;        memory[37597] <=  8'h62;        memory[37598] <=  8'h6e;        memory[37599] <=  8'h61;        memory[37600] <=  8'h73;        memory[37601] <=  8'h66;        memory[37602] <=  8'h6c;        memory[37603] <=  8'h6b;        memory[37604] <=  8'h64;        memory[37605] <=  8'h6a;        memory[37606] <=  8'h68;        memory[37607] <=  8'h63;        memory[37608] <=  8'h67;        memory[37609] <=  8'h6a;        memory[37610] <=  8'h76;        memory[37611] <=  8'h73;        memory[37612] <=  8'h64;        memory[37613] <=  8'h62;        memory[37614] <=  8'h62;        memory[37615] <=  8'h61;        memory[37616] <=  8'h72;        memory[37617] <=  8'h62;        memory[37618] <=  8'h62;        memory[37619] <=  8'h73;        memory[37620] <=  8'h62;        memory[37621] <=  8'h67;        memory[37622] <=  8'h73;        memory[37623] <=  8'h66;        memory[37624] <=  8'h67;        memory[37625] <=  8'h61;        memory[37626] <=  8'h68;        memory[37627] <=  8'h66;        memory[37628] <=  8'h73;        memory[37629] <=  8'h68;        memory[37630] <=  8'h61;        memory[37631] <=  8'h66;        memory[37632] <=  8'h73;        memory[37633] <=  8'h66;        memory[37634] <=  8'h68;        memory[37635] <=  8'h61;        memory[37636] <=  8'h69;        memory[37637] <=  8'h64;        memory[37638] <=  8'h75;        memory[37639] <=  8'h67;        memory[37640] <=  8'h64;        memory[37641] <=  8'h77;        memory[37642] <=  8'h62;        memory[37643] <=  8'h61;        memory[37644] <=  8'h62;        memory[37645] <=  8'h72;        memory[37646] <=  8'h62;        memory[37647] <=  8'h61;        memory[37648] <=  8'h62;        memory[37649] <=  8'h62;        memory[37650] <=  8'h74;        memory[37651] <=  8'h62;        memory[37652] <=  8'h62;        memory[37653] <=  8'h62;        memory[37654] <=  8'h62;        memory[37655] <=  8'h62;        memory[37656] <=  8'h62;        memory[37657] <=  8'h62;        memory[37658] <=  8'h62;        memory[37659] <=  8'h61;        memory[37660] <=  8'h62;        memory[37661] <=  8'h62;        memory[37662] <=  8'h72;        memory[37663] <=  8'h74;        memory[37664] <=  8'h62;        memory[37665] <=  8'h62;        memory[37666] <=  8'h61;        memory[37667] <=  8'h62;        memory[37668] <=  8'h72;        memory[37669] <=  8'h62;        memory[37670] <=  8'h74;        memory[37671] <=  8'h62;        memory[37672] <=  8'h62;        memory[37673] <=  8'h62;        memory[37674] <=  8'h63;        memory[37675] <=  8'h61;        memory[37676] <=  8'h72;        memory[37677] <=  8'h74;        memory[37678] <=  8'h73;        memory[37679] <=  8'h62;        memory[37680] <=  8'h61;        memory[37681] <=  8'h72;        memory[37682] <=  8'h74;        memory[37683] <=  8'h74;        memory[37684] <=  8'h62;        memory[37685] <=  8'h61;        memory[37686] <=  8'h72;        memory[37687] <=  8'h74;        memory[37688] <=  8'h78;        memory[37689] <=  8'h61;        memory[37690] <=  8'h74;        memory[37691] <=  8'h6b;        memory[37692] <=  8'h73;        memory[37693] <=  8'h68;        memory[37694] <=  8'h63;        memory[37695] <=  8'h66;        memory[37696] <=  8'h69;        memory[37697] <=  8'h77;        memory[37698] <=  8'h68;        memory[37699] <=  8'h61;        memory[37700] <=  8'h74;        memory[37701] <=  8'h61;        memory[37702] <=  8'h6e;        memory[37703] <=  8'h61;        memory[37704] <=  8'h62;        memory[37705] <=  8'h61;        memory[37706] <=  8'h63;        memory[37707] <=  8'h61;        memory[37708] <=  8'h74;        memory[37709] <=  8'h61;        memory[37710] <=  8'h62;        memory[37711] <=  8'h61;        memory[37712] <=  8'h72;        memory[37713] <=  8'h63;        memory[37714] <=  8'h61;        memory[37715] <=  8'h68;        memory[37716] <=  8'h64;        memory[37717] <=  8'h75;        memory[37718] <=  8'h63;        memory[37719] <=  8'h74;        memory[37720] <=  8'h61;        memory[37721] <=  8'h64;        memory[37722] <=  8'h61;        memory[37723] <=  8'h61;        memory[37724] <=  8'h63;        memory[37725] <=  8'h61;        memory[37726] <=  8'h72;        memory[37727] <=  8'h63;        memory[37728] <=  8'h74;        memory[37729] <=  8'h72;        memory[37730] <=  8'h63;        memory[37731] <=  8'h61;        memory[37732] <=  8'h74;        memory[37733] <=  8'h72;        memory[37734] <=  8'h63;        memory[37735] <=  8'h61;        memory[37736] <=  8'h74;        memory[37737] <=  8'h63;        memory[37738] <=  8'h62;        memory[37739] <=  8'h61;        memory[37740] <=  8'h74;        memory[37741] <=  8'h62;        memory[37742] <=  8'h72;        memory[37743] <=  8'h63;        memory[37744] <=  8'h61;        memory[37745] <=  8'h74;        memory[37746] <=  8'h72;        memory[37747] <=  8'h6e;        memory[37748] <=  8'h62;        memory[37749] <=  8'h61;        memory[37750] <=  8'h63;        memory[37751] <=  8'h61;        memory[37752] <=  8'h74;        memory[37753] <=  8'h79;        memory[37754] <=  8'h73;        memory[37755] <=  8'h6e;        memory[37756] <=  8'h63;        memory[37757] <=  8'h74;        memory[37758] <=  8'h61;        memory[37759] <=  8'h6e;        memory[37760] <=  8'h62;        memory[37761] <=  8'h61;        memory[37762] <=  8'h63;        memory[37763] <=  8'h72;        memory[37764] <=  8'h6e;        memory[37765] <=  8'h74;        memory[37766] <=  8'h61;        memory[37767] <=  8'h62;        memory[37768] <=  8'h74;        memory[37769] <=  8'h6e;        memory[37770] <=  8'h61;        memory[37771] <=  8'h72;        memory[37772] <=  8'h62;        memory[37773] <=  8'h78;        memory[37774] <=  8'h74;        memory[37775] <=  8'h61;        memory[37776] <=  8'h72;        memory[37777] <=  8'h62;        memory[37778] <=  8'h61;        memory[37779] <=  8'h72;        memory[37780] <=  8'h74;        memory[37781] <=  8'h74;        memory[37782] <=  8'h62;        memory[37783] <=  8'h61;        memory[37784] <=  8'h72;        memory[37785] <=  8'h74;        memory[37786] <=  8'h78;        memory[37787] <=  8'h61;        memory[37788] <=  8'h74;        memory[37789] <=  8'h6b;        memory[37790] <=  8'h73;        memory[37791] <=  8'h68;        memory[37792] <=  8'h63;        memory[37793] <=  8'h66;        memory[37794] <=  8'h69;        memory[37795] <=  8'h77;        memory[37796] <=  8'h68;        memory[37797] <=  8'h61;        memory[37798] <=  8'h74;        memory[37799] <=  8'h61;        memory[37800] <=  8'h6e;        memory[37801] <=  8'h61;        memory[37802] <=  8'h62;        memory[37803] <=  8'h61;        memory[37804] <=  8'h63;        memory[37805] <=  8'h61;        memory[37806] <=  8'h74;        memory[37807] <=  8'h61;        memory[37808] <=  8'h62;        memory[37809] <=  8'h61;        memory[37810] <=  8'h72;        memory[37811] <=  8'h63;        memory[37812] <=  8'h61;        memory[37813] <=  8'h68;        memory[37814] <=  8'h64;        memory[37815] <=  8'h75;        memory[37816] <=  8'h63;        memory[37817] <=  8'h74;        memory[37818] <=  8'h61;        memory[37819] <=  8'h64;        memory[37820] <=  8'h61;        memory[37821] <=  8'h61;        memory[37822] <=  8'h63;        memory[37823] <=  8'h61;        memory[37824] <=  8'h72;        memory[37825] <=  8'h63;        memory[37826] <=  8'h74;        memory[37827] <=  8'h72;        memory[37828] <=  8'h63;        memory[37829] <=  8'h61;        memory[37830] <=  8'h74;        memory[37831] <=  8'h72;        memory[37832] <=  8'h63;        memory[37833] <=  8'h61;        memory[37834] <=  8'h74;        memory[37835] <=  8'h63;        memory[37836] <=  8'h62;        memory[37837] <=  8'h61;        memory[37838] <=  8'h74;        memory[37839] <=  8'h62;        memory[37840] <=  8'h72;        memory[37841] <=  8'h63;        memory[37842] <=  8'h61;        memory[37843] <=  8'h74;        memory[37844] <=  8'h72;        memory[37845] <=  8'h6e;        memory[37846] <=  8'h62;        memory[37847] <=  8'h61;        memory[37848] <=  8'h63;        memory[37849] <=  8'h61;        memory[37850] <=  8'h74;        memory[37851] <=  8'h79;        memory[37852] <=  8'h73;        memory[37853] <=  8'h6e;        memory[37854] <=  8'h63;        memory[37855] <=  8'h74;        memory[37856] <=  8'h61;        memory[37857] <=  8'h6e;        memory[37858] <=  8'h62;        memory[37859] <=  8'h61;        memory[37860] <=  8'h63;        memory[37861] <=  8'h72;        memory[37862] <=  8'h6e;        memory[37863] <=  8'h74;        memory[37864] <=  8'h61;        memory[37865] <=  8'h62;        memory[37866] <=  8'h74;        memory[37867] <=  8'h6e;        memory[37868] <=  8'h61;        memory[37869] <=  8'h72;        memory[37870] <=  8'h62;        memory[37871] <=  8'h78;        memory[37872] <=  8'h74;        memory[37873] <=  8'h61;        memory[37874] <=  8'h72;        memory[37875] <=  8'h62;        memory[37876] <=  8'h61;        memory[37877] <=  8'h72;        memory[37878] <=  8'h74;        memory[37879] <=  8'h74;        memory[37880] <=  8'h62;        memory[37881] <=  8'h61;        memory[37882] <=  8'h72;        memory[37883] <=  8'h74;        memory[37884] <=  8'h78;        memory[37885] <=  8'h61;        memory[37886] <=  8'h74;        memory[37887] <=  8'h6b;        memory[37888] <=  8'h73;        memory[37889] <=  8'h68;        memory[37890] <=  8'h63;        memory[37891] <=  8'h66;        memory[37892] <=  8'h69;        memory[37893] <=  8'h77;        memory[37894] <=  8'h68;        memory[37895] <=  8'h61;        memory[37896] <=  8'h74;        memory[37897] <=  8'h61;        memory[37898] <=  8'h6e;        memory[37899] <=  8'h61;        memory[37900] <=  8'h62;        memory[37901] <=  8'h61;        memory[37902] <=  8'h63;        memory[37903] <=  8'h61;        memory[37904] <=  8'h74;        memory[37905] <=  8'h61;        memory[37906] <=  8'h62;        memory[37907] <=  8'h61;        memory[37908] <=  8'h72;        memory[37909] <=  8'h63;        memory[37910] <=  8'h61;        memory[37911] <=  8'h68;        memory[37912] <=  8'h64;        memory[37913] <=  8'h75;        memory[37914] <=  8'h63;        memory[37915] <=  8'h74;        memory[37916] <=  8'h61;        memory[37917] <=  8'h64;        memory[37918] <=  8'h61;        memory[37919] <=  8'h61;        memory[37920] <=  8'h63;        memory[37921] <=  8'h61;        memory[37922] <=  8'h72;        memory[37923] <=  8'h63;        memory[37924] <=  8'h74;        memory[37925] <=  8'h72;        memory[37926] <=  8'h63;        memory[37927] <=  8'h61;        memory[37928] <=  8'h74;        memory[37929] <=  8'h72;        memory[37930] <=  8'h63;        memory[37931] <=  8'h61;        memory[37932] <=  8'h74;        memory[37933] <=  8'h63;        memory[37934] <=  8'h62;        memory[37935] <=  8'h61;        memory[37936] <=  8'h74;        memory[37937] <=  8'h62;        memory[37938] <=  8'h72;        memory[37939] <=  8'h63;        memory[37940] <=  8'h61;        memory[37941] <=  8'h74;        memory[37942] <=  8'h72;        memory[37943] <=  8'h6e;        memory[37944] <=  8'h62;        memory[37945] <=  8'h61;        memory[37946] <=  8'h63;        memory[37947] <=  8'h61;        memory[37948] <=  8'h74;        memory[37949] <=  8'h79;        memory[37950] <=  8'h73;        memory[37951] <=  8'h6e;        memory[37952] <=  8'h63;        memory[37953] <=  8'h74;        memory[37954] <=  8'h61;        memory[37955] <=  8'h6e;        memory[37956] <=  8'h62;        memory[37957] <=  8'h61;        memory[37958] <=  8'h63;        memory[37959] <=  8'h72;        memory[37960] <=  8'h6e;        memory[37961] <=  8'h74;        memory[37962] <=  8'h61;        memory[37963] <=  8'h62;        memory[37964] <=  8'h74;        memory[37965] <=  8'h6e;        memory[37966] <=  8'h61;        memory[37967] <=  8'h72;        memory[37968] <=  8'h62;        memory[37969] <=  8'h78;        memory[37970] <=  8'h74;        memory[37971] <=  8'h61;        memory[37972] <=  8'h72;        memory[37973] <=  8'h5d;        memory[37974] <=  8'h5d;        memory[37975] <=  8'h65;        memory[37976] <=  8'h66;        memory[37977] <=  8'h77;        memory[37978] <=  8'h65;        memory[37979] <=  8'h5d;        memory[37980] <=  8'h65;        memory[37981] <=  8'h67;        memory[37982] <=  8'h73;        memory[37983] <=  8'h67;        memory[37984] <=  8'h66;        memory[37985] <=  8'h62;        memory[37986] <=  8'h61;        memory[37987] <=  8'h72;        memory[37988] <=  8'h74;        memory[37989] <=  8'h74;        memory[37990] <=  8'h62;        memory[37991] <=  8'h61;        memory[37992] <=  8'h72;        memory[37993] <=  8'h74;        memory[37994] <=  8'h78;        memory[37995] <=  8'h61;        memory[37996] <=  8'h74;        memory[37997] <=  8'h6b;        memory[37998] <=  8'h73;        memory[37999] <=  8'h68;        memory[38000] <=  8'h63;        memory[38001] <=  8'h66;        memory[38002] <=  8'h69;        memory[38003] <=  8'h77;        memory[38004] <=  8'h68;        memory[38005] <=  8'h61;        memory[38006] <=  8'h74;        memory[38007] <=  8'h61;        memory[38008] <=  8'h6e;        memory[38009] <=  8'h61;        memory[38010] <=  8'h62;        memory[38011] <=  8'h61;        memory[38012] <=  8'h63;        memory[38013] <=  8'h61;        memory[38014] <=  8'h74;        memory[38015] <=  8'h61;        memory[38016] <=  8'h62;        memory[38017] <=  8'h61;        memory[38018] <=  8'h72;        memory[38019] <=  8'h63;        memory[38020] <=  8'h61;        memory[38021] <=  8'h68;        memory[38022] <=  8'h64;        memory[38023] <=  8'h75;        memory[38024] <=  8'h63;        memory[38025] <=  8'h74;        memory[38026] <=  8'h61;        memory[38027] <=  8'h64;        memory[38028] <=  8'h61;        memory[38029] <=  8'h61;        memory[38030] <=  8'h63;        memory[38031] <=  8'h61;        memory[38032] <=  8'h72;        memory[38033] <=  8'h63;        memory[38034] <=  8'h74;        memory[38035] <=  8'h72;        memory[38036] <=  8'h63;        memory[38037] <=  8'h61;        memory[38038] <=  8'h74;        memory[38039] <=  8'h72;        memory[38040] <=  8'h63;        memory[38041] <=  8'h61;        memory[38042] <=  8'h74;        memory[38043] <=  8'h63;        memory[38044] <=  8'h62;        memory[38045] <=  8'h61;        memory[38046] <=  8'h74;        memory[38047] <=  8'h62;        memory[38048] <=  8'h72;        memory[38049] <=  8'h63;        memory[38050] <=  8'h61;        memory[38051] <=  8'h74;        memory[38052] <=  8'h72;        memory[38053] <=  8'h6e;        memory[38054] <=  8'h62;        memory[38055] <=  8'h61;        memory[38056] <=  8'h63;        memory[38057] <=  8'h61;        memory[38058] <=  8'h74;        memory[38059] <=  8'h79;        memory[38060] <=  8'h73;        memory[38061] <=  8'h6e;        memory[38062] <=  8'h63;        memory[38063] <=  8'h74;        memory[38064] <=  8'h61;        memory[38065] <=  8'h6e;        memory[38066] <=  8'h62;        memory[38067] <=  8'h61;        memory[38068] <=  8'h63;        memory[38069] <=  8'h72;        memory[38070] <=  8'h6e;        memory[38071] <=  8'h74;        memory[38072] <=  8'h61;        memory[38073] <=  8'h62;        memory[38074] <=  8'h74;        memory[38075] <=  8'h6e;        memory[38076] <=  8'h61;        memory[38077] <=  8'h72;        memory[38078] <=  8'h62;        memory[38079] <=  8'h78;        memory[38080] <=  8'h74;        memory[38081] <=  8'h61;        memory[38082] <=  8'h72;        memory[38083] <=  8'h62;        memory[38084] <=  8'h61;        memory[38085] <=  8'h72;        memory[38086] <=  8'h74;        memory[38087] <=  8'h74;        memory[38088] <=  8'h62;        memory[38089] <=  8'h61;        memory[38090] <=  8'h72;        memory[38091] <=  8'h74;        memory[38092] <=  8'h78;        memory[38093] <=  8'h61;        memory[38094] <=  8'h74;        memory[38095] <=  8'h6b;        memory[38096] <=  8'h73;        memory[38097] <=  8'h68;        memory[38098] <=  8'h63;        memory[38099] <=  8'h66;        memory[38100] <=  8'h69;        memory[38101] <=  8'h77;        memory[38102] <=  8'h68;        memory[38103] <=  8'h61;        memory[38104] <=  8'h74;        memory[38105] <=  8'h61;        memory[38106] <=  8'h6e;        memory[38107] <=  8'h61;        memory[38108] <=  8'h62;        memory[38109] <=  8'h61;        memory[38110] <=  8'h63;        memory[38111] <=  8'h61;        memory[38112] <=  8'h74;        memory[38113] <=  8'h61;        memory[38114] <=  8'h62;        memory[38115] <=  8'h61;        memory[38116] <=  8'h72;        memory[38117] <=  8'h63;        memory[38118] <=  8'h61;        memory[38119] <=  8'h68;        memory[38120] <=  8'h64;        memory[38121] <=  8'h75;        memory[38122] <=  8'h63;        memory[38123] <=  8'h74;        memory[38124] <=  8'h61;        memory[38125] <=  8'h64;        memory[38126] <=  8'h61;        memory[38127] <=  8'h61;        memory[38128] <=  8'h63;        memory[38129] <=  8'h61;        memory[38130] <=  8'h72;        memory[38131] <=  8'h63;        memory[38132] <=  8'h74;        memory[38133] <=  8'h72;        memory[38134] <=  8'h63;        memory[38135] <=  8'h61;        memory[38136] <=  8'h74;        memory[38137] <=  8'h72;        memory[38138] <=  8'h63;        memory[38139] <=  8'h61;        memory[38140] <=  8'h74;        memory[38141] <=  8'h63;        memory[38142] <=  8'h62;        memory[38143] <=  8'h61;        memory[38144] <=  8'h74;        memory[38145] <=  8'h62;        memory[38146] <=  8'h72;        memory[38147] <=  8'h63;        memory[38148] <=  8'h61;        memory[38149] <=  8'h74;        memory[38150] <=  8'h72;        memory[38151] <=  8'h6e;        memory[38152] <=  8'h62;        memory[38153] <=  8'h61;        memory[38154] <=  8'h63;        memory[38155] <=  8'h61;        memory[38156] <=  8'h74;        memory[38157] <=  8'h79;        memory[38158] <=  8'h73;        memory[38159] <=  8'h6e;        memory[38160] <=  8'h63;        memory[38161] <=  8'h74;        memory[38162] <=  8'h61;        memory[38163] <=  8'h6e;        memory[38164] <=  8'h62;        memory[38165] <=  8'h61;        memory[38166] <=  8'h63;        memory[38167] <=  8'h72;        memory[38168] <=  8'h6e;        memory[38169] <=  8'h74;        memory[38170] <=  8'h61;        memory[38171] <=  8'h62;        memory[38172] <=  8'h74;        memory[38173] <=  8'h6e;        memory[38174] <=  8'h61;        memory[38175] <=  8'h72;        memory[38176] <=  8'h62;        memory[38177] <=  8'h78;        memory[38178] <=  8'h74;        memory[38179] <=  8'h61;        memory[38180] <=  8'h72;        memory[38181] <=  8'h64;        memory[38182] <=  8'h66;        memory[38183] <=  8'h73;        memory[38184] <=  8'h67;        memory[38185] <=  8'h76;        memory[38186] <=  8'h68;        memory[38187] <=  8'h62;        memory[38188] <=  8'h6b;        memory[38189] <=  8'h6a;        memory[38190] <=  8'h6e;        memory[38191] <=  8'h6d;        memory[38192] <=  8'h62;        memory[38193] <=  8'h76;        memory[38194] <=  8'h78;        memory[38195] <=  8'h63;        memory[38196] <=  8'h73;        memory[38197] <=  8'h66;        memory[38198] <=  8'h72;        memory[38199] <=  8'h74;        memory[38200] <=  8'h79;        memory[38201] <=  8'h75;        memory[38202] <=  8'h6a;        memory[38203] <=  8'h6e;        memory[38204] <=  8'h62;        memory[38205] <=  8'h76;        memory[38206] <=  8'h63;        memory[38207] <=  8'h64;        memory[38208] <=  8'h74;        memory[38209] <=  8'h79;        memory[38210] <=  8'h75;        memory[38211] <=  8'h69;        memory[38212] <=  8'h6b;        memory[38213] <=  8'h6d;        memory[38214] <=  8'h6e;        memory[38215] <=  8'h62;        memory[38216] <=  8'h76;        memory[38217] <=  8'h63;        memory[38218] <=  8'h78;        memory[38219] <=  8'h73;        memory[38220] <=  8'h64;        memory[38221] <=  8'h72;        memory[38222] <=  8'h74;        memory[38223] <=  8'h79;        memory[38224] <=  8'h75;        memory[38225] <=  8'h69;        memory[38226] <=  8'h6b;        memory[38227] <=  8'h6d;        memory[38228] <=  8'h6e;        memory[38229] <=  8'h62;        memory[38230] <=  8'h76;        memory[38231] <=  8'h63;        memory[38232] <=  8'h73;        memory[38233] <=  8'h77;        memory[38234] <=  8'h33;        memory[38235] <=  8'h34;        memory[38236] <=  8'h35;        memory[38237] <=  8'h36;        memory[38238] <=  8'h37;        memory[38239] <=  8'h38;        memory[38240] <=  8'h69;        memory[38241] <=  8'h6b;        memory[38242] <=  8'h6d;        memory[38243] <=  8'h6e;        memory[38244] <=  8'h62;        memory[38245] <=  8'h76;        memory[38246] <=  8'h63;        memory[38247] <=  8'h64;        memory[38248] <=  8'h65;        memory[38249] <=  8'h72;        memory[38250] <=  8'h36;        memory[38251] <=  8'h37;        memory[38252] <=  8'h38;        memory[38253] <=  8'h69;        memory[38254] <=  8'h6f;        memory[38255] <=  8'h6b;        memory[38256] <=  8'h6a;        memory[38257] <=  8'h6e;        memory[38258] <=  8'h62;        memory[38259] <=  8'h76;        memory[38260] <=  8'h63;        memory[38261] <=  8'h64;        memory[38262] <=  8'h72;        memory[38263] <=  8'h74;        memory[38264] <=  8'h79;        memory[38265] <=  8'h75;        memory[38266] <=  8'h73;        memory[38267] <=  8'h6a;        memory[38268] <=  8'h63;        memory[38269] <=  8'h6e;        memory[38270] <=  8'h62;        memory[38271] <=  8'h64;        memory[38272] <=  8'h66;        memory[38273] <=  8'h73;        memory[38274] <=  8'h74;        memory[38275] <=  8'h79;        memory[38276] <=  8'h75;        memory[38277] <=  8'h61;        memory[38278] <=  8'h69;        memory[38279] <=  8'h6b;        memory[38280] <=  8'h78;        memory[38281] <=  8'h6d;        memory[38282] <=  8'h6e;        memory[38283] <=  8'h73;        memory[38284] <=  8'h6a;        memory[38285] <=  8'h6f;        memory[38286] <=  8'h64;        memory[38287] <=  8'h6c;        memory[38288] <=  8'h63;        memory[38289] <=  8'h78;        memory[38290] <=  8'h62;        memory[38291] <=  8'h61;        memory[38292] <=  8'h72;        memory[38293] <=  8'h74;        memory[38294] <=  8'h78;        memory[38295] <=  8'h61;        memory[38296] <=  8'h74;        memory[38297] <=  8'h6b;        memory[38298] <=  8'h73;        memory[38299] <=  8'h68;        memory[38300] <=  8'h63;        memory[38301] <=  8'h66;        memory[38302] <=  8'h69;        memory[38303] <=  8'h77;        memory[38304] <=  8'h68;        memory[38305] <=  8'h61;        memory[38306] <=  8'h74;        memory[38307] <=  8'h61;        memory[38308] <=  8'h6e;        memory[38309] <=  8'h61;        memory[38310] <=  8'h62;        memory[38311] <=  8'h61;        memory[38312] <=  8'h63;        memory[38313] <=  8'h61;        memory[38314] <=  8'h74;        memory[38315] <=  8'h61;        memory[38316] <=  8'h62;        memory[38317] <=  8'h61;        memory[38318] <=  8'h72;        memory[38319] <=  8'h63;        memory[38320] <=  8'h61;        memory[38321] <=  8'h68;        memory[38322] <=  8'h64;        memory[38323] <=  8'h75;        memory[38324] <=  8'h63;        memory[38325] <=  8'h74;        memory[38326] <=  8'h61;        memory[38327] <=  8'h64;        memory[38328] <=  8'h61;        memory[38329] <=  8'h61;        memory[38330] <=  8'h63;        memory[38331] <=  8'h61;        memory[38332] <=  8'h72;        memory[38333] <=  8'h62;        memory[38334] <=  8'h61;        memory[38335] <=  8'h72;        memory[38336] <=  8'h74;        memory[38337] <=  8'h78;        memory[38338] <=  8'h61;        memory[38339] <=  8'h74;        memory[38340] <=  8'h6b;        memory[38341] <=  8'h73;        memory[38342] <=  8'h68;        memory[38343] <=  8'h63;        memory[38344] <=  8'h66;        memory[38345] <=  8'h69;        memory[38346] <=  8'h77;        memory[38347] <=  8'h68;        memory[38348] <=  8'h61;        memory[38349] <=  8'h74;        memory[38350] <=  8'h61;        memory[38351] <=  8'h6e;        memory[38352] <=  8'h61;        memory[38353] <=  8'h62;        memory[38354] <=  8'h61;        memory[38355] <=  8'h63;        memory[38356] <=  8'h61;        memory[38357] <=  8'h74;        memory[38358] <=  8'h61;        memory[38359] <=  8'h62;        memory[38360] <=  8'h61;        memory[38361] <=  8'h72;        memory[38362] <=  8'h63;        memory[38363] <=  8'h61;        memory[38364] <=  8'h68;        memory[38365] <=  8'h64;        memory[38366] <=  8'h75;        memory[38367] <=  8'h63;        memory[38368] <=  8'h74;        memory[38369] <=  8'h61;        memory[38370] <=  8'h64;        memory[38371] <=  8'h61;        memory[38372] <=  8'h61;        memory[38373] <=  8'h63;        memory[38374] <=  8'h61;        memory[38375] <=  8'h72;        memory[38376] <=  8'h62;        memory[38377] <=  8'h61;        memory[38378] <=  8'h72;        memory[38379] <=  8'h74;        memory[38380] <=  8'h78;        memory[38381] <=  8'h61;        memory[38382] <=  8'h74;        memory[38383] <=  8'h6b;        memory[38384] <=  8'h73;        memory[38385] <=  8'h68;        memory[38386] <=  8'h63;        memory[38387] <=  8'h66;        memory[38388] <=  8'h69;        memory[38389] <=  8'h77;        memory[38390] <=  8'h68;        memory[38391] <=  8'h61;        memory[38392] <=  8'h74;        memory[38393] <=  8'h61;        memory[38394] <=  8'h6e;        memory[38395] <=  8'h61;        memory[38396] <=  8'h62;        memory[38397] <=  8'h61;        memory[38398] <=  8'h63;        memory[38399] <=  8'h61;        memory[38400] <=  8'h74;        memory[38401] <=  8'h61;        memory[38402] <=  8'h62;        memory[38403] <=  8'h61;        memory[38404] <=  8'h72;        memory[38405] <=  8'h63;        memory[38406] <=  8'h61;        memory[38407] <=  8'h68;        memory[38408] <=  8'h64;        memory[38409] <=  8'h75;        memory[38410] <=  8'h63;        memory[38411] <=  8'h74;        memory[38412] <=  8'h61;        memory[38413] <=  8'h64;        memory[38414] <=  8'h61;        memory[38415] <=  8'h61;        memory[38416] <=  8'h63;        memory[38417] <=  8'h61;        memory[38418] <=  8'h72;        memory[38419] <=  8'h62;        memory[38420] <=  8'h61;        memory[38421] <=  8'h72;        memory[38422] <=  8'h74;        memory[38423] <=  8'h78;        memory[38424] <=  8'h61;        memory[38425] <=  8'h74;        memory[38426] <=  8'h6b;        memory[38427] <=  8'h73;        memory[38428] <=  8'h68;        memory[38429] <=  8'h63;        memory[38430] <=  8'h66;        memory[38431] <=  8'h69;        memory[38432] <=  8'h77;        memory[38433] <=  8'h68;        memory[38434] <=  8'h61;        memory[38435] <=  8'h74;        memory[38436] <=  8'h61;        memory[38437] <=  8'h6e;        memory[38438] <=  8'h61;        memory[38439] <=  8'h62;        memory[38440] <=  8'h61;        memory[38441] <=  8'h63;        memory[38442] <=  8'h61;        memory[38443] <=  8'h74;        memory[38444] <=  8'h61;        memory[38445] <=  8'h62;        memory[38446] <=  8'h61;        memory[38447] <=  8'h72;        memory[38448] <=  8'h63;        memory[38449] <=  8'h61;        memory[38450] <=  8'h68;        memory[38451] <=  8'h64;        memory[38452] <=  8'h75;        memory[38453] <=  8'h63;        memory[38454] <=  8'h74;        memory[38455] <=  8'h61;        memory[38456] <=  8'h64;        memory[38457] <=  8'h61;        memory[38458] <=  8'h61;        memory[38459] <=  8'h63;        memory[38460] <=  8'h61;        memory[38461] <=  8'h72;        memory[38462] <=  8'h62;        memory[38463] <=  8'h61;        memory[38464] <=  8'h72;        memory[38465] <=  8'h74;        memory[38466] <=  8'h78;        memory[38467] <=  8'h61;        memory[38468] <=  8'h74;        memory[38469] <=  8'h6b;        memory[38470] <=  8'h73;        memory[38471] <=  8'h68;        memory[38472] <=  8'h63;        memory[38473] <=  8'h66;        memory[38474] <=  8'h69;        memory[38475] <=  8'h77;        memory[38476] <=  8'h68;        memory[38477] <=  8'h61;        memory[38478] <=  8'h74;        memory[38479] <=  8'h61;        memory[38480] <=  8'h6e;        memory[38481] <=  8'h61;        memory[38482] <=  8'h62;        memory[38483] <=  8'h61;        memory[38484] <=  8'h63;        memory[38485] <=  8'h61;        memory[38486] <=  8'h74;        memory[38487] <=  8'h61;        memory[38488] <=  8'h62;        memory[38489] <=  8'h61;        memory[38490] <=  8'h72;        memory[38491] <=  8'h63;        memory[38492] <=  8'h61;        memory[38493] <=  8'h68;        memory[38494] <=  8'h64;        memory[38495] <=  8'h75;        memory[38496] <=  8'h63;        memory[38497] <=  8'h74;        memory[38498] <=  8'h61;        memory[38499] <=  8'h64;        memory[38500] <=  8'h61;        memory[38501] <=  8'h61;        memory[38502] <=  8'h63;        memory[38503] <=  8'h61;        memory[38504] <=  8'h72;        memory[38505] <=  8'h62;        memory[38506] <=  8'h61;        memory[38507] <=  8'h72;        memory[38508] <=  8'h74;        memory[38509] <=  8'h78;        memory[38510] <=  8'h61;        memory[38511] <=  8'h74;        memory[38512] <=  8'h6b;        memory[38513] <=  8'h73;        memory[38514] <=  8'h68;        memory[38515] <=  8'h63;        memory[38516] <=  8'h66;        memory[38517] <=  8'h69;        memory[38518] <=  8'h77;        memory[38519] <=  8'h68;        memory[38520] <=  8'h61;        memory[38521] <=  8'h74;        memory[38522] <=  8'h61;        memory[38523] <=  8'h6e;        memory[38524] <=  8'h61;        memory[38525] <=  8'h62;        memory[38526] <=  8'h61;        memory[38527] <=  8'h63;        memory[38528] <=  8'h61;        memory[38529] <=  8'h74;        memory[38530] <=  8'h61;        memory[38531] <=  8'h62;        memory[38532] <=  8'h61;        memory[38533] <=  8'h72;        memory[38534] <=  8'h63;        memory[38535] <=  8'h61;        memory[38536] <=  8'h68;        memory[38537] <=  8'h64;        memory[38538] <=  8'h75;        memory[38539] <=  8'h63;        memory[38540] <=  8'h74;        memory[38541] <=  8'h61;        memory[38542] <=  8'h64;        memory[38543] <=  8'h61;        memory[38544] <=  8'h61;        memory[38545] <=  8'h63;        memory[38546] <=  8'h61;        memory[38547] <=  8'h72;        memory[38548] <=  8'h62;        memory[38549] <=  8'h61;        memory[38550] <=  8'h72;        memory[38551] <=  8'h74;        memory[38552] <=  8'h78;        memory[38553] <=  8'h61;        memory[38554] <=  8'h74;        memory[38555] <=  8'h6b;        memory[38556] <=  8'h73;        memory[38557] <=  8'h68;        memory[38558] <=  8'h63;        memory[38559] <=  8'h66;        memory[38560] <=  8'h69;        memory[38561] <=  8'h77;        memory[38562] <=  8'h68;        memory[38563] <=  8'h61;        memory[38564] <=  8'h74;        memory[38565] <=  8'h61;        memory[38566] <=  8'h6e;        memory[38567] <=  8'h61;        memory[38568] <=  8'h62;        memory[38569] <=  8'h61;        memory[38570] <=  8'h63;        memory[38571] <=  8'h61;        memory[38572] <=  8'h74;        memory[38573] <=  8'h61;        memory[38574] <=  8'h62;        memory[38575] <=  8'h61;        memory[38576] <=  8'h72;        memory[38577] <=  8'h63;        memory[38578] <=  8'h61;        memory[38579] <=  8'h68;        memory[38580] <=  8'h64;        memory[38581] <=  8'h75;        memory[38582] <=  8'h63;        memory[38583] <=  8'h74;        memory[38584] <=  8'h61;        memory[38585] <=  8'h64;        memory[38586] <=  8'h61;        memory[38587] <=  8'h61;        memory[38588] <=  8'h63;        memory[38589] <=  8'h61;        memory[38590] <=  8'h72;        memory[38591] <=  8'h62;        memory[38592] <=  8'h61;        memory[38593] <=  8'h72;        memory[38594] <=  8'h74;        memory[38595] <=  8'h78;        memory[38596] <=  8'h61;        memory[38597] <=  8'h74;        memory[38598] <=  8'h6b;        memory[38599] <=  8'h73;        memory[38600] <=  8'h68;        memory[38601] <=  8'h63;        memory[38602] <=  8'h66;        memory[38603] <=  8'h69;        memory[38604] <=  8'h77;        memory[38605] <=  8'h68;        memory[38606] <=  8'h61;        memory[38607] <=  8'h74;        memory[38608] <=  8'h61;        memory[38609] <=  8'h6e;        memory[38610] <=  8'h61;        memory[38611] <=  8'h62;        memory[38612] <=  8'h61;        memory[38613] <=  8'h63;        memory[38614] <=  8'h61;        memory[38615] <=  8'h74;        memory[38616] <=  8'h61;        memory[38617] <=  8'h62;        memory[38618] <=  8'h61;        memory[38619] <=  8'h72;        memory[38620] <=  8'h63;        memory[38621] <=  8'h61;        memory[38622] <=  8'h68;        memory[38623] <=  8'h64;        memory[38624] <=  8'h75;        memory[38625] <=  8'h63;        memory[38626] <=  8'h74;        memory[38627] <=  8'h61;        memory[38628] <=  8'h64;        memory[38629] <=  8'h61;        memory[38630] <=  8'h61;        memory[38631] <=  8'h63;        memory[38632] <=  8'h61;        memory[38633] <=  8'h72;        memory[38634] <=  8'h62;        memory[38635] <=  8'h61;        memory[38636] <=  8'h72;        memory[38637] <=  8'h74;        memory[38638] <=  8'h78;        memory[38639] <=  8'h61;        memory[38640] <=  8'h74;        memory[38641] <=  8'h6b;        memory[38642] <=  8'h73;        memory[38643] <=  8'h68;        memory[38644] <=  8'h63;        memory[38645] <=  8'h66;        memory[38646] <=  8'h69;        memory[38647] <=  8'h77;        memory[38648] <=  8'h68;        memory[38649] <=  8'h61;        memory[38650] <=  8'h74;        memory[38651] <=  8'h61;        memory[38652] <=  8'h6e;        memory[38653] <=  8'h61;        memory[38654] <=  8'h62;        memory[38655] <=  8'h61;        memory[38656] <=  8'h63;        memory[38657] <=  8'h61;        memory[38658] <=  8'h74;        memory[38659] <=  8'h61;        memory[38660] <=  8'h62;        memory[38661] <=  8'h61;        memory[38662] <=  8'h72;        memory[38663] <=  8'h63;        memory[38664] <=  8'h61;        memory[38665] <=  8'h68;        memory[38666] <=  8'h64;        memory[38667] <=  8'h75;        memory[38668] <=  8'h63;        memory[38669] <=  8'h74;        memory[38670] <=  8'h61;        memory[38671] <=  8'h64;        memory[38672] <=  8'h61;        memory[38673] <=  8'h61;        memory[38674] <=  8'h63;        memory[38675] <=  8'h61;        memory[38676] <=  8'h72;        memory[38677] <=  8'h62;        memory[38678] <=  8'h61;        memory[38679] <=  8'h72;        memory[38680] <=  8'h74;        memory[38681] <=  8'h74;        memory[38682] <=  8'h62;        memory[38683] <=  8'h61;        memory[38684] <=  8'h72;        memory[38685] <=  8'h74;        memory[38686] <=  8'h78;        memory[38687] <=  8'h61;        memory[38688] <=  8'h74;        memory[38689] <=  8'h6b;        memory[38690] <=  8'h73;        memory[38691] <=  8'h68;        memory[38692] <=  8'h63;        memory[38693] <=  8'h66;        memory[38694] <=  8'h69;        memory[38695] <=  8'h77;        memory[38696] <=  8'h68;        memory[38697] <=  8'h61;        memory[38698] <=  8'h74;        memory[38699] <=  8'h61;        memory[38700] <=  8'h6e;        memory[38701] <=  8'h61;        memory[38702] <=  8'h62;        memory[38703] <=  8'h61;        memory[38704] <=  8'h63;        memory[38705] <=  8'h61;        memory[38706] <=  8'h74;        memory[38707] <=  8'h61;        memory[38708] <=  8'h62;        memory[38709] <=  8'h61;        memory[38710] <=  8'h72;        memory[38711] <=  8'h63;        memory[38712] <=  8'h61;        memory[38713] <=  8'h68;        memory[38714] <=  8'h64;        memory[38715] <=  8'h75;        memory[38716] <=  8'h63;        memory[38717] <=  8'h74;        memory[38718] <=  8'h61;        memory[38719] <=  8'h64;        memory[38720] <=  8'h61;        memory[38721] <=  8'h61;        memory[38722] <=  8'h63;        memory[38723] <=  8'h61;        memory[38724] <=  8'h72;        memory[38725] <=  8'h63;        memory[38726] <=  8'h74;        memory[38727] <=  8'h72;        memory[38728] <=  8'h63;        memory[38729] <=  8'h61;        memory[38730] <=  8'h74;        memory[38731] <=  8'h72;        memory[38732] <=  8'h63;        memory[38733] <=  8'h61;        memory[38734] <=  8'h74;        memory[38735] <=  8'h63;        memory[38736] <=  8'h62;        memory[38737] <=  8'h61;        memory[38738] <=  8'h74;        memory[38739] <=  8'h62;        memory[38740] <=  8'h72;        memory[38741] <=  8'h63;        memory[38742] <=  8'h61;        memory[38743] <=  8'h72;        memory[38744] <=  8'h62;        memory[38745] <=  8'h78;        memory[38746] <=  8'h74;        memory[38747] <=  8'h61;        memory[38748] <=  8'h72;        memory[38749] <=  8'h64;        memory[38750] <=  8'h66;        memory[38751] <=  8'h73;        memory[38752] <=  8'h67;        memory[38753] <=  8'h76;        memory[38754] <=  8'h68;        memory[38755] <=  8'h62;        memory[38756] <=  8'h6b;        memory[38757] <=  8'h6a;        memory[38758] <=  8'h6e;        memory[38759] <=  8'h6d;        memory[38760] <=  8'h62;        memory[38761] <=  8'h76;        memory[38762] <=  8'h78;        memory[38763] <=  8'h63;        memory[38764] <=  8'h73;        memory[38765] <=  8'h66;        memory[38766] <=  8'h72;        memory[38767] <=  8'h74;        memory[38768] <=  8'h79;        memory[38769] <=  8'h75;        memory[38770] <=  8'h6a;        memory[38771] <=  8'h6e;        memory[38772] <=  8'h62;        memory[38773] <=  8'h76;        memory[38774] <=  8'h63;        memory[38775] <=  8'h64;        memory[38776] <=  8'h74;        memory[38777] <=  8'h79;        memory[38778] <=  8'h75;        memory[38779] <=  8'h69;        memory[38780] <=  8'h6b;        memory[38781] <=  8'h6d;        memory[38782] <=  8'h6e;        memory[38783] <=  8'h62;        memory[38784] <=  8'h76;        memory[38785] <=  8'h63;        memory[38786] <=  8'h78;        memory[38787] <=  8'h73;        memory[38788] <=  8'h64;        memory[38789] <=  8'h72;        memory[38790] <=  8'h74;        memory[38791] <=  8'h79;        memory[38792] <=  8'h75;        memory[38793] <=  8'h69;        memory[38794] <=  8'h6b;        memory[38795] <=  8'h6d;        memory[38796] <=  8'h6e;        memory[38797] <=  8'h62;        memory[38798] <=  8'h76;        memory[38799] <=  8'h63;        memory[38800] <=  8'h73;        memory[38801] <=  8'h77;        memory[38802] <=  8'h33;        memory[38803] <=  8'h34;        memory[38804] <=  8'h35;        memory[38805] <=  8'h36;        memory[38806] <=  8'h37;        memory[38807] <=  8'h38;        memory[38808] <=  8'h69;        memory[38809] <=  8'h6b;        memory[38810] <=  8'h6d;        memory[38811] <=  8'h6e;        memory[38812] <=  8'h62;        memory[38813] <=  8'h76;        memory[38814] <=  8'h63;        memory[38815] <=  8'h64;        memory[38816] <=  8'h65;        memory[38817] <=  8'h72;        memory[38818] <=  8'h36;        memory[38819] <=  8'h37;        memory[38820] <=  8'h38;        memory[38821] <=  8'h69;        memory[38822] <=  8'h6f;        memory[38823] <=  8'h6b;        memory[38824] <=  8'h6a;        memory[38825] <=  8'h6e;        memory[38826] <=  8'h62;        memory[38827] <=  8'h76;        memory[38828] <=  8'h63;        memory[38829] <=  8'h64;        memory[38830] <=  8'h72;        memory[38831] <=  8'h74;        memory[38832] <=  8'h79;        memory[38833] <=  8'h75;        memory[38834] <=  8'h73;        memory[38835] <=  8'h6a;        memory[38836] <=  8'h63;        memory[38837] <=  8'h6e;        memory[38838] <=  8'h62;        memory[38839] <=  8'h64;        memory[38840] <=  8'h66;        memory[38841] <=  8'h73;        memory[38842] <=  8'h74;        memory[38843] <=  8'h79;        memory[38844] <=  8'h75;        memory[38845] <=  8'h61;        memory[38846] <=  8'h69;        memory[38847] <=  8'h6b;        memory[38848] <=  8'h78;        memory[38849] <=  8'h6d;        memory[38850] <=  8'h6e;        memory[38851] <=  8'h73;        memory[38852] <=  8'h6a;        memory[38853] <=  8'h6f;        memory[38854] <=  8'h64;        memory[38855] <=  8'h6c;        memory[38856] <=  8'h63;        memory[38857] <=  8'h78;        memory[38858] <=  8'h2c;        memory[38859] <=  8'h6d;        memory[38860] <=  8'h73;        memory[38861] <=  8'h6b;        memory[38862] <=  8'h64;        memory[38863] <=  8'h6c;        memory[38864] <=  8'h70;        memory[38865] <=  8'h5b;        memory[38866] <=  8'h3b;        memory[38867] <=  8'h73;        memory[38868] <=  8'h6c;        memory[38869] <=  8'h64;        memory[38870] <=  8'h70;        memory[38871] <=  8'h76;        memory[38872] <=  8'h63;        memory[38873] <=  8'h5b;        memory[38874] <=  8'h78;        memory[38875] <=  8'h76;        memory[38876] <=  8'h63;        memory[38877] <=  8'h5b;        memory[38878] <=  8'h78;        memory[38879] <=  8'h70;        memory[38880] <=  8'h6f;        memory[38881] <=  8'h20;        memory[38882] <=  8'h62;        memory[38883] <=  8'h61;        memory[38884] <=  8'h72;        memory[38885] <=  8'h74;        memory[38886] <=  8'h74;        memory[38887] <=  8'h62;        memory[38888] <=  8'h61;        memory[38889] <=  8'h72;        memory[38890] <=  8'h74;        memory[38891] <=  8'h78;        memory[38892] <=  8'h61;        memory[38893] <=  8'h74;        memory[38894] <=  8'h6b;        memory[38895] <=  8'h73;        memory[38896] <=  8'h68;        memory[38897] <=  8'h63;        memory[38898] <=  8'h66;        memory[38899] <=  8'h69;        memory[38900] <=  8'h77;        memory[38901] <=  8'h68;        memory[38902] <=  8'h61;        memory[38903] <=  8'h69;        memory[38904] <=  8'h6a;        memory[38905] <=  8'h78;        memory[38906] <=  8'h5d;        memory[38907] <=  8'h65;        memory[38908] <=  8'h6b;        memory[38909] <=  8'h6f;        memory[38910] <=  8'h39;        memory[38911] <=  8'h64;        memory[38912] <=  8'h75;        memory[38913] <=  8'h38;        memory[38914] <=  8'h79;        memory[38915] <=  8'h20;        memory[38916] <=  8'h37;        memory[38917] <=  8'h63;        memory[38918] <=  8'h67;        memory[38919] <=  8'h78;        memory[38920] <=  8'h63;        memory[38921] <=  8'h75;        memory[38922] <=  8'h68;        memory[38923] <=  8'h69;        memory[38924] <=  8'h6a;        memory[38925] <=  8'h77;        memory[38926] <=  8'h69;        memory[38927] <=  8'h64;        memory[38928] <=  8'h66;        memory[38929] <=  8'h68;        memory[38930] <=  8'h75;        memory[38931] <=  8'h76;        memory[38932] <=  8'h64;        memory[38933] <=  8'h62;        memory[38934] <=  8'h66;        memory[38935] <=  8'h6a;        memory[38936] <=  8'h6e;        memory[38937] <=  8'h6b;        memory[38938] <=  8'h6a;        memory[38939] <=  8'h65;        memory[38940] <=  8'h38;        memory[38941] <=  8'h66;        memory[38942] <=  8'h37;        memory[38943] <=  8'h67;        memory[38944] <=  8'h79;        memory[38945] <=  8'h76;        memory[38946] <=  8'h63;        memory[38947] <=  8'h68;        memory[38948] <=  8'h69;        memory[38949] <=  8'h6a;        memory[38950] <=  8'h33;        memory[38951] <=  8'h65;        memory[38952] <=  8'h67;        memory[38953] <=  8'h79;        memory[38954] <=  8'h72;        memory[38955] <=  8'h64;        memory[38956] <=  8'h62;        memory[38957] <=  8'h6e;        memory[38958] <=  8'h63;        memory[38959] <=  8'h7a;        memory[38960] <=  8'h6a;        memory[38961] <=  8'h6f;        memory[38962] <=  8'h66;        memory[38963] <=  8'h78;        memory[38964] <=  8'h6a;        memory[38965] <=  8'h69;        memory[38966] <=  8'h63;        memory[38967] <=  8'h68;        memory[38968] <=  8'h62;        memory[38969] <=  8'h6e;        memory[38970] <=  8'h6d;        memory[38971] <=  8'h63;        memory[38972] <=  8'h73;        memory[38973] <=  8'h6c;        memory[38974] <=  8'h6b;        memory[38975] <=  8'h6a;        memory[38976] <=  8'h69;        memory[38977] <=  8'h68;        memory[38978] <=  8'h76;        memory[38979] <=  8'h75;        memory[38980] <=  8'h69;        memory[38981] <=  8'h64;        memory[38982] <=  8'h68;        memory[38983] <=  8'h75;        memory[38984] <=  8'h67;        memory[38985] <=  8'h79;        memory[38986] <=  8'h62;        memory[38987] <=  8'h68;        memory[38988] <=  8'h65;        memory[38989] <=  8'h6a;        memory[38990] <=  8'h72;        memory[38991] <=  8'h6b;        memory[38992] <=  8'h6a;        memory[38993] <=  8'h6f;        memory[38994] <=  8'h64;        memory[38995] <=  8'h67;        memory[38996] <=  8'h69;        memory[38997] <=  8'h75;        memory[38998] <=  8'h69;        memory[38999] <=  8'h67;        memory[39000] <=  8'h76;        memory[39001] <=  8'h79;        memory[39002] <=  8'h75;        memory[39003] <=  8'h67;        memory[39004] <=  8'h78;        memory[39005] <=  8'h68;        memory[39006] <=  8'h63;        memory[39007] <=  8'h20;        memory[39008] <=  8'h20;        memory[39009] <=  8'h20;        memory[39010] <=  8'h78;        memory[39011] <=  8'h76;        memory[39012] <=  8'h20;        memory[39013] <=  8'h63;        memory[39014] <=  8'h78;        memory[39015] <=  8'h67;        memory[39016] <=  8'h79;        memory[39017] <=  8'h63;        memory[39018] <=  8'h75;        memory[39019] <=  8'h68;        memory[39020] <=  8'h6a;        memory[39021] <=  8'h6b;        memory[39022] <=  8'h61;        memory[39023] <=  8'h6c;        memory[39024] <=  8'h78;        memory[39025] <=  8'h76;        memory[39026] <=  8'h70;        memory[39027] <=  8'h6f;        memory[39028] <=  8'h69;        memory[39029] <=  8'h6a;        memory[39030] <=  8'h69;        memory[39031] <=  8'h68;        memory[39032] <=  8'h6a;        memory[39033] <=  8'h62;        memory[39034] <=  8'h77;        memory[39035] <=  8'h65;        memory[39036] <=  8'h6e;        memory[39037] <=  8'h61;        memory[39038] <=  8'h66;        memory[39039] <=  8'h6d;        memory[39040] <=  8'h64;        memory[39041] <=  8'h6b;        memory[39042] <=  8'h6d;        memory[39043] <=  8'h76;        memory[39044] <=  8'h6c;        memory[39045] <=  8'h63;        memory[39046] <=  8'h6f;        memory[39047] <=  8'h64;        memory[39048] <=  8'h69;        memory[39049] <=  8'h75;        memory[39050] <=  8'h68;        memory[39051] <=  8'h73;        memory[39052] <=  8'h66;        memory[39053] <=  8'h65;        memory[39054] <=  8'h62;        memory[39055] <=  8'h6e;        memory[39056] <=  8'h64;        memory[39057] <=  8'h73;        memory[39058] <=  8'h63;        memory[39059] <=  8'h6b;        memory[39060] <=  8'h20;        memory[39061] <=  8'h78;        memory[39062] <=  8'h6a;        memory[39063] <=  8'h78;        memory[39064] <=  8'h63;        memory[39065] <=  8'h73;        memory[39066] <=  8'h64;        memory[39067] <=  8'h66;        memory[39068] <=  8'h6b;        memory[39069] <=  8'h64;        memory[39070] <=  8'h6e;        memory[39071] <=  8'h6d;        memory[39072] <=  8'h64;        memory[39073] <=  8'h73;        memory[39074] <=  8'h63;        memory[39075] <=  8'h6b;        memory[39076] <=  8'h78;        memory[39077] <=  8'h6c;        memory[39078] <=  8'h6f;        memory[39079] <=  8'h66;        memory[39080] <=  8'h6a;        memory[39081] <=  8'h69;        memory[39082] <=  8'h61;        memory[39083] <=  8'h62;        memory[39084] <=  8'h6e;        memory[39085] <=  8'h20;        memory[39086] <=  8'h78;        memory[39087] <=  8'h6b;        memory[39088] <=  8'h6d;        memory[39089] <=  8'h20;        memory[39090] <=  8'h6f;        memory[39091] <=  8'h63;        memory[39092] <=  8'h76;        memory[39093] <=  8'h73;        memory[39094] <=  8'h64;        memory[39095] <=  8'h69;        memory[39096] <=  8'h66;        memory[39097] <=  8'h68;        memory[39098] <=  8'h65;        memory[39099] <=  8'h71;        memory[39100] <=  8'h6a;        memory[39101] <=  8'h77;        memory[39102] <=  8'h62;        memory[39103] <=  8'h65;        memory[39104] <=  8'h6e;        memory[39105] <=  8'h20;        memory[39106] <=  8'h6d;        memory[39107] <=  8'h64;        memory[39108] <=  8'h73;        memory[39109] <=  8'h6c;        memory[39110] <=  8'h76;        memory[39111] <=  8'h6b;        memory[39112] <=  8'h63;        memory[39113] <=  8'h78;        memory[39114] <=  8'h20;        memory[39115] <=  8'h6f;        memory[39116] <=  8'h78;        memory[39117] <=  8'h69;        memory[39118] <=  8'h63;        memory[39119] <=  8'h6a;        memory[39120] <=  8'h76;        memory[39121] <=  8'h64;        memory[39122] <=  8'h66;        memory[39123] <=  8'h65;        memory[39124] <=  8'h71;        memory[39125] <=  8'h6e;        memory[39126] <=  8'h20;        memory[39127] <=  8'h64;        memory[39128] <=  8'h6d;        memory[39129] <=  8'h73;        memory[39130] <=  8'h6c;        memory[39131] <=  8'h63;        memory[39132] <=  8'h78;        memory[39133] <=  8'h6b;        memory[39134] <=  8'h20;        memory[39135] <=  8'h6f;        memory[39136] <=  8'h78;        memory[39137] <=  8'h63;        memory[39138] <=  8'h76;        memory[39139] <=  8'h6a;        memory[39140] <=  8'h64;        memory[39141] <=  8'h62;        memory[39142] <=  8'h71;        memory[39143] <=  8'h77;        memory[39144] <=  8'h65;        memory[39145] <=  8'h6e;        memory[39146] <=  8'h6d;        memory[39147] <=  8'h64;        memory[39148] <=  8'h6c;        memory[39149] <=  8'h73;        memory[39150] <=  8'h2c;        memory[39151] <=  8'h76;        memory[39152] <=  8'h63;        memory[39153] <=  8'h78;        memory[39154] <=  8'h20;        memory[39155] <=  8'h63;        memory[39156] <=  8'h6f;        memory[39157] <=  8'h69;        memory[39158] <=  8'h76;        memory[39159] <=  8'h68;        memory[39160] <=  8'h73;        memory[39161] <=  8'h64;        memory[39162] <=  8'h62;        memory[39163] <=  8'h71;        memory[39164] <=  8'h77;        memory[39165] <=  8'h65;        memory[39166] <=  8'h6e;        memory[39167] <=  8'h64;        memory[39168] <=  8'h6b;        memory[39169] <=  8'h73;        memory[39170] <=  8'h76;        memory[39171] <=  8'h6f;        memory[39172] <=  8'h63;        memory[39173] <=  8'h20;        memory[39174] <=  8'h76;        memory[39175] <=  8'h69;        memory[39176] <=  8'h75;        memory[39177] <=  8'h69;        memory[39178] <=  8'h68;        memory[39179] <=  8'h63;        memory[39180] <=  8'h78;        memory[39181] <=  8'h69;        memory[39182] <=  8'h6f;        memory[39183] <=  8'h76;        memory[39184] <=  8'h73;        memory[39185] <=  8'h64;        memory[39186] <=  8'h61;        memory[39187] <=  8'h64;        memory[39188] <=  8'h6e;        memory[39189] <=  8'h77;        memory[39190] <=  8'h71;        memory[39191] <=  8'h6b;        memory[39192] <=  8'h6c;        memory[39193] <=  8'h73;        memory[39194] <=  8'h76;        memory[39195] <=  8'h6e;        memory[39196] <=  8'h62;        memory[39197] <=  8'h20;        memory[39198] <=  8'h64;        memory[39199] <=  8'h66;        memory[39200] <=  8'h6a;        memory[39201] <=  8'h6b;        memory[39202] <=  8'h71;        memory[39203] <=  8'h64;        memory[39204] <=  8'h77;        memory[39205] <=  8'h65;        memory[39206] <=  8'h6e;        memory[39207] <=  8'h62;        memory[39208] <=  8'h20;        memory[39209] <=  8'h64;        memory[39210] <=  8'h73;        memory[39211] <=  8'h76;        memory[39212] <=  8'h68;        memory[39213] <=  8'h64;        memory[39214] <=  8'h61;        memory[39215] <=  8'h71;        memory[39216] <=  8'h77;        memory[39217] <=  8'h6a;        memory[39218] <=  8'h65;        memory[39219] <=  8'h6e;        memory[39220] <=  8'h64;        memory[39221] <=  8'h20;        memory[39222] <=  8'h61;        memory[39223] <=  8'h63;        memory[39224] <=  8'h62;        memory[39225] <=  8'h68;        memory[39226] <=  8'h64;        memory[39227] <=  8'h61;        memory[39228] <=  8'h77;        memory[39229] <=  8'h71;        memory[39230] <=  8'h6e;        memory[39231] <=  8'h20;        memory[39232] <=  8'h62;        memory[39233] <=  8'h73;        memory[39234] <=  8'h76;        memory[39235] <=  8'h61;        memory[39236] <=  8'h67;        memory[39237] <=  8'h76;        memory[39238] <=  8'h68;        memory[39239] <=  8'h67;        memory[39240] <=  8'h61;        memory[39241] <=  8'h73;        memory[39242] <=  8'h6a;        memory[39243] <=  8'h6b;        memory[39244] <=  8'h63;        memory[39245] <=  8'h78;        memory[39246] <=  8'h76;        memory[39247] <=  8'h6e;        memory[39248] <=  8'h73;        memory[39249] <=  8'h64;        memory[39250] <=  8'h20;        memory[39251] <=  8'h66;        memory[39252] <=  8'h62;        memory[39253] <=  8'h64;        memory[39254] <=  8'h61;        memory[39255] <=  8'h73;        memory[39256] <=  8'h76;        memory[39257] <=  8'h67;        memory[39258] <=  8'h63;        memory[39259] <=  8'h79;        memory[39260] <=  8'h7a;        memory[39261] <=  8'h78;        memory[39262] <=  8'h79;        memory[39263] <=  8'h75;        memory[39264] <=  8'h20;        memory[39265] <=  8'h69;        memory[39266] <=  8'h6a;        memory[39267] <=  8'h64;        memory[39268] <=  8'h66;        memory[39269] <=  8'h6b;        memory[39270] <=  8'h61;        memory[39271] <=  8'h64;        memory[39272] <=  8'h63;        memory[39273] <=  8'h78;        memory[39274] <=  8'h68;        memory[39275] <=  8'h20;        memory[39276] <=  8'h67;        memory[39277] <=  8'h61;        memory[39278] <=  8'h68;        memory[39279] <=  8'h75;        memory[39280] <=  8'h64;        memory[39281] <=  8'h73;        memory[39282] <=  8'h69;        memory[39283] <=  8'h6a;        memory[39284] <=  8'h61;        memory[39285] <=  8'h6b;        memory[39286] <=  8'h63;        memory[39287] <=  8'h62;        memory[39288] <=  8'h61;        memory[39289] <=  8'h72;        memory[39290] <=  8'h73;        memory[39291] <=  8'h68;        memory[39292] <=  8'h64;        memory[39293] <=  8'h66;        memory[39294] <=  8'h67;        memory[39295] <=  8'h73;        memory[39296] <=  8'h68;        memory[39297] <=  8'h64;        memory[39298] <=  8'h66;        memory[39299] <=  8'h68;        memory[39300] <=  8'h64;        memory[39301] <=  8'h6a;        memory[39302] <=  8'h68;        memory[39303] <=  8'h62;        memory[39304] <=  8'h67;        memory[39305] <=  8'h63;        memory[39306] <=  8'h61;        memory[39307] <=  8'h66;        memory[39308] <=  8'h73;        memory[39309] <=  8'h79;        memory[39310] <=  8'h67;        memory[39311] <=  8'h6b;        memory[39312] <=  8'h75;        memory[39313] <=  8'h64;        memory[39314] <=  8'h68;        memory[39315] <=  8'h62;        memory[39316] <=  8'h77;        memory[39317] <=  8'h76;        memory[39318] <=  8'h67;        memory[39319] <=  8'h61;        memory[39320] <=  8'h66;        memory[39321] <=  8'h64;        memory[39322] <=  8'h74;        memory[39323] <=  8'h75;        memory[39324] <=  8'h66;        memory[39325] <=  8'h79;        memory[39326] <=  8'h67;        memory[39327] <=  8'h69;        memory[39328] <=  8'h75;        memory[39329] <=  8'h68;        memory[39330] <=  8'h6c;        memory[39331] <=  8'h6a;        memory[39332] <=  8'h62;        memory[39333] <=  8'h6b;        memory[39334] <=  8'h68;        memory[39335] <=  8'h76;        memory[39336] <=  8'h67;        memory[39337] <=  8'h63;        memory[39338] <=  8'h66;        memory[39339] <=  8'h78;        memory[39340] <=  8'h64;        memory[39341] <=  8'h74;        memory[39342] <=  8'h75;        memory[39343] <=  8'h79;        memory[39344] <=  8'h69;        memory[39345] <=  8'h75;        memory[39346] <=  8'h68;        memory[39347] <=  8'h6c;        memory[39348] <=  8'h6a;        memory[39349] <=  8'h6b;        memory[39350] <=  8'h67;        memory[39351] <=  8'h6a;        memory[39352] <=  8'h63;        memory[39353] <=  8'h66;        memory[39354] <=  8'h68;        memory[39355] <=  8'h64;        memory[39356] <=  8'h67;        memory[39357] <=  8'h72;        memory[39358] <=  8'h79;        memory[39359] <=  8'h74;        memory[39360] <=  8'h66;        memory[39361] <=  8'h75;        memory[39362] <=  8'h79;        memory[39363] <=  8'h69;        memory[39364] <=  8'h68;        memory[39365] <=  8'h6c;        memory[39366] <=  8'h62;        memory[39367] <=  8'h6d;        memory[39368] <=  8'h76;        memory[39369] <=  8'h6e;        memory[39370] <=  8'h63;        memory[39371] <=  8'h66;        memory[39372] <=  8'h68;        memory[39373] <=  8'h64;        memory[39374] <=  8'h74;        memory[39375] <=  8'h75;        memory[39376] <=  8'h67;        memory[39377] <=  8'h79;        memory[39378] <=  8'h69;        memory[39379] <=  8'h68;        memory[39380] <=  8'h75;        memory[39381] <=  8'h6a;        memory[39382] <=  8'h6c;        memory[39383] <=  8'h62;        memory[39384] <=  8'h6d;        memory[39385] <=  8'h76;        memory[39386] <=  8'h6e;        memory[39387] <=  8'h63;        memory[39388] <=  8'h66;        memory[39389] <=  8'h68;        memory[39390] <=  8'h67;        memory[39391] <=  8'h79;        memory[39392] <=  8'h68;        memory[39393] <=  8'h75;        memory[39394] <=  8'h6a;        memory[39395] <=  8'h6e;        memory[39396] <=  8'h2c;        memory[39397] <=  8'h62;        memory[39398] <=  8'h6e;        memory[39399] <=  8'h6d;        memory[39400] <=  8'h76;        memory[39401] <=  8'h6e;        memory[39402] <=  8'h63;        memory[39403] <=  8'h66;        memory[39404] <=  8'h68;        memory[39405] <=  8'h74;        memory[39406] <=  8'h79;        memory[39407] <=  8'h69;        memory[39408] <=  8'h75;        memory[39409] <=  8'h6c;        memory[39410] <=  8'h6a;        memory[39411] <=  8'h62;        memory[39412] <=  8'h6d;        memory[39413] <=  8'h76;        memory[39414] <=  8'h6e;        memory[39415] <=  8'h63;        memory[39416] <=  8'h66;        memory[39417] <=  8'h74;        memory[39418] <=  8'h75;        memory[39419] <=  8'h79;        memory[39420] <=  8'h69;        memory[39421] <=  8'h68;        memory[39422] <=  8'h6b;        memory[39423] <=  8'h62;        memory[39424] <=  8'h76;        memory[39425] <=  8'h63;        memory[39426] <=  8'h66;        memory[39427] <=  8'h67;        memory[39428] <=  8'h74;        memory[39429] <=  8'h75;        memory[39430] <=  8'h79;        memory[39431] <=  8'h69;        memory[39432] <=  8'h75;        memory[39433] <=  8'h68;        memory[39434] <=  8'h6a;        memory[39435] <=  8'h6b;        memory[39436] <=  8'h62;        memory[39437] <=  8'h76;        memory[39438] <=  8'h63;        memory[39439] <=  8'h66;        memory[39440] <=  8'h74;        memory[39441] <=  8'h75;        memory[39442] <=  8'h79;        memory[39443] <=  8'h69;        memory[39444] <=  8'h75;        memory[39445] <=  8'h6a;        memory[39446] <=  8'h6b;        memory[39447] <=  8'h6e;        memory[39448] <=  8'h62;        memory[39449] <=  8'h76;        memory[39450] <=  8'h67;        memory[39451] <=  8'h66;        memory[39452] <=  8'h74;        memory[39453] <=  8'h79;        memory[39454] <=  8'h75;        memory[39455] <=  8'h75;        memory[39456] <=  8'h69;        memory[39457] <=  8'h6a;        memory[39458] <=  8'h6b;        memory[39459] <=  8'h68;        memory[39460] <=  8'h62;        memory[39461] <=  8'h6a;        memory[39462] <=  8'h67;        memory[39463] <=  8'h68;        memory[39464] <=  8'h66;        memory[39465] <=  8'h79;        memory[39466] <=  8'h74;        memory[39467] <=  8'h79;        memory[39468] <=  8'h69;        memory[39469] <=  8'h75;        memory[39470] <=  8'h64;        memory[39471] <=  8'h6a;        memory[39472] <=  8'h6b;        memory[39473] <=  8'h68;        memory[39474] <=  8'h63;        memory[39475] <=  8'h7a;        memory[39476] <=  8'h67;        memory[39477] <=  8'h68;        memory[39478] <=  8'h74;        memory[39479] <=  8'h75;        memory[39480] <=  8'h79;        memory[39481] <=  8'h69;        memory[39482] <=  8'h61;        memory[39483] <=  8'h73;        memory[39484] <=  8'h75;        memory[39485] <=  8'h6a;        memory[39486] <=  8'h6b;        memory[39487] <=  8'h62;        memory[39488] <=  8'h6e;        memory[39489] <=  8'h61;        memory[39490] <=  8'h76;        memory[39491] <=  8'h63;        memory[39492] <=  8'h66;        memory[39493] <=  8'h68;        memory[39494] <=  8'h75;        memory[39495] <=  8'h61;        memory[39496] <=  8'h73;        memory[39497] <=  8'h79;        memory[39498] <=  8'h64;        memory[39499] <=  8'h75;        memory[39500] <=  8'h69;        memory[39501] <=  8'h6a;        memory[39502] <=  8'h61;        memory[39503] <=  8'h6b;        memory[39504] <=  8'h62;        memory[39505] <=  8'h63;        memory[39506] <=  8'h78;        memory[39507] <=  8'h68;        memory[39508] <=  8'h67;        memory[39509] <=  8'h79;        memory[39510] <=  8'h75;        memory[39511] <=  8'h7a;        memory[39512] <=  8'h63;        memory[39513] <=  8'h61;        memory[39514] <=  8'h73;        memory[39515] <=  8'h69;        memory[39516] <=  8'h75;        memory[39517] <=  8'h6f;        memory[39518] <=  8'h69;        memory[39519] <=  8'h6a;        memory[39520] <=  8'h61;        memory[39521] <=  8'h6c;        memory[39522] <=  8'h63;        memory[39523] <=  8'h78;        memory[39524] <=  8'h62;        memory[39525] <=  8'h63;        memory[39526] <=  8'h20;        memory[39527] <=  8'h6e;        memory[39528] <=  8'h76;        memory[39529] <=  8'h63;        memory[39530] <=  8'h61;        memory[39531] <=  8'h64;        memory[39532] <=  8'h73;        memory[39533] <=  8'h67;        memory[39534] <=  8'h79;        memory[39535] <=  8'h68;        memory[39536] <=  8'h75;        memory[39537] <=  8'h61;        memory[39538] <=  8'h6a;        memory[39539] <=  8'h6b;        memory[39540] <=  8'h78;        memory[39541] <=  8'h62;        memory[39542] <=  8'h20;        memory[39543] <=  8'h6e;        memory[39544] <=  8'h76;        memory[39545] <=  8'h63;        memory[39546] <=  8'h61;        memory[39547] <=  8'h73;        memory[39548] <=  8'h67;        memory[39549] <=  8'h68;        memory[39550] <=  8'h75;        memory[39551] <=  8'h6a;        memory[39552] <=  8'h6c;        memory[39553] <=  8'h6b;        memory[39554] <=  8'h63;        memory[39555] <=  8'h78;        memory[39556] <=  8'h20;        memory[39557] <=  8'h6a;        memory[39558] <=  8'h6b;        memory[39559] <=  8'h68;        memory[39560] <=  8'h61;        memory[39561] <=  8'h73;        memory[39562] <=  8'h76;        memory[39563] <=  8'h64;        memory[39564] <=  8'h6e;        memory[39565] <=  8'h20;        memory[39566] <=  8'h62;        memory[39567] <=  8'h6e;        memory[39568] <=  8'h6d;        memory[39569] <=  8'h6b;        memory[39570] <=  8'h77;        memory[39571] <=  8'h64;        memory[39572] <=  8'h6f;        memory[39573] <=  8'h77;        memory[39574] <=  8'h69;        memory[39575] <=  8'h6f;        memory[39576] <=  8'h75;        memory[39577] <=  8'h69;        memory[39578] <=  8'h68;        memory[39579] <=  8'h62;        memory[39580] <=  8'h6e;        memory[39581] <=  8'h6b;        memory[39582] <=  8'h77;        memory[39583] <=  8'h69;        memory[39584] <=  8'h6f;        memory[39585] <=  8'h75;        memory[39586] <=  8'h71;        memory[39587] <=  8'h69;        memory[39588] <=  8'h79;        memory[39589] <=  8'h67;        memory[39590] <=  8'h6a;        memory[39591] <=  8'h64;        memory[39592] <=  8'h61;        memory[39593] <=  8'h76;        memory[39594] <=  8'h62;        memory[39595] <=  8'h6e;        memory[39596] <=  8'h6b;        memory[39597] <=  8'h6f;        memory[39598] <=  8'h70;        memory[39599] <=  8'h64;        memory[39600] <=  8'h76;        memory[39601] <=  8'h69;        memory[39602] <=  8'h6f;        memory[39603] <=  8'h75;        memory[39604] <=  8'h69;        memory[39605] <=  8'h48;        memory[39606] <=  8'h42;        memory[39607] <=  8'h6b;        memory[39608] <=  8'h64;        memory[39609] <=  8'h6e;        memory[39610] <=  8'h6c;        memory[39611] <=  8'h71;        memory[39612] <=  8'h6b;        memory[39613] <=  8'h6d;        memory[39614] <=  8'h6a;        memory[39615] <=  8'h70;        memory[39616] <=  8'h69;        memory[39617] <=  8'h6f;        memory[39618] <=  8'h68;        memory[39619] <=  8'h65;        memory[39620] <=  8'h66;        memory[39621] <=  8'h75;        memory[39622] <=  8'h67;        memory[39623] <=  8'h69;        memory[39624] <=  8'h73;        memory[39625] <=  8'h61;        memory[39626] <=  8'h62;        memory[39627] <=  8'h64;        memory[39628] <=  8'h6b;        memory[39629] <=  8'h6a;        memory[39630] <=  8'h6b;        memory[39631] <=  8'h6c;        memory[39632] <=  8'h6a;        memory[39633] <=  8'h69;        memory[39634] <=  8'h73;        memory[39635] <=  8'h6f;        memory[39636] <=  8'h71;        memory[39637] <=  8'h68;        memory[39638] <=  8'h77;        memory[39639] <=  8'h67;        memory[39640] <=  8'h69;        memory[39641] <=  8'h79;        memory[39642] <=  8'h6a;        memory[39643] <=  8'h64;        memory[39644] <=  8'h76;        memory[39645] <=  8'h62;        memory[39646] <=  8'h6e;        memory[39647] <=  8'h61;        memory[39648] <=  8'h73;        memory[39649] <=  8'h66;        memory[39650] <=  8'h6c;        memory[39651] <=  8'h6b;        memory[39652] <=  8'h64;        memory[39653] <=  8'h6a;        memory[39654] <=  8'h68;        memory[39655] <=  8'h63;        memory[39656] <=  8'h67;        memory[39657] <=  8'h6a;        memory[39658] <=  8'h76;        memory[39659] <=  8'h73;        memory[39660] <=  8'h64;        memory[39661] <=  8'h62;        memory[39662] <=  8'h62;        memory[39663] <=  8'h61;        memory[39664] <=  8'h72;        memory[39665] <=  8'h62;        memory[39666] <=  8'h62;        memory[39667] <=  8'h73;        memory[39668] <=  8'h62;        memory[39669] <=  8'h67;        memory[39670] <=  8'h73;        memory[39671] <=  8'h66;        memory[39672] <=  8'h67;        memory[39673] <=  8'h61;        memory[39674] <=  8'h68;        memory[39675] <=  8'h66;        memory[39676] <=  8'h73;        memory[39677] <=  8'h68;        memory[39678] <=  8'h61;        memory[39679] <=  8'h66;        memory[39680] <=  8'h73;        memory[39681] <=  8'h66;        memory[39682] <=  8'h68;        memory[39683] <=  8'h61;        memory[39684] <=  8'h69;        memory[39685] <=  8'h64;        memory[39686] <=  8'h75;        memory[39687] <=  8'h67;        memory[39688] <=  8'h64;        memory[39689] <=  8'h77;        memory[39690] <=  8'h62;        memory[39691] <=  8'h61;        memory[39692] <=  8'h62;        memory[39693] <=  8'h72;        memory[39694] <=  8'h62;        memory[39695] <=  8'h61;        memory[39696] <=  8'h62;        memory[39697] <=  8'h62;        memory[39698] <=  8'h74;        memory[39699] <=  8'h62;        memory[39700] <=  8'h62;        memory[39701] <=  8'h62;        memory[39702] <=  8'h62;        memory[39703] <=  8'h62;        memory[39704] <=  8'h62;        memory[39705] <=  8'h62;        memory[39706] <=  8'h62;        memory[39707] <=  8'h61;        memory[39708] <=  8'h62;        memory[39709] <=  8'h62;        memory[39710] <=  8'h72;        memory[39711] <=  8'h74;        memory[39712] <=  8'h62;        memory[39713] <=  8'h62;        memory[39714] <=  8'h61;        memory[39715] <=  8'h62;        memory[39716] <=  8'h72;        memory[39717] <=  8'h62;        memory[39718] <=  8'h74;        memory[39719] <=  8'h62;        memory[39720] <=  8'h62;        memory[39721] <=  8'h62;        memory[39722] <=  8'h63;        memory[39723] <=  8'h61;        memory[39724] <=  8'h72;        memory[39725] <=  8'h74;        memory[39726] <=  8'h73;        memory[39727] <=  8'h62;        memory[39728] <=  8'h61;        memory[39729] <=  8'h72;        memory[39730] <=  8'h74;        memory[39731] <=  8'h74;        memory[39732] <=  8'h62;        memory[39733] <=  8'h61;        memory[39734] <=  8'h72;        memory[39735] <=  8'h74;        memory[39736] <=  8'h78;        memory[39737] <=  8'h61;        memory[39738] <=  8'h74;        memory[39739] <=  8'h6b;        memory[39740] <=  8'h73;        memory[39741] <=  8'h68;        memory[39742] <=  8'h63;        memory[39743] <=  8'h66;        memory[39744] <=  8'h69;        memory[39745] <=  8'h77;        memory[39746] <=  8'h68;        memory[39747] <=  8'h61;        memory[39748] <=  8'h74;        memory[39749] <=  8'h61;        memory[39750] <=  8'h6e;        memory[39751] <=  8'h61;        memory[39752] <=  8'h62;        memory[39753] <=  8'h61;        memory[39754] <=  8'h63;        memory[39755] <=  8'h61;        memory[39756] <=  8'h74;        memory[39757] <=  8'h61;        memory[39758] <=  8'h62;        memory[39759] <=  8'h61;        memory[39760] <=  8'h72;        memory[39761] <=  8'h63;        memory[39762] <=  8'h61;        memory[39763] <=  8'h68;        memory[39764] <=  8'h64;        memory[39765] <=  8'h75;        memory[39766] <=  8'h63;        memory[39767] <=  8'h74;        memory[39768] <=  8'h61;        memory[39769] <=  8'h64;        memory[39770] <=  8'h61;        memory[39771] <=  8'h61;        memory[39772] <=  8'h63;        memory[39773] <=  8'h61;        memory[39774] <=  8'h72;        memory[39775] <=  8'h63;        memory[39776] <=  8'h74;        memory[39777] <=  8'h72;        memory[39778] <=  8'h63;        memory[39779] <=  8'h61;        memory[39780] <=  8'h74;        memory[39781] <=  8'h72;        memory[39782] <=  8'h63;        memory[39783] <=  8'h61;        memory[39784] <=  8'h74;        memory[39785] <=  8'h63;        memory[39786] <=  8'h62;        memory[39787] <=  8'h61;        memory[39788] <=  8'h74;        memory[39789] <=  8'h62;        memory[39790] <=  8'h72;        memory[39791] <=  8'h63;        memory[39792] <=  8'h61;        memory[39793] <=  8'h74;        memory[39794] <=  8'h72;        memory[39795] <=  8'h6e;        memory[39796] <=  8'h62;        memory[39797] <=  8'h61;        memory[39798] <=  8'h63;        memory[39799] <=  8'h61;        memory[39800] <=  8'h74;        memory[39801] <=  8'h79;        memory[39802] <=  8'h73;        memory[39803] <=  8'h6e;        memory[39804] <=  8'h63;        memory[39805] <=  8'h74;        memory[39806] <=  8'h61;        memory[39807] <=  8'h6e;        memory[39808] <=  8'h62;        memory[39809] <=  8'h61;        memory[39810] <=  8'h63;        memory[39811] <=  8'h72;        memory[39812] <=  8'h6e;        memory[39813] <=  8'h74;        memory[39814] <=  8'h61;        memory[39815] <=  8'h62;        memory[39816] <=  8'h74;        memory[39817] <=  8'h6e;        memory[39818] <=  8'h61;        memory[39819] <=  8'h72;        memory[39820] <=  8'h62;        memory[39821] <=  8'h78;        memory[39822] <=  8'h74;        memory[39823] <=  8'h61;        memory[39824] <=  8'h72;        memory[39825] <=  8'h62;        memory[39826] <=  8'h61;        memory[39827] <=  8'h72;        memory[39828] <=  8'h74;        memory[39829] <=  8'h74;        memory[39830] <=  8'h62;        memory[39831] <=  8'h61;        memory[39832] <=  8'h72;        memory[39833] <=  8'h74;        memory[39834] <=  8'h78;        memory[39835] <=  8'h61;        memory[39836] <=  8'h74;        memory[39837] <=  8'h6b;        memory[39838] <=  8'h73;        memory[39839] <=  8'h68;        memory[39840] <=  8'h63;        memory[39841] <=  8'h66;        memory[39842] <=  8'h69;        memory[39843] <=  8'h77;        memory[39844] <=  8'h68;        memory[39845] <=  8'h61;        memory[39846] <=  8'h74;        memory[39847] <=  8'h61;        memory[39848] <=  8'h6e;        memory[39849] <=  8'h61;        memory[39850] <=  8'h62;        memory[39851] <=  8'h61;        memory[39852] <=  8'h63;        memory[39853] <=  8'h61;        memory[39854] <=  8'h74;        memory[39855] <=  8'h61;        memory[39856] <=  8'h62;        memory[39857] <=  8'h61;        memory[39858] <=  8'h72;        memory[39859] <=  8'h63;        memory[39860] <=  8'h61;        memory[39861] <=  8'h68;        memory[39862] <=  8'h64;        memory[39863] <=  8'h75;        memory[39864] <=  8'h63;        memory[39865] <=  8'h74;        memory[39866] <=  8'h61;        memory[39867] <=  8'h64;        memory[39868] <=  8'h61;        memory[39869] <=  8'h61;        memory[39870] <=  8'h63;        memory[39871] <=  8'h61;        memory[39872] <=  8'h72;        memory[39873] <=  8'h63;        memory[39874] <=  8'h74;        memory[39875] <=  8'h72;        memory[39876] <=  8'h63;        memory[39877] <=  8'h61;        memory[39878] <=  8'h74;        memory[39879] <=  8'h72;        memory[39880] <=  8'h63;        memory[39881] <=  8'h61;        memory[39882] <=  8'h74;        memory[39883] <=  8'h63;        memory[39884] <=  8'h62;        memory[39885] <=  8'h61;        memory[39886] <=  8'h74;        memory[39887] <=  8'h62;        memory[39888] <=  8'h72;        memory[39889] <=  8'h63;        memory[39890] <=  8'h61;        memory[39891] <=  8'h74;        memory[39892] <=  8'h72;        memory[39893] <=  8'h6e;        memory[39894] <=  8'h62;        memory[39895] <=  8'h61;        memory[39896] <=  8'h63;        memory[39897] <=  8'h61;        memory[39898] <=  8'h74;        memory[39899] <=  8'h79;        memory[39900] <=  8'h73;        memory[39901] <=  8'h6e;        memory[39902] <=  8'h63;        memory[39903] <=  8'h74;        memory[39904] <=  8'h61;        memory[39905] <=  8'h6e;        memory[39906] <=  8'h62;        memory[39907] <=  8'h61;        memory[39908] <=  8'h63;        memory[39909] <=  8'h72;        memory[39910] <=  8'h6e;        memory[39911] <=  8'h74;        memory[39912] <=  8'h61;        memory[39913] <=  8'h62;        memory[39914] <=  8'h74;        memory[39915] <=  8'h6e;        memory[39916] <=  8'h61;        memory[39917] <=  8'h72;        memory[39918] <=  8'h62;        memory[39919] <=  8'h78;        memory[39920] <=  8'h74;        memory[39921] <=  8'h61;        memory[39922] <=  8'h72;        memory[39923] <=  8'h62;        memory[39924] <=  8'h61;        memory[39925] <=  8'h72;        memory[39926] <=  8'h74;        memory[39927] <=  8'h74;        memory[39928] <=  8'h62;        memory[39929] <=  8'h61;        memory[39930] <=  8'h72;        memory[39931] <=  8'h74;        memory[39932] <=  8'h78;        memory[39933] <=  8'h61;        memory[39934] <=  8'h74;        memory[39935] <=  8'h6b;        memory[39936] <=  8'h73;        memory[39937] <=  8'h68;        memory[39938] <=  8'h63;        memory[39939] <=  8'h66;        memory[39940] <=  8'h69;        memory[39941] <=  8'h77;        memory[39942] <=  8'h68;        memory[39943] <=  8'h61;        memory[39944] <=  8'h74;        memory[39945] <=  8'h61;        memory[39946] <=  8'h6e;        memory[39947] <=  8'h61;        memory[39948] <=  8'h62;        memory[39949] <=  8'h61;        memory[39950] <=  8'h63;        memory[39951] <=  8'h61;        memory[39952] <=  8'h74;        memory[39953] <=  8'h61;        memory[39954] <=  8'h62;        memory[39955] <=  8'h61;        memory[39956] <=  8'h72;        memory[39957] <=  8'h63;        memory[39958] <=  8'h61;        memory[39959] <=  8'h68;        memory[39960] <=  8'h64;        memory[39961] <=  8'h75;        memory[39962] <=  8'h63;        memory[39963] <=  8'h74;        memory[39964] <=  8'h61;        memory[39965] <=  8'h64;        memory[39966] <=  8'h61;        memory[39967] <=  8'h61;        memory[39968] <=  8'h63;        memory[39969] <=  8'h61;        memory[39970] <=  8'h72;        memory[39971] <=  8'h63;        memory[39972] <=  8'h74;        memory[39973] <=  8'h72;        memory[39974] <=  8'h63;        memory[39975] <=  8'h61;        memory[39976] <=  8'h74;        memory[39977] <=  8'h72;        memory[39978] <=  8'h63;        memory[39979] <=  8'h61;        memory[39980] <=  8'h74;        memory[39981] <=  8'h63;        memory[39982] <=  8'h62;        memory[39983] <=  8'h61;        memory[39984] <=  8'h74;        memory[39985] <=  8'h62;        memory[39986] <=  8'h72;        memory[39987] <=  8'h63;        memory[39988] <=  8'h61;        memory[39989] <=  8'h74;        memory[39990] <=  8'h72;        memory[39991] <=  8'h6e;        memory[39992] <=  8'h62;        memory[39993] <=  8'h61;        memory[39994] <=  8'h63;        memory[39995] <=  8'h61;        memory[39996] <=  8'h74;        memory[39997] <=  8'h79;        memory[39998] <=  8'h73;        memory[39999] <=  8'h6e;        memory[40000] <=  8'h63;        memory[40001] <=  8'h74;        memory[40002] <=  8'h61;        memory[40003] <=  8'h6e;        memory[40004] <=  8'h62;        memory[40005] <=  8'h61;        memory[40006] <=  8'h63;        memory[40007] <=  8'h72;        memory[40008] <=  8'h6e;        memory[40009] <=  8'h74;        memory[40010] <=  8'h61;        memory[40011] <=  8'h62;        memory[40012] <=  8'h74;        memory[40013] <=  8'h6e;        memory[40014] <=  8'h61;        memory[40015] <=  8'h72;        memory[40016] <=  8'h62;        memory[40017] <=  8'h78;        memory[40018] <=  8'h74;        memory[40019] <=  8'h61;        memory[40020] <=  8'h72;        memory[40021] <=  8'h5d;        memory[40022] <=  8'h5d;        memory[40023] <=  8'h65;        memory[40024] <=  8'h66;        memory[40025] <=  8'h77;        memory[40026] <=  8'h65;        memory[40027] <=  8'h5d;        memory[40028] <=  8'h65;        memory[40029] <=  8'h67;        memory[40030] <=  8'h73;        memory[40031] <=  8'h67;        memory[40032] <=  8'h66;        memory[40033] <=  8'h62;        memory[40034] <=  8'h61;        memory[40035] <=  8'h72;        memory[40036] <=  8'h74;        memory[40037] <=  8'h74;        memory[40038] <=  8'h62;        memory[40039] <=  8'h61;        memory[40040] <=  8'h72;        memory[40041] <=  8'h74;        memory[40042] <=  8'h78;        memory[40043] <=  8'h61;        memory[40044] <=  8'h74;        memory[40045] <=  8'h6b;        memory[40046] <=  8'h73;        memory[40047] <=  8'h68;        memory[40048] <=  8'h63;        memory[40049] <=  8'h66;        memory[40050] <=  8'h69;        memory[40051] <=  8'h77;        memory[40052] <=  8'h68;        memory[40053] <=  8'h61;        memory[40054] <=  8'h74;        memory[40055] <=  8'h61;        memory[40056] <=  8'h6e;        memory[40057] <=  8'h61;        memory[40058] <=  8'h62;        memory[40059] <=  8'h61;        memory[40060] <=  8'h63;        memory[40061] <=  8'h61;        memory[40062] <=  8'h74;        memory[40063] <=  8'h61;        memory[40064] <=  8'h62;        memory[40065] <=  8'h61;        memory[40066] <=  8'h72;        memory[40067] <=  8'h63;        memory[40068] <=  8'h61;        memory[40069] <=  8'h68;        memory[40070] <=  8'h64;        memory[40071] <=  8'h75;        memory[40072] <=  8'h63;        memory[40073] <=  8'h74;        memory[40074] <=  8'h61;        memory[40075] <=  8'h64;        memory[40076] <=  8'h61;        memory[40077] <=  8'h61;        memory[40078] <=  8'h63;        memory[40079] <=  8'h61;        memory[40080] <=  8'h72;        memory[40081] <=  8'h63;        memory[40082] <=  8'h74;        memory[40083] <=  8'h72;        memory[40084] <=  8'h63;        memory[40085] <=  8'h61;        memory[40086] <=  8'h74;        memory[40087] <=  8'h72;        memory[40088] <=  8'h63;        memory[40089] <=  8'h61;        memory[40090] <=  8'h74;        memory[40091] <=  8'h63;        memory[40092] <=  8'h62;        memory[40093] <=  8'h61;        memory[40094] <=  8'h74;        memory[40095] <=  8'h62;        memory[40096] <=  8'h72;        memory[40097] <=  8'h63;        memory[40098] <=  8'h61;        memory[40099] <=  8'h74;        memory[40100] <=  8'h72;        memory[40101] <=  8'h6e;        memory[40102] <=  8'h62;        memory[40103] <=  8'h61;        memory[40104] <=  8'h63;        memory[40105] <=  8'h61;        memory[40106] <=  8'h74;        memory[40107] <=  8'h79;        memory[40108] <=  8'h73;        memory[40109] <=  8'h6e;        memory[40110] <=  8'h63;        memory[40111] <=  8'h74;        memory[40112] <=  8'h61;        memory[40113] <=  8'h6e;        memory[40114] <=  8'h62;        memory[40115] <=  8'h61;        memory[40116] <=  8'h63;        memory[40117] <=  8'h72;        memory[40118] <=  8'h6e;        memory[40119] <=  8'h74;        memory[40120] <=  8'h61;        memory[40121] <=  8'h62;        memory[40122] <=  8'h74;        memory[40123] <=  8'h6e;        memory[40124] <=  8'h61;        memory[40125] <=  8'h72;        memory[40126] <=  8'h62;        memory[40127] <=  8'h78;        memory[40128] <=  8'h74;        memory[40129] <=  8'h61;        memory[40130] <=  8'h72;        memory[40131] <=  8'h62;        memory[40132] <=  8'h61;        memory[40133] <=  8'h72;        memory[40134] <=  8'h74;        memory[40135] <=  8'h74;        memory[40136] <=  8'h62;        memory[40137] <=  8'h61;        memory[40138] <=  8'h72;        memory[40139] <=  8'h74;        memory[40140] <=  8'h78;        memory[40141] <=  8'h61;        memory[40142] <=  8'h74;        memory[40143] <=  8'h6b;        memory[40144] <=  8'h73;        memory[40145] <=  8'h68;        memory[40146] <=  8'h63;        memory[40147] <=  8'h66;        memory[40148] <=  8'h69;        memory[40149] <=  8'h77;        memory[40150] <=  8'h68;        memory[40151] <=  8'h61;        memory[40152] <=  8'h74;        memory[40153] <=  8'h61;        memory[40154] <=  8'h6e;        memory[40155] <=  8'h61;        memory[40156] <=  8'h62;        memory[40157] <=  8'h61;        memory[40158] <=  8'h63;        memory[40159] <=  8'h61;        memory[40160] <=  8'h74;        memory[40161] <=  8'h61;        memory[40162] <=  8'h62;        memory[40163] <=  8'h61;        memory[40164] <=  8'h72;        memory[40165] <=  8'h63;        memory[40166] <=  8'h61;        memory[40167] <=  8'h68;        memory[40168] <=  8'h64;        memory[40169] <=  8'h75;        memory[40170] <=  8'h63;        memory[40171] <=  8'h74;        memory[40172] <=  8'h61;        memory[40173] <=  8'h64;        memory[40174] <=  8'h61;        memory[40175] <=  8'h61;        memory[40176] <=  8'h63;        memory[40177] <=  8'h61;        memory[40178] <=  8'h72;        memory[40179] <=  8'h63;        memory[40180] <=  8'h74;        memory[40181] <=  8'h72;        memory[40182] <=  8'h63;        memory[40183] <=  8'h61;        memory[40184] <=  8'h74;        memory[40185] <=  8'h72;        memory[40186] <=  8'h63;        memory[40187] <=  8'h61;        memory[40188] <=  8'h74;        memory[40189] <=  8'h63;        memory[40190] <=  8'h62;        memory[40191] <=  8'h61;        memory[40192] <=  8'h74;        memory[40193] <=  8'h62;        memory[40194] <=  8'h72;        memory[40195] <=  8'h63;        memory[40196] <=  8'h61;        memory[40197] <=  8'h74;        memory[40198] <=  8'h72;        memory[40199] <=  8'h6e;        memory[40200] <=  8'h62;        memory[40201] <=  8'h61;        memory[40202] <=  8'h63;        memory[40203] <=  8'h61;        memory[40204] <=  8'h74;        memory[40205] <=  8'h79;        memory[40206] <=  8'h73;        memory[40207] <=  8'h6e;        memory[40208] <=  8'h63;        memory[40209] <=  8'h74;        memory[40210] <=  8'h61;        memory[40211] <=  8'h6e;        memory[40212] <=  8'h62;        memory[40213] <=  8'h61;        memory[40214] <=  8'h63;        memory[40215] <=  8'h72;        memory[40216] <=  8'h6e;        memory[40217] <=  8'h74;        memory[40218] <=  8'h61;        memory[40219] <=  8'h62;        memory[40220] <=  8'h74;        memory[40221] <=  8'h6e;        memory[40222] <=  8'h61;        memory[40223] <=  8'h72;        memory[40224] <=  8'h62;        memory[40225] <=  8'h78;        memory[40226] <=  8'h74;        memory[40227] <=  8'h61;        memory[40228] <=  8'h72;        memory[40229] <=  8'h64;        memory[40230] <=  8'h66;        memory[40231] <=  8'h73;        memory[40232] <=  8'h67;        memory[40233] <=  8'h76;        memory[40234] <=  8'h68;        memory[40235] <=  8'h62;        memory[40236] <=  8'h6b;        memory[40237] <=  8'h6a;        memory[40238] <=  8'h6e;        memory[40239] <=  8'h6d;        memory[40240] <=  8'h62;        memory[40241] <=  8'h76;        memory[40242] <=  8'h78;        memory[40243] <=  8'h63;        memory[40244] <=  8'h73;        memory[40245] <=  8'h66;        memory[40246] <=  8'h72;        memory[40247] <=  8'h74;        memory[40248] <=  8'h79;        memory[40249] <=  8'h75;        memory[40250] <=  8'h6a;        memory[40251] <=  8'h6e;        memory[40252] <=  8'h62;        memory[40253] <=  8'h76;        memory[40254] <=  8'h63;        memory[40255] <=  8'h64;        memory[40256] <=  8'h74;        memory[40257] <=  8'h79;        memory[40258] <=  8'h75;        memory[40259] <=  8'h69;        memory[40260] <=  8'h6b;        memory[40261] <=  8'h6d;        memory[40262] <=  8'h6e;        memory[40263] <=  8'h62;        memory[40264] <=  8'h76;        memory[40265] <=  8'h63;        memory[40266] <=  8'h78;        memory[40267] <=  8'h73;        memory[40268] <=  8'h64;        memory[40269] <=  8'h72;        memory[40270] <=  8'h74;        memory[40271] <=  8'h79;        memory[40272] <=  8'h75;        memory[40273] <=  8'h69;        memory[40274] <=  8'h6b;        memory[40275] <=  8'h6d;        memory[40276] <=  8'h6e;        memory[40277] <=  8'h62;        memory[40278] <=  8'h76;        memory[40279] <=  8'h63;        memory[40280] <=  8'h73;        memory[40281] <=  8'h77;        memory[40282] <=  8'h33;        memory[40283] <=  8'h34;        memory[40284] <=  8'h35;        memory[40285] <=  8'h36;        memory[40286] <=  8'h37;        memory[40287] <=  8'h38;        memory[40288] <=  8'h69;        memory[40289] <=  8'h6b;        memory[40290] <=  8'h6d;        memory[40291] <=  8'h6e;        memory[40292] <=  8'h62;        memory[40293] <=  8'h76;        memory[40294] <=  8'h63;        memory[40295] <=  8'h64;        memory[40296] <=  8'h65;        memory[40297] <=  8'h72;        memory[40298] <=  8'h36;        memory[40299] <=  8'h37;        memory[40300] <=  8'h38;        memory[40301] <=  8'h69;        memory[40302] <=  8'h6f;        memory[40303] <=  8'h6b;        memory[40304] <=  8'h6a;        memory[40305] <=  8'h6e;        memory[40306] <=  8'h62;        memory[40307] <=  8'h76;        memory[40308] <=  8'h63;        memory[40309] <=  8'h64;        memory[40310] <=  8'h72;        memory[40311] <=  8'h74;        memory[40312] <=  8'h79;        memory[40313] <=  8'h75;        memory[40314] <=  8'h73;        memory[40315] <=  8'h6a;        memory[40316] <=  8'h63;        memory[40317] <=  8'h6e;        memory[40318] <=  8'h62;        memory[40319] <=  8'h64;        memory[40320] <=  8'h66;        memory[40321] <=  8'h73;        memory[40322] <=  8'h74;        memory[40323] <=  8'h79;        memory[40324] <=  8'h75;        memory[40325] <=  8'h61;        memory[40326] <=  8'h69;        memory[40327] <=  8'h6b;        memory[40328] <=  8'h78;        memory[40329] <=  8'h6d;        memory[40330] <=  8'h6e;        memory[40331] <=  8'h73;        memory[40332] <=  8'h6a;        memory[40333] <=  8'h6f;        memory[40334] <=  8'h64;        memory[40335] <=  8'h6c;        memory[40336] <=  8'h63;        memory[40337] <=  8'h78;        memory[40338] <=  8'h62;        memory[40339] <=  8'h61;        memory[40340] <=  8'h72;        memory[40341] <=  8'h74;        memory[40342] <=  8'h78;        memory[40343] <=  8'h61;        memory[40344] <=  8'h74;        memory[40345] <=  8'h6b;        memory[40346] <=  8'h73;        memory[40347] <=  8'h68;        memory[40348] <=  8'h63;        memory[40349] <=  8'h66;        memory[40350] <=  8'h69;        memory[40351] <=  8'h77;        memory[40352] <=  8'h68;        memory[40353] <=  8'h61;        memory[40354] <=  8'h74;        memory[40355] <=  8'h61;        memory[40356] <=  8'h6e;        memory[40357] <=  8'h61;        memory[40358] <=  8'h62;        memory[40359] <=  8'h61;        memory[40360] <=  8'h63;        memory[40361] <=  8'h61;        memory[40362] <=  8'h74;        memory[40363] <=  8'h61;        memory[40364] <=  8'h62;        memory[40365] <=  8'h61;        memory[40366] <=  8'h72;        memory[40367] <=  8'h63;        memory[40368] <=  8'h61;        memory[40369] <=  8'h68;        memory[40370] <=  8'h64;        memory[40371] <=  8'h75;        memory[40372] <=  8'h63;        memory[40373] <=  8'h74;        memory[40374] <=  8'h61;        memory[40375] <=  8'h64;        memory[40376] <=  8'h61;        memory[40377] <=  8'h61;        memory[40378] <=  8'h63;        memory[40379] <=  8'h61;        memory[40380] <=  8'h72;        memory[40381] <=  8'h62;        memory[40382] <=  8'h61;        memory[40383] <=  8'h72;        memory[40384] <=  8'h74;        memory[40385] <=  8'h78;        memory[40386] <=  8'h61;        memory[40387] <=  8'h74;        memory[40388] <=  8'h6b;        memory[40389] <=  8'h73;        memory[40390] <=  8'h68;        memory[40391] <=  8'h63;        memory[40392] <=  8'h66;        memory[40393] <=  8'h69;        memory[40394] <=  8'h77;        memory[40395] <=  8'h68;        memory[40396] <=  8'h61;        memory[40397] <=  8'h74;        memory[40398] <=  8'h61;        memory[40399] <=  8'h6e;        memory[40400] <=  8'h61;        memory[40401] <=  8'h62;        memory[40402] <=  8'h61;        memory[40403] <=  8'h63;        memory[40404] <=  8'h61;        memory[40405] <=  8'h74;        memory[40406] <=  8'h61;        memory[40407] <=  8'h62;        memory[40408] <=  8'h61;        memory[40409] <=  8'h72;        memory[40410] <=  8'h63;        memory[40411] <=  8'h61;        memory[40412] <=  8'h68;        memory[40413] <=  8'h64;        memory[40414] <=  8'h75;        memory[40415] <=  8'h63;        memory[40416] <=  8'h74;        memory[40417] <=  8'h61;        memory[40418] <=  8'h64;        memory[40419] <=  8'h61;        memory[40420] <=  8'h61;        memory[40421] <=  8'h63;        memory[40422] <=  8'h61;        memory[40423] <=  8'h72;        memory[40424] <=  8'h62;        memory[40425] <=  8'h61;        memory[40426] <=  8'h72;        memory[40427] <=  8'h74;        memory[40428] <=  8'h78;        memory[40429] <=  8'h61;        memory[40430] <=  8'h74;        memory[40431] <=  8'h6b;        memory[40432] <=  8'h73;        memory[40433] <=  8'h68;        memory[40434] <=  8'h63;        memory[40435] <=  8'h66;        memory[40436] <=  8'h69;        memory[40437] <=  8'h77;        memory[40438] <=  8'h68;        memory[40439] <=  8'h61;        memory[40440] <=  8'h74;        memory[40441] <=  8'h61;        memory[40442] <=  8'h6e;        memory[40443] <=  8'h61;        memory[40444] <=  8'h62;        memory[40445] <=  8'h61;        memory[40446] <=  8'h63;        memory[40447] <=  8'h61;        memory[40448] <=  8'h74;        memory[40449] <=  8'h61;        memory[40450] <=  8'h62;        memory[40451] <=  8'h61;        memory[40452] <=  8'h72;        memory[40453] <=  8'h63;        memory[40454] <=  8'h61;        memory[40455] <=  8'h68;        memory[40456] <=  8'h64;        memory[40457] <=  8'h75;        memory[40458] <=  8'h63;        memory[40459] <=  8'h74;        memory[40460] <=  8'h61;        memory[40461] <=  8'h64;        memory[40462] <=  8'h61;        memory[40463] <=  8'h61;        memory[40464] <=  8'h63;        memory[40465] <=  8'h61;        memory[40466] <=  8'h72;        memory[40467] <=  8'h62;        memory[40468] <=  8'h61;        memory[40469] <=  8'h72;        memory[40470] <=  8'h74;        memory[40471] <=  8'h78;        memory[40472] <=  8'h61;        memory[40473] <=  8'h74;        memory[40474] <=  8'h6b;        memory[40475] <=  8'h73;        memory[40476] <=  8'h68;        memory[40477] <=  8'h63;        memory[40478] <=  8'h66;        memory[40479] <=  8'h69;        memory[40480] <=  8'h77;        memory[40481] <=  8'h68;        memory[40482] <=  8'h61;        memory[40483] <=  8'h74;        memory[40484] <=  8'h61;        memory[40485] <=  8'h6e;        memory[40486] <=  8'h61;        memory[40487] <=  8'h62;        memory[40488] <=  8'h61;        memory[40489] <=  8'h63;        memory[40490] <=  8'h61;        memory[40491] <=  8'h74;        memory[40492] <=  8'h61;        memory[40493] <=  8'h62;        memory[40494] <=  8'h61;        memory[40495] <=  8'h72;        memory[40496] <=  8'h63;        memory[40497] <=  8'h61;        memory[40498] <=  8'h68;        memory[40499] <=  8'h64;        memory[40500] <=  8'h75;        memory[40501] <=  8'h63;        memory[40502] <=  8'h74;        memory[40503] <=  8'h61;        memory[40504] <=  8'h64;        memory[40505] <=  8'h61;        memory[40506] <=  8'h61;        memory[40507] <=  8'h63;        memory[40508] <=  8'h61;        memory[40509] <=  8'h72;        memory[40510] <=  8'h62;        memory[40511] <=  8'h61;        memory[40512] <=  8'h72;        memory[40513] <=  8'h74;        memory[40514] <=  8'h78;        memory[40515] <=  8'h61;        memory[40516] <=  8'h74;        memory[40517] <=  8'h6b;        memory[40518] <=  8'h73;        memory[40519] <=  8'h68;        memory[40520] <=  8'h63;        memory[40521] <=  8'h66;        memory[40522] <=  8'h69;        memory[40523] <=  8'h77;        memory[40524] <=  8'h68;        memory[40525] <=  8'h61;        memory[40526] <=  8'h74;        memory[40527] <=  8'h61;        memory[40528] <=  8'h6e;        memory[40529] <=  8'h61;        memory[40530] <=  8'h62;        memory[40531] <=  8'h61;        memory[40532] <=  8'h63;        memory[40533] <=  8'h61;        memory[40534] <=  8'h74;        memory[40535] <=  8'h61;        memory[40536] <=  8'h62;        memory[40537] <=  8'h61;        memory[40538] <=  8'h72;        memory[40539] <=  8'h63;        memory[40540] <=  8'h61;        memory[40541] <=  8'h68;        memory[40542] <=  8'h64;        memory[40543] <=  8'h75;        memory[40544] <=  8'h63;        memory[40545] <=  8'h74;        memory[40546] <=  8'h61;        memory[40547] <=  8'h64;        memory[40548] <=  8'h61;        memory[40549] <=  8'h61;        memory[40550] <=  8'h63;        memory[40551] <=  8'h61;        memory[40552] <=  8'h72;        memory[40553] <=  8'h62;        memory[40554] <=  8'h61;        memory[40555] <=  8'h72;        memory[40556] <=  8'h74;        memory[40557] <=  8'h78;        memory[40558] <=  8'h61;        memory[40559] <=  8'h74;        memory[40560] <=  8'h6b;        memory[40561] <=  8'h73;        memory[40562] <=  8'h68;        memory[40563] <=  8'h63;        memory[40564] <=  8'h66;        memory[40565] <=  8'h69;        memory[40566] <=  8'h77;        memory[40567] <=  8'h68;        memory[40568] <=  8'h61;        memory[40569] <=  8'h74;        memory[40570] <=  8'h61;        memory[40571] <=  8'h6e;        memory[40572] <=  8'h61;        memory[40573] <=  8'h62;        memory[40574] <=  8'h61;        memory[40575] <=  8'h63;        memory[40576] <=  8'h61;        memory[40577] <=  8'h74;        memory[40578] <=  8'h61;        memory[40579] <=  8'h62;        memory[40580] <=  8'h61;        memory[40581] <=  8'h72;        memory[40582] <=  8'h63;        memory[40583] <=  8'h61;        memory[40584] <=  8'h68;        memory[40585] <=  8'h64;        memory[40586] <=  8'h75;        memory[40587] <=  8'h63;        memory[40588] <=  8'h74;        memory[40589] <=  8'h61;        memory[40590] <=  8'h64;        memory[40591] <=  8'h61;        memory[40592] <=  8'h61;        memory[40593] <=  8'h63;        memory[40594] <=  8'h61;        memory[40595] <=  8'h72;        memory[40596] <=  8'h62;        memory[40597] <=  8'h61;        memory[40598] <=  8'h72;        memory[40599] <=  8'h74;        memory[40600] <=  8'h78;        memory[40601] <=  8'h61;        memory[40602] <=  8'h74;        memory[40603] <=  8'h6b;        memory[40604] <=  8'h73;        memory[40605] <=  8'h68;        memory[40606] <=  8'h63;        memory[40607] <=  8'h66;        memory[40608] <=  8'h69;        memory[40609] <=  8'h77;        memory[40610] <=  8'h68;        memory[40611] <=  8'h61;        memory[40612] <=  8'h74;        memory[40613] <=  8'h61;        memory[40614] <=  8'h6e;        memory[40615] <=  8'h61;        memory[40616] <=  8'h62;        memory[40617] <=  8'h61;        memory[40618] <=  8'h63;        memory[40619] <=  8'h61;        memory[40620] <=  8'h74;        memory[40621] <=  8'h61;        memory[40622] <=  8'h62;        memory[40623] <=  8'h61;        memory[40624] <=  8'h72;        memory[40625] <=  8'h63;        memory[40626] <=  8'h61;        memory[40627] <=  8'h68;        memory[40628] <=  8'h64;        memory[40629] <=  8'h75;        memory[40630] <=  8'h63;        memory[40631] <=  8'h74;        memory[40632] <=  8'h61;        memory[40633] <=  8'h64;        memory[40634] <=  8'h61;        memory[40635] <=  8'h61;        memory[40636] <=  8'h63;        memory[40637] <=  8'h61;        memory[40638] <=  8'h72;        memory[40639] <=  8'h62;        memory[40640] <=  8'h61;        memory[40641] <=  8'h72;        memory[40642] <=  8'h74;        memory[40643] <=  8'h78;        memory[40644] <=  8'h61;        memory[40645] <=  8'h74;        memory[40646] <=  8'h6b;        memory[40647] <=  8'h73;        memory[40648] <=  8'h68;        memory[40649] <=  8'h63;        memory[40650] <=  8'h66;        memory[40651] <=  8'h69;        memory[40652] <=  8'h77;        memory[40653] <=  8'h68;        memory[40654] <=  8'h61;        memory[40655] <=  8'h74;        memory[40656] <=  8'h61;        memory[40657] <=  8'h6e;        memory[40658] <=  8'h61;        memory[40659] <=  8'h62;        memory[40660] <=  8'h61;        memory[40661] <=  8'h63;        memory[40662] <=  8'h61;        memory[40663] <=  8'h74;        memory[40664] <=  8'h61;        memory[40665] <=  8'h62;        memory[40666] <=  8'h61;        memory[40667] <=  8'h72;        memory[40668] <=  8'h63;        memory[40669] <=  8'h61;        memory[40670] <=  8'h68;        memory[40671] <=  8'h64;        memory[40672] <=  8'h75;        memory[40673] <=  8'h63;        memory[40674] <=  8'h74;        memory[40675] <=  8'h61;        memory[40676] <=  8'h64;        memory[40677] <=  8'h61;        memory[40678] <=  8'h61;        memory[40679] <=  8'h63;        memory[40680] <=  8'h61;        memory[40681] <=  8'h72;        memory[40682] <=  8'h62;        memory[40683] <=  8'h61;        memory[40684] <=  8'h72;        memory[40685] <=  8'h74;        memory[40686] <=  8'h78;        memory[40687] <=  8'h61;        memory[40688] <=  8'h74;        memory[40689] <=  8'h6b;        memory[40690] <=  8'h73;        memory[40691] <=  8'h68;        memory[40692] <=  8'h63;        memory[40693] <=  8'h66;        memory[40694] <=  8'h69;        memory[40695] <=  8'h77;        memory[40696] <=  8'h68;        memory[40697] <=  8'h61;        memory[40698] <=  8'h74;        memory[40699] <=  8'h61;        memory[40700] <=  8'h6e;        memory[40701] <=  8'h61;        memory[40702] <=  8'h62;        memory[40703] <=  8'h61;        memory[40704] <=  8'h63;        memory[40705] <=  8'h61;        memory[40706] <=  8'h74;        memory[40707] <=  8'h61;        memory[40708] <=  8'h62;        memory[40709] <=  8'h61;        memory[40710] <=  8'h72;        memory[40711] <=  8'h63;        memory[40712] <=  8'h61;        memory[40713] <=  8'h68;        memory[40714] <=  8'h64;        memory[40715] <=  8'h75;        memory[40716] <=  8'h63;        memory[40717] <=  8'h74;        memory[40718] <=  8'h61;        memory[40719] <=  8'h64;        memory[40720] <=  8'h61;        memory[40721] <=  8'h61;        memory[40722] <=  8'h63;        memory[40723] <=  8'h61;        memory[40724] <=  8'h72;        memory[40725] <=  8'h62;        memory[40726] <=  8'h61;        memory[40727] <=  8'h72;        memory[40728] <=  8'h74;        memory[40729] <=  8'h74;        memory[40730] <=  8'h62;        memory[40731] <=  8'h61;        memory[40732] <=  8'h72;        memory[40733] <=  8'h74;        memory[40734] <=  8'h78;        memory[40735] <=  8'h61;        memory[40736] <=  8'h74;        memory[40737] <=  8'h6b;        memory[40738] <=  8'h73;        memory[40739] <=  8'h68;        memory[40740] <=  8'h63;        memory[40741] <=  8'h66;        memory[40742] <=  8'h69;        memory[40743] <=  8'h77;        memory[40744] <=  8'h68;        memory[40745] <=  8'h61;        memory[40746] <=  8'h74;        memory[40747] <=  8'h61;        memory[40748] <=  8'h6e;        memory[40749] <=  8'h61;        memory[40750] <=  8'h62;        memory[40751] <=  8'h61;        memory[40752] <=  8'h63;        memory[40753] <=  8'h61;        memory[40754] <=  8'h74;        memory[40755] <=  8'h61;        memory[40756] <=  8'h62;        memory[40757] <=  8'h61;        memory[40758] <=  8'h72;        memory[40759] <=  8'h63;        memory[40760] <=  8'h61;        memory[40761] <=  8'h68;        memory[40762] <=  8'h64;        memory[40763] <=  8'h75;        memory[40764] <=  8'h63;        memory[40765] <=  8'h74;        memory[40766] <=  8'h61;        memory[40767] <=  8'h64;        memory[40768] <=  8'h61;        memory[40769] <=  8'h61;        memory[40770] <=  8'h63;        memory[40771] <=  8'h61;        memory[40772] <=  8'h72;        memory[40773] <=  8'h63;        memory[40774] <=  8'h74;        memory[40775] <=  8'h72;        memory[40776] <=  8'h63;        memory[40777] <=  8'h61;        memory[40778] <=  8'h74;        memory[40779] <=  8'h72;        memory[40780] <=  8'h63;        memory[40781] <=  8'h61;        memory[40782] <=  8'h74;        memory[40783] <=  8'h63;        memory[40784] <=  8'h62;        memory[40785] <=  8'h61;        memory[40786] <=  8'h74;        memory[40787] <=  8'h62;        memory[40788] <=  8'h72;        memory[40789] <=  8'h63;        memory[40790] <=  8'h61;        memory[40791] <=  8'h72;        memory[40792] <=  8'h62;        memory[40793] <=  8'h78;        memory[40794] <=  8'h74;        memory[40795] <=  8'h61;        memory[40796] <=  8'h72;        memory[40797] <=  8'h64;        memory[40798] <=  8'h66;        memory[40799] <=  8'h73;        memory[40800] <=  8'h67;        memory[40801] <=  8'h76;        memory[40802] <=  8'h68;        memory[40803] <=  8'h62;        memory[40804] <=  8'h6b;        memory[40805] <=  8'h6a;        memory[40806] <=  8'h6e;        memory[40807] <=  8'h6d;        memory[40808] <=  8'h62;        memory[40809] <=  8'h76;        memory[40810] <=  8'h78;        memory[40811] <=  8'h63;        memory[40812] <=  8'h73;        memory[40813] <=  8'h66;        memory[40814] <=  8'h72;        memory[40815] <=  8'h74;        memory[40816] <=  8'h79;        memory[40817] <=  8'h75;        memory[40818] <=  8'h6a;        memory[40819] <=  8'h6e;        memory[40820] <=  8'h62;        memory[40821] <=  8'h76;        memory[40822] <=  8'h63;        memory[40823] <=  8'h64;        memory[40824] <=  8'h74;        memory[40825] <=  8'h79;        memory[40826] <=  8'h75;        memory[40827] <=  8'h69;        memory[40828] <=  8'h6b;        memory[40829] <=  8'h6d;        memory[40830] <=  8'h6e;        memory[40831] <=  8'h62;        memory[40832] <=  8'h76;        memory[40833] <=  8'h63;        memory[40834] <=  8'h78;        memory[40835] <=  8'h73;        memory[40836] <=  8'h64;        memory[40837] <=  8'h72;        memory[40838] <=  8'h74;        memory[40839] <=  8'h79;        memory[40840] <=  8'h75;        memory[40841] <=  8'h69;        memory[40842] <=  8'h6b;        memory[40843] <=  8'h6d;        memory[40844] <=  8'h6e;        memory[40845] <=  8'h62;        memory[40846] <=  8'h76;        memory[40847] <=  8'h63;        memory[40848] <=  8'h73;        memory[40849] <=  8'h77;        memory[40850] <=  8'h33;        memory[40851] <=  8'h34;        memory[40852] <=  8'h35;        memory[40853] <=  8'h36;        memory[40854] <=  8'h37;        memory[40855] <=  8'h38;        memory[40856] <=  8'h69;        memory[40857] <=  8'h6b;        memory[40858] <=  8'h6d;        memory[40859] <=  8'h6e;        memory[40860] <=  8'h62;        memory[40861] <=  8'h76;        memory[40862] <=  8'h63;        memory[40863] <=  8'h64;        memory[40864] <=  8'h65;        memory[40865] <=  8'h72;        memory[40866] <=  8'h36;        memory[40867] <=  8'h37;        memory[40868] <=  8'h38;        memory[40869] <=  8'h69;        memory[40870] <=  8'h6f;        memory[40871] <=  8'h6b;        memory[40872] <=  8'h6a;        memory[40873] <=  8'h6e;        memory[40874] <=  8'h62;        memory[40875] <=  8'h76;        memory[40876] <=  8'h63;        memory[40877] <=  8'h64;        memory[40878] <=  8'h72;        memory[40879] <=  8'h74;        memory[40880] <=  8'h79;        memory[40881] <=  8'h75;        memory[40882] <=  8'h73;        memory[40883] <=  8'h6a;        memory[40884] <=  8'h63;        memory[40885] <=  8'h6e;        memory[40886] <=  8'h62;        memory[40887] <=  8'h64;        memory[40888] <=  8'h66;        memory[40889] <=  8'h73;        memory[40890] <=  8'h74;        memory[40891] <=  8'h79;        memory[40892] <=  8'h75;        memory[40893] <=  8'h61;        memory[40894] <=  8'h69;        memory[40895] <=  8'h6b;        memory[40896] <=  8'h78;        memory[40897] <=  8'h6d;        memory[40898] <=  8'h6e;        memory[40899] <=  8'h73;        memory[40900] <=  8'h6a;        memory[40901] <=  8'h6f;        memory[40902] <=  8'h64;        memory[40903] <=  8'h6c;        memory[40904] <=  8'h63;        memory[40905] <=  8'h78;        memory[40906] <=  8'h2c;        memory[40907] <=  8'h6d;        memory[40908] <=  8'h73;        memory[40909] <=  8'h6b;        memory[40910] <=  8'h64;        memory[40911] <=  8'h6c;        memory[40912] <=  8'h70;        memory[40913] <=  8'h5b;        memory[40914] <=  8'h3b;        memory[40915] <=  8'h73;        memory[40916] <=  8'h6c;        memory[40917] <=  8'h64;        memory[40918] <=  8'h70;        memory[40919] <=  8'h76;        memory[40920] <=  8'h63;        memory[40921] <=  8'h5b;        memory[40922] <=  8'h78;        memory[40923] <=  8'h76;        memory[40924] <=  8'h63;        memory[40925] <=  8'h5b;        memory[40926] <=  8'h78;        memory[40927] <=  8'h70;        memory[40928] <=  8'h6f;        memory[40929] <=  8'h20;        memory[40930] <=  8'h62;        memory[40931] <=  8'h61;        memory[40932] <=  8'h72;        memory[40933] <=  8'h74;        memory[40934] <=  8'h74;        memory[40935] <=  8'h62;        memory[40936] <=  8'h61;        memory[40937] <=  8'h72;        memory[40938] <=  8'h74;        memory[40939] <=  8'h78;        memory[40940] <=  8'h61;        memory[40941] <=  8'h74;        memory[40942] <=  8'h6b;        memory[40943] <=  8'h73;        memory[40944] <=  8'h68;        memory[40945] <=  8'h63;        memory[40946] <=  8'h66;        memory[40947] <=  8'h69;        memory[40948] <=  8'h77;        memory[40949] <=  8'h68;        memory[40950] <=  8'h61;        memory[40951] <=  8'h69;        memory[40952] <=  8'h6a;        memory[40953] <=  8'h78;        memory[40954] <=  8'h5d;        memory[40955] <=  8'h65;        memory[40956] <=  8'h6b;        memory[40957] <=  8'h6f;        memory[40958] <=  8'h39;        memory[40959] <=  8'h64;        memory[40960] <=  8'h75;        memory[40961] <=  8'h38;        memory[40962] <=  8'h79;        memory[40963] <=  8'h20;        memory[40964] <=  8'h37;        memory[40965] <=  8'h63;        memory[40966] <=  8'h67;        memory[40967] <=  8'h78;        memory[40968] <=  8'h63;        memory[40969] <=  8'h75;        memory[40970] <=  8'h68;        memory[40971] <=  8'h69;        memory[40972] <=  8'h6a;        memory[40973] <=  8'h77;        memory[40974] <=  8'h69;        memory[40975] <=  8'h64;        memory[40976] <=  8'h66;        memory[40977] <=  8'h68;        memory[40978] <=  8'h75;        memory[40979] <=  8'h76;        memory[40980] <=  8'h64;        memory[40981] <=  8'h62;        memory[40982] <=  8'h66;        memory[40983] <=  8'h6a;        memory[40984] <=  8'h6e;        memory[40985] <=  8'h6b;        memory[40986] <=  8'h6a;        memory[40987] <=  8'h65;        memory[40988] <=  8'h38;        memory[40989] <=  8'h66;        memory[40990] <=  8'h37;        memory[40991] <=  8'h67;        memory[40992] <=  8'h79;        memory[40993] <=  8'h76;        memory[40994] <=  8'h63;        memory[40995] <=  8'h68;        memory[40996] <=  8'h69;        memory[40997] <=  8'h6a;        memory[40998] <=  8'h33;        memory[40999] <=  8'h65;        memory[41000] <=  8'h67;        memory[41001] <=  8'h79;        memory[41002] <=  8'h72;        memory[41003] <=  8'h64;        memory[41004] <=  8'h62;        memory[41005] <=  8'h6e;        memory[41006] <=  8'h63;        memory[41007] <=  8'h7a;        memory[41008] <=  8'h6a;        memory[41009] <=  8'h6f;        memory[41010] <=  8'h66;        memory[41011] <=  8'h78;        memory[41012] <=  8'h6a;        memory[41013] <=  8'h69;        memory[41014] <=  8'h63;        memory[41015] <=  8'h68;        memory[41016] <=  8'h62;        memory[41017] <=  8'h6e;        memory[41018] <=  8'h6d;        memory[41019] <=  8'h63;        memory[41020] <=  8'h73;        memory[41021] <=  8'h6c;        memory[41022] <=  8'h6b;        memory[41023] <=  8'h6a;        memory[41024] <=  8'h69;        memory[41025] <=  8'h68;        memory[41026] <=  8'h76;        memory[41027] <=  8'h75;        memory[41028] <=  8'h69;        memory[41029] <=  8'h64;        memory[41030] <=  8'h68;        memory[41031] <=  8'h75;        memory[41032] <=  8'h67;        memory[41033] <=  8'h79;        memory[41034] <=  8'h62;        memory[41035] <=  8'h68;        memory[41036] <=  8'h65;        memory[41037] <=  8'h6a;        memory[41038] <=  8'h72;        memory[41039] <=  8'h6b;        memory[41040] <=  8'h6a;        memory[41041] <=  8'h6f;        memory[41042] <=  8'h64;        memory[41043] <=  8'h67;        memory[41044] <=  8'h69;        memory[41045] <=  8'h75;        memory[41046] <=  8'h69;        memory[41047] <=  8'h67;        memory[41048] <=  8'h76;        memory[41049] <=  8'h79;        memory[41050] <=  8'h75;        memory[41051] <=  8'h67;        memory[41052] <=  8'h78;        memory[41053] <=  8'h68;        memory[41054] <=  8'h63;        memory[41055] <=  8'h20;        memory[41056] <=  8'h20;        memory[41057] <=  8'h20;        memory[41058] <=  8'h78;        memory[41059] <=  8'h76;        memory[41060] <=  8'h20;        memory[41061] <=  8'h63;        memory[41062] <=  8'h78;        memory[41063] <=  8'h67;        memory[41064] <=  8'h79;        memory[41065] <=  8'h63;        memory[41066] <=  8'h75;        memory[41067] <=  8'h68;        memory[41068] <=  8'h6a;        memory[41069] <=  8'h6b;        memory[41070] <=  8'h61;        memory[41071] <=  8'h6c;        memory[41072] <=  8'h78;        memory[41073] <=  8'h76;        memory[41074] <=  8'h70;        memory[41075] <=  8'h6f;        memory[41076] <=  8'h69;        memory[41077] <=  8'h6a;        memory[41078] <=  8'h69;        memory[41079] <=  8'h68;        memory[41080] <=  8'h6a;        memory[41081] <=  8'h62;        memory[41082] <=  8'h77;        memory[41083] <=  8'h65;        memory[41084] <=  8'h6e;        memory[41085] <=  8'h61;        memory[41086] <=  8'h66;        memory[41087] <=  8'h6d;        memory[41088] <=  8'h64;        memory[41089] <=  8'h6b;        memory[41090] <=  8'h6d;        memory[41091] <=  8'h76;        memory[41092] <=  8'h6c;        memory[41093] <=  8'h63;        memory[41094] <=  8'h6f;        memory[41095] <=  8'h64;        memory[41096] <=  8'h69;        memory[41097] <=  8'h75;        memory[41098] <=  8'h68;        memory[41099] <=  8'h73;        memory[41100] <=  8'h66;        memory[41101] <=  8'h65;        memory[41102] <=  8'h62;        memory[41103] <=  8'h6e;        memory[41104] <=  8'h64;        memory[41105] <=  8'h73;        memory[41106] <=  8'h63;        memory[41107] <=  8'h6b;        memory[41108] <=  8'h20;        memory[41109] <=  8'h78;        memory[41110] <=  8'h6a;        memory[41111] <=  8'h78;        memory[41112] <=  8'h63;        memory[41113] <=  8'h73;        memory[41114] <=  8'h64;        memory[41115] <=  8'h66;        memory[41116] <=  8'h6b;        memory[41117] <=  8'h64;        memory[41118] <=  8'h6e;        memory[41119] <=  8'h6d;        memory[41120] <=  8'h64;        memory[41121] <=  8'h73;        memory[41122] <=  8'h63;        memory[41123] <=  8'h6b;        memory[41124] <=  8'h78;        memory[41125] <=  8'h6c;        memory[41126] <=  8'h6f;        memory[41127] <=  8'h66;        memory[41128] <=  8'h6a;        memory[41129] <=  8'h69;        memory[41130] <=  8'h61;        memory[41131] <=  8'h62;        memory[41132] <=  8'h6e;        memory[41133] <=  8'h20;        memory[41134] <=  8'h78;        memory[41135] <=  8'h6b;        memory[41136] <=  8'h6d;        memory[41137] <=  8'h20;        memory[41138] <=  8'h6f;        memory[41139] <=  8'h63;        memory[41140] <=  8'h76;        memory[41141] <=  8'h73;        memory[41142] <=  8'h64;        memory[41143] <=  8'h69;        memory[41144] <=  8'h66;        memory[41145] <=  8'h68;        memory[41146] <=  8'h65;        memory[41147] <=  8'h71;        memory[41148] <=  8'h6a;        memory[41149] <=  8'h77;        memory[41150] <=  8'h62;        memory[41151] <=  8'h65;        memory[41152] <=  8'h6e;        memory[41153] <=  8'h20;        memory[41154] <=  8'h6d;        memory[41155] <=  8'h64;        memory[41156] <=  8'h73;        memory[41157] <=  8'h6c;        memory[41158] <=  8'h76;        memory[41159] <=  8'h6b;        memory[41160] <=  8'h63;        memory[41161] <=  8'h78;        memory[41162] <=  8'h20;        memory[41163] <=  8'h6f;        memory[41164] <=  8'h78;        memory[41165] <=  8'h69;        memory[41166] <=  8'h63;        memory[41167] <=  8'h6a;        memory[41168] <=  8'h76;        memory[41169] <=  8'h64;        memory[41170] <=  8'h66;        memory[41171] <=  8'h65;        memory[41172] <=  8'h71;        memory[41173] <=  8'h6e;        memory[41174] <=  8'h20;        memory[41175] <=  8'h64;        memory[41176] <=  8'h6d;        memory[41177] <=  8'h73;        memory[41178] <=  8'h6c;        memory[41179] <=  8'h63;        memory[41180] <=  8'h78;        memory[41181] <=  8'h6b;        memory[41182] <=  8'h20;        memory[41183] <=  8'h6f;        memory[41184] <=  8'h78;        memory[41185] <=  8'h63;        memory[41186] <=  8'h76;        memory[41187] <=  8'h6a;        memory[41188] <=  8'h64;        memory[41189] <=  8'h62;        memory[41190] <=  8'h71;        memory[41191] <=  8'h77;        memory[41192] <=  8'h65;        memory[41193] <=  8'h6e;        memory[41194] <=  8'h6d;        memory[41195] <=  8'h64;        memory[41196] <=  8'h6c;        memory[41197] <=  8'h73;        memory[41198] <=  8'h2c;        memory[41199] <=  8'h76;        memory[41200] <=  8'h63;        memory[41201] <=  8'h78;        memory[41202] <=  8'h20;        memory[41203] <=  8'h63;        memory[41204] <=  8'h6f;        memory[41205] <=  8'h69;        memory[41206] <=  8'h76;        memory[41207] <=  8'h68;        memory[41208] <=  8'h73;        memory[41209] <=  8'h64;        memory[41210] <=  8'h62;        memory[41211] <=  8'h71;        memory[41212] <=  8'h77;        memory[41213] <=  8'h65;        memory[41214] <=  8'h6e;        memory[41215] <=  8'h64;        memory[41216] <=  8'h6b;        memory[41217] <=  8'h73;        memory[41218] <=  8'h76;        memory[41219] <=  8'h6f;        memory[41220] <=  8'h63;        memory[41221] <=  8'h20;        memory[41222] <=  8'h76;        memory[41223] <=  8'h69;        memory[41224] <=  8'h75;        memory[41225] <=  8'h69;        memory[41226] <=  8'h68;        memory[41227] <=  8'h63;        memory[41228] <=  8'h78;        memory[41229] <=  8'h69;        memory[41230] <=  8'h6f;        memory[41231] <=  8'h76;        memory[41232] <=  8'h73;        memory[41233] <=  8'h64;        memory[41234] <=  8'h61;        memory[41235] <=  8'h64;        memory[41236] <=  8'h6e;        memory[41237] <=  8'h77;        memory[41238] <=  8'h71;        memory[41239] <=  8'h6b;        memory[41240] <=  8'h6c;        memory[41241] <=  8'h73;        memory[41242] <=  8'h76;        memory[41243] <=  8'h6e;        memory[41244] <=  8'h62;        memory[41245] <=  8'h20;        memory[41246] <=  8'h64;        memory[41247] <=  8'h66;        memory[41248] <=  8'h6a;        memory[41249] <=  8'h6b;        memory[41250] <=  8'h71;        memory[41251] <=  8'h64;        memory[41252] <=  8'h77;        memory[41253] <=  8'h65;        memory[41254] <=  8'h6e;        memory[41255] <=  8'h62;        memory[41256] <=  8'h20;        memory[41257] <=  8'h64;        memory[41258] <=  8'h73;        memory[41259] <=  8'h76;        memory[41260] <=  8'h68;        memory[41261] <=  8'h64;        memory[41262] <=  8'h61;        memory[41263] <=  8'h71;        memory[41264] <=  8'h77;        memory[41265] <=  8'h6a;        memory[41266] <=  8'h65;        memory[41267] <=  8'h6e;        memory[41268] <=  8'h64;        memory[41269] <=  8'h20;        memory[41270] <=  8'h61;        memory[41271] <=  8'h63;        memory[41272] <=  8'h62;        memory[41273] <=  8'h68;        memory[41274] <=  8'h64;        memory[41275] <=  8'h61;        memory[41276] <=  8'h77;        memory[41277] <=  8'h71;        memory[41278] <=  8'h6e;        memory[41279] <=  8'h20;        memory[41280] <=  8'h62;        memory[41281] <=  8'h73;        memory[41282] <=  8'h76;        memory[41283] <=  8'h61;        memory[41284] <=  8'h67;        memory[41285] <=  8'h76;        memory[41286] <=  8'h68;        memory[41287] <=  8'h67;        memory[41288] <=  8'h61;        memory[41289] <=  8'h73;        memory[41290] <=  8'h6a;        memory[41291] <=  8'h6b;        memory[41292] <=  8'h63;        memory[41293] <=  8'h78;        memory[41294] <=  8'h76;        memory[41295] <=  8'h6e;        memory[41296] <=  8'h73;        memory[41297] <=  8'h64;        memory[41298] <=  8'h20;        memory[41299] <=  8'h66;        memory[41300] <=  8'h62;        memory[41301] <=  8'h64;        memory[41302] <=  8'h61;        memory[41303] <=  8'h73;        memory[41304] <=  8'h76;        memory[41305] <=  8'h67;        memory[41306] <=  8'h63;        memory[41307] <=  8'h79;        memory[41308] <=  8'h7a;        memory[41309] <=  8'h78;        memory[41310] <=  8'h79;        memory[41311] <=  8'h75;        memory[41312] <=  8'h20;        memory[41313] <=  8'h69;        memory[41314] <=  8'h6a;        memory[41315] <=  8'h64;        memory[41316] <=  8'h66;        memory[41317] <=  8'h6b;        memory[41318] <=  8'h61;        memory[41319] <=  8'h64;        memory[41320] <=  8'h63;        memory[41321] <=  8'h78;        memory[41322] <=  8'h68;        memory[41323] <=  8'h20;        memory[41324] <=  8'h67;        memory[41325] <=  8'h61;        memory[41326] <=  8'h68;        memory[41327] <=  8'h75;        memory[41328] <=  8'h64;        memory[41329] <=  8'h73;        memory[41330] <=  8'h69;        memory[41331] <=  8'h6a;        memory[41332] <=  8'h61;        memory[41333] <=  8'h6b;        memory[41334] <=  8'h63;        memory[41335] <=  8'h62;        memory[41336] <=  8'h61;        memory[41337] <=  8'h72;        memory[41338] <=  8'h73;        memory[41339] <=  8'h68;        memory[41340] <=  8'h64;        memory[41341] <=  8'h66;        memory[41342] <=  8'h67;        memory[41343] <=  8'h73;        memory[41344] <=  8'h68;        memory[41345] <=  8'h64;        memory[41346] <=  8'h66;        memory[41347] <=  8'h68;        memory[41348] <=  8'h64;        memory[41349] <=  8'h6a;        memory[41350] <=  8'h68;        memory[41351] <=  8'h62;        memory[41352] <=  8'h67;        memory[41353] <=  8'h63;        memory[41354] <=  8'h61;        memory[41355] <=  8'h66;        memory[41356] <=  8'h73;        memory[41357] <=  8'h79;        memory[41358] <=  8'h67;        memory[41359] <=  8'h6b;        memory[41360] <=  8'h75;        memory[41361] <=  8'h64;        memory[41362] <=  8'h68;        memory[41363] <=  8'h62;        memory[41364] <=  8'h77;        memory[41365] <=  8'h76;        memory[41366] <=  8'h67;        memory[41367] <=  8'h61;        memory[41368] <=  8'h66;        memory[41369] <=  8'h64;        memory[41370] <=  8'h74;        memory[41371] <=  8'h75;        memory[41372] <=  8'h66;        memory[41373] <=  8'h79;        memory[41374] <=  8'h67;        memory[41375] <=  8'h69;        memory[41376] <=  8'h75;        memory[41377] <=  8'h68;        memory[41378] <=  8'h6c;        memory[41379] <=  8'h6a;        memory[41380] <=  8'h62;        memory[41381] <=  8'h6b;        memory[41382] <=  8'h68;        memory[41383] <=  8'h76;        memory[41384] <=  8'h67;        memory[41385] <=  8'h63;        memory[41386] <=  8'h66;        memory[41387] <=  8'h78;        memory[41388] <=  8'h64;        memory[41389] <=  8'h74;        memory[41390] <=  8'h75;        memory[41391] <=  8'h79;        memory[41392] <=  8'h69;        memory[41393] <=  8'h75;        memory[41394] <=  8'h68;        memory[41395] <=  8'h6c;        memory[41396] <=  8'h6a;        memory[41397] <=  8'h6b;        memory[41398] <=  8'h67;        memory[41399] <=  8'h6a;        memory[41400] <=  8'h63;        memory[41401] <=  8'h66;        memory[41402] <=  8'h68;        memory[41403] <=  8'h64;        memory[41404] <=  8'h67;        memory[41405] <=  8'h72;        memory[41406] <=  8'h79;        memory[41407] <=  8'h74;        memory[41408] <=  8'h66;        memory[41409] <=  8'h75;        memory[41410] <=  8'h79;        memory[41411] <=  8'h69;        memory[41412] <=  8'h68;        memory[41413] <=  8'h6c;        memory[41414] <=  8'h62;        memory[41415] <=  8'h6d;        memory[41416] <=  8'h76;        memory[41417] <=  8'h6e;        memory[41418] <=  8'h63;        memory[41419] <=  8'h66;        memory[41420] <=  8'h68;        memory[41421] <=  8'h64;        memory[41422] <=  8'h74;        memory[41423] <=  8'h75;        memory[41424] <=  8'h67;        memory[41425] <=  8'h79;        memory[41426] <=  8'h69;        memory[41427] <=  8'h68;        memory[41428] <=  8'h75;        memory[41429] <=  8'h6a;        memory[41430] <=  8'h6c;        memory[41431] <=  8'h62;        memory[41432] <=  8'h6d;        memory[41433] <=  8'h76;        memory[41434] <=  8'h6e;        memory[41435] <=  8'h63;        memory[41436] <=  8'h66;        memory[41437] <=  8'h68;        memory[41438] <=  8'h67;        memory[41439] <=  8'h79;        memory[41440] <=  8'h68;        memory[41441] <=  8'h75;        memory[41442] <=  8'h6a;        memory[41443] <=  8'h6e;        memory[41444] <=  8'h2c;        memory[41445] <=  8'h62;        memory[41446] <=  8'h6e;        memory[41447] <=  8'h6d;        memory[41448] <=  8'h76;        memory[41449] <=  8'h6e;        memory[41450] <=  8'h63;        memory[41451] <=  8'h66;        memory[41452] <=  8'h68;        memory[41453] <=  8'h74;        memory[41454] <=  8'h79;        memory[41455] <=  8'h69;        memory[41456] <=  8'h75;        memory[41457] <=  8'h6c;        memory[41458] <=  8'h6a;        memory[41459] <=  8'h62;        memory[41460] <=  8'h6d;        memory[41461] <=  8'h76;        memory[41462] <=  8'h6e;        memory[41463] <=  8'h63;        memory[41464] <=  8'h66;        memory[41465] <=  8'h74;        memory[41466] <=  8'h75;        memory[41467] <=  8'h79;        memory[41468] <=  8'h69;        memory[41469] <=  8'h68;        memory[41470] <=  8'h6b;        memory[41471] <=  8'h62;        memory[41472] <=  8'h76;        memory[41473] <=  8'h63;        memory[41474] <=  8'h66;        memory[41475] <=  8'h67;        memory[41476] <=  8'h74;        memory[41477] <=  8'h75;        memory[41478] <=  8'h79;        memory[41479] <=  8'h69;        memory[41480] <=  8'h75;        memory[41481] <=  8'h68;        memory[41482] <=  8'h6a;        memory[41483] <=  8'h6b;        memory[41484] <=  8'h62;        memory[41485] <=  8'h76;        memory[41486] <=  8'h63;        memory[41487] <=  8'h66;        memory[41488] <=  8'h74;        memory[41489] <=  8'h75;        memory[41490] <=  8'h79;        memory[41491] <=  8'h69;        memory[41492] <=  8'h75;        memory[41493] <=  8'h6a;        memory[41494] <=  8'h6b;        memory[41495] <=  8'h6e;        memory[41496] <=  8'h62;        memory[41497] <=  8'h76;        memory[41498] <=  8'h67;        memory[41499] <=  8'h66;        memory[41500] <=  8'h74;        memory[41501] <=  8'h79;        memory[41502] <=  8'h75;        memory[41503] <=  8'h75;        memory[41504] <=  8'h69;        memory[41505] <=  8'h6a;        memory[41506] <=  8'h6b;        memory[41507] <=  8'h68;        memory[41508] <=  8'h62;        memory[41509] <=  8'h6a;        memory[41510] <=  8'h67;        memory[41511] <=  8'h68;        memory[41512] <=  8'h66;        memory[41513] <=  8'h79;        memory[41514] <=  8'h74;        memory[41515] <=  8'h79;        memory[41516] <=  8'h69;        memory[41517] <=  8'h75;        memory[41518] <=  8'h64;        memory[41519] <=  8'h6a;        memory[41520] <=  8'h6b;        memory[41521] <=  8'h68;        memory[41522] <=  8'h63;        memory[41523] <=  8'h7a;        memory[41524] <=  8'h67;        memory[41525] <=  8'h68;        memory[41526] <=  8'h74;        memory[41527] <=  8'h75;        memory[41528] <=  8'h79;        memory[41529] <=  8'h69;        memory[41530] <=  8'h61;        memory[41531] <=  8'h73;        memory[41532] <=  8'h75;        memory[41533] <=  8'h6a;        memory[41534] <=  8'h6b;        memory[41535] <=  8'h62;        memory[41536] <=  8'h6e;        memory[41537] <=  8'h61;        memory[41538] <=  8'h76;        memory[41539] <=  8'h63;        memory[41540] <=  8'h66;        memory[41541] <=  8'h68;        memory[41542] <=  8'h75;        memory[41543] <=  8'h61;        memory[41544] <=  8'h73;        memory[41545] <=  8'h79;        memory[41546] <=  8'h64;        memory[41547] <=  8'h75;        memory[41548] <=  8'h69;        memory[41549] <=  8'h6a;        memory[41550] <=  8'h61;        memory[41551] <=  8'h6b;        memory[41552] <=  8'h62;        memory[41553] <=  8'h63;        memory[41554] <=  8'h78;        memory[41555] <=  8'h68;        memory[41556] <=  8'h67;        memory[41557] <=  8'h79;        memory[41558] <=  8'h75;        memory[41559] <=  8'h7a;        memory[41560] <=  8'h63;        memory[41561] <=  8'h61;        memory[41562] <=  8'h73;        memory[41563] <=  8'h69;        memory[41564] <=  8'h75;        memory[41565] <=  8'h6f;        memory[41566] <=  8'h69;        memory[41567] <=  8'h6a;        memory[41568] <=  8'h61;        memory[41569] <=  8'h6c;        memory[41570] <=  8'h63;        memory[41571] <=  8'h78;        memory[41572] <=  8'h62;        memory[41573] <=  8'h63;        memory[41574] <=  8'h20;        memory[41575] <=  8'h6e;        memory[41576] <=  8'h76;        memory[41577] <=  8'h63;        memory[41578] <=  8'h61;        memory[41579] <=  8'h64;        memory[41580] <=  8'h73;        memory[41581] <=  8'h67;        memory[41582] <=  8'h79;        memory[41583] <=  8'h68;        memory[41584] <=  8'h75;        memory[41585] <=  8'h61;        memory[41586] <=  8'h6a;        memory[41587] <=  8'h6b;        memory[41588] <=  8'h78;        memory[41589] <=  8'h62;        memory[41590] <=  8'h20;        memory[41591] <=  8'h6e;        memory[41592] <=  8'h76;        memory[41593] <=  8'h63;        memory[41594] <=  8'h61;        memory[41595] <=  8'h73;        memory[41596] <=  8'h67;        memory[41597] <=  8'h68;        memory[41598] <=  8'h75;        memory[41599] <=  8'h6a;        memory[41600] <=  8'h6c;        memory[41601] <=  8'h6b;        memory[41602] <=  8'h63;        memory[41603] <=  8'h78;        memory[41604] <=  8'h20;        memory[41605] <=  8'h6a;        memory[41606] <=  8'h6b;        memory[41607] <=  8'h68;        memory[41608] <=  8'h61;        memory[41609] <=  8'h73;        memory[41610] <=  8'h76;        memory[41611] <=  8'h64;        memory[41612] <=  8'h6e;        memory[41613] <=  8'h20;        memory[41614] <=  8'h62;        memory[41615] <=  8'h6e;        memory[41616] <=  8'h6d;        memory[41617] <=  8'h6b;        memory[41618] <=  8'h77;        memory[41619] <=  8'h64;        memory[41620] <=  8'h6f;        memory[41621] <=  8'h77;        memory[41622] <=  8'h69;        memory[41623] <=  8'h6f;        memory[41624] <=  8'h75;        memory[41625] <=  8'h69;        memory[41626] <=  8'h68;        memory[41627] <=  8'h62;        memory[41628] <=  8'h6e;        memory[41629] <=  8'h6b;        memory[41630] <=  8'h77;        memory[41631] <=  8'h69;        memory[41632] <=  8'h6f;        memory[41633] <=  8'h75;        memory[41634] <=  8'h71;        memory[41635] <=  8'h69;        memory[41636] <=  8'h79;        memory[41637] <=  8'h67;        memory[41638] <=  8'h6a;        memory[41639] <=  8'h64;        memory[41640] <=  8'h61;        memory[41641] <=  8'h76;        memory[41642] <=  8'h62;        memory[41643] <=  8'h6e;        memory[41644] <=  8'h6b;        memory[41645] <=  8'h6f;        memory[41646] <=  8'h70;        memory[41647] <=  8'h64;        memory[41648] <=  8'h76;        memory[41649] <=  8'h69;        memory[41650] <=  8'h6f;        memory[41651] <=  8'h75;        memory[41652] <=  8'h69;        memory[41653] <=  8'h48;        memory[41654] <=  8'h42;        memory[41655] <=  8'h6b;        memory[41656] <=  8'h64;        memory[41657] <=  8'h6e;        memory[41658] <=  8'h6c;        memory[41659] <=  8'h71;        memory[41660] <=  8'h6b;        memory[41661] <=  8'h6d;        memory[41662] <=  8'h6a;        memory[41663] <=  8'h70;        memory[41664] <=  8'h69;        memory[41665] <=  8'h6f;        memory[41666] <=  8'h68;        memory[41667] <=  8'h65;        memory[41668] <=  8'h66;        memory[41669] <=  8'h75;        memory[41670] <=  8'h67;        memory[41671] <=  8'h69;        memory[41672] <=  8'h73;        memory[41673] <=  8'h61;        memory[41674] <=  8'h62;        memory[41675] <=  8'h64;        memory[41676] <=  8'h6b;        memory[41677] <=  8'h6a;        memory[41678] <=  8'h6b;        memory[41679] <=  8'h6c;        memory[41680] <=  8'h6a;        memory[41681] <=  8'h69;        memory[41682] <=  8'h73;        memory[41683] <=  8'h6f;        memory[41684] <=  8'h71;        memory[41685] <=  8'h68;        memory[41686] <=  8'h77;        memory[41687] <=  8'h67;        memory[41688] <=  8'h69;        memory[41689] <=  8'h79;        memory[41690] <=  8'h6a;        memory[41691] <=  8'h64;        memory[41692] <=  8'h76;        memory[41693] <=  8'h62;        memory[41694] <=  8'h6e;        memory[41695] <=  8'h61;        memory[41696] <=  8'h73;        memory[41697] <=  8'h66;        memory[41698] <=  8'h6c;        memory[41699] <=  8'h6b;        memory[41700] <=  8'h64;        memory[41701] <=  8'h6a;        memory[41702] <=  8'h68;        memory[41703] <=  8'h63;        memory[41704] <=  8'h67;        memory[41705] <=  8'h6a;        memory[41706] <=  8'h76;        memory[41707] <=  8'h73;        memory[41708] <=  8'h64;        memory[41709] <=  8'h62;        memory[41710] <=  8'h62;        memory[41711] <=  8'h61;        memory[41712] <=  8'h72;        memory[41713] <=  8'h62;        memory[41714] <=  8'h62;        memory[41715] <=  8'h73;        memory[41716] <=  8'h62;        memory[41717] <=  8'h67;        memory[41718] <=  8'h73;        memory[41719] <=  8'h66;        memory[41720] <=  8'h67;        memory[41721] <=  8'h61;        memory[41722] <=  8'h68;        memory[41723] <=  8'h66;        memory[41724] <=  8'h73;        memory[41725] <=  8'h68;        memory[41726] <=  8'h61;        memory[41727] <=  8'h66;        memory[41728] <=  8'h73;        memory[41729] <=  8'h66;        memory[41730] <=  8'h68;        memory[41731] <=  8'h61;        memory[41732] <=  8'h69;        memory[41733] <=  8'h64;        memory[41734] <=  8'h75;        memory[41735] <=  8'h67;        memory[41736] <=  8'h64;        memory[41737] <=  8'h77;        memory[41738] <=  8'h62;        memory[41739] <=  8'h61;        memory[41740] <=  8'h62;        memory[41741] <=  8'h72;        memory[41742] <=  8'h62;        memory[41743] <=  8'h61;        memory[41744] <=  8'h62;        memory[41745] <=  8'h62;        memory[41746] <=  8'h74;        memory[41747] <=  8'h62;        memory[41748] <=  8'h62;        memory[41749] <=  8'h62;        memory[41750] <=  8'h62;        memory[41751] <=  8'h62;        memory[41752] <=  8'h62;        memory[41753] <=  8'h62;        memory[41754] <=  8'h62;        memory[41755] <=  8'h61;        memory[41756] <=  8'h62;        memory[41757] <=  8'h62;        memory[41758] <=  8'h72;        memory[41759] <=  8'h74;        memory[41760] <=  8'h62;        memory[41761] <=  8'h62;        memory[41762] <=  8'h61;        memory[41763] <=  8'h62;        memory[41764] <=  8'h72;        memory[41765] <=  8'h62;        memory[41766] <=  8'h74;        memory[41767] <=  8'h62;        memory[41768] <=  8'h62;        memory[41769] <=  8'h62;        memory[41770] <=  8'h63;        memory[41771] <=  8'h61;        memory[41772] <=  8'h72;        memory[41773] <=  8'h74;        memory[41774] <=  8'h73;        memory[41775] <=  8'h62;        memory[41776] <=  8'h61;        memory[41777] <=  8'h72;        memory[41778] <=  8'h74;        memory[41779] <=  8'h74;        memory[41780] <=  8'h62;        memory[41781] <=  8'h61;        memory[41782] <=  8'h72;        memory[41783] <=  8'h74;        memory[41784] <=  8'h78;        memory[41785] <=  8'h61;        memory[41786] <=  8'h74;        memory[41787] <=  8'h6b;        memory[41788] <=  8'h73;        memory[41789] <=  8'h68;        memory[41790] <=  8'h63;        memory[41791] <=  8'h66;        memory[41792] <=  8'h69;        memory[41793] <=  8'h77;        memory[41794] <=  8'h68;        memory[41795] <=  8'h61;        memory[41796] <=  8'h74;        memory[41797] <=  8'h61;        memory[41798] <=  8'h6e;        memory[41799] <=  8'h61;        memory[41800] <=  8'h62;        memory[41801] <=  8'h61;        memory[41802] <=  8'h63;        memory[41803] <=  8'h61;        memory[41804] <=  8'h74;        memory[41805] <=  8'h61;        memory[41806] <=  8'h62;        memory[41807] <=  8'h61;        memory[41808] <=  8'h72;        memory[41809] <=  8'h63;        memory[41810] <=  8'h61;        memory[41811] <=  8'h68;        memory[41812] <=  8'h64;        memory[41813] <=  8'h75;        memory[41814] <=  8'h63;        memory[41815] <=  8'h74;        memory[41816] <=  8'h61;        memory[41817] <=  8'h64;        memory[41818] <=  8'h61;        memory[41819] <=  8'h61;        memory[41820] <=  8'h63;        memory[41821] <=  8'h61;        memory[41822] <=  8'h72;        memory[41823] <=  8'h63;        memory[41824] <=  8'h74;        memory[41825] <=  8'h72;        memory[41826] <=  8'h63;        memory[41827] <=  8'h61;        memory[41828] <=  8'h74;        memory[41829] <=  8'h72;        memory[41830] <=  8'h63;        memory[41831] <=  8'h61;        memory[41832] <=  8'h74;        memory[41833] <=  8'h63;        memory[41834] <=  8'h62;        memory[41835] <=  8'h61;        memory[41836] <=  8'h74;        memory[41837] <=  8'h62;        memory[41838] <=  8'h72;        memory[41839] <=  8'h63;        memory[41840] <=  8'h61;        memory[41841] <=  8'h74;        memory[41842] <=  8'h72;        memory[41843] <=  8'h6e;        memory[41844] <=  8'h62;        memory[41845] <=  8'h61;        memory[41846] <=  8'h63;        memory[41847] <=  8'h61;        memory[41848] <=  8'h74;        memory[41849] <=  8'h79;        memory[41850] <=  8'h73;        memory[41851] <=  8'h6e;        memory[41852] <=  8'h63;        memory[41853] <=  8'h74;        memory[41854] <=  8'h61;        memory[41855] <=  8'h6e;        memory[41856] <=  8'h62;        memory[41857] <=  8'h61;        memory[41858] <=  8'h63;        memory[41859] <=  8'h72;        memory[41860] <=  8'h6e;        memory[41861] <=  8'h74;        memory[41862] <=  8'h61;        memory[41863] <=  8'h62;        memory[41864] <=  8'h74;        memory[41865] <=  8'h6e;        memory[41866] <=  8'h61;        memory[41867] <=  8'h72;        memory[41868] <=  8'h62;        memory[41869] <=  8'h78;        memory[41870] <=  8'h74;        memory[41871] <=  8'h61;        memory[41872] <=  8'h72;        memory[41873] <=  8'h62;        memory[41874] <=  8'h61;        memory[41875] <=  8'h72;        memory[41876] <=  8'h74;        memory[41877] <=  8'h74;        memory[41878] <=  8'h62;        memory[41879] <=  8'h61;        memory[41880] <=  8'h72;        memory[41881] <=  8'h74;        memory[41882] <=  8'h78;        memory[41883] <=  8'h61;        memory[41884] <=  8'h74;        memory[41885] <=  8'h6b;        memory[41886] <=  8'h73;        memory[41887] <=  8'h68;        memory[41888] <=  8'h63;        memory[41889] <=  8'h66;        memory[41890] <=  8'h69;        memory[41891] <=  8'h77;        memory[41892] <=  8'h68;        memory[41893] <=  8'h61;        memory[41894] <=  8'h74;        memory[41895] <=  8'h61;        memory[41896] <=  8'h6e;        memory[41897] <=  8'h61;        memory[41898] <=  8'h62;        memory[41899] <=  8'h61;        memory[41900] <=  8'h63;        memory[41901] <=  8'h61;        memory[41902] <=  8'h74;        memory[41903] <=  8'h61;        memory[41904] <=  8'h62;        memory[41905] <=  8'h61;        memory[41906] <=  8'h72;        memory[41907] <=  8'h63;        memory[41908] <=  8'h61;        memory[41909] <=  8'h68;        memory[41910] <=  8'h64;        memory[41911] <=  8'h75;        memory[41912] <=  8'h63;        memory[41913] <=  8'h74;        memory[41914] <=  8'h61;        memory[41915] <=  8'h64;        memory[41916] <=  8'h61;        memory[41917] <=  8'h61;        memory[41918] <=  8'h63;        memory[41919] <=  8'h61;        memory[41920] <=  8'h72;        memory[41921] <=  8'h63;        memory[41922] <=  8'h74;        memory[41923] <=  8'h72;        memory[41924] <=  8'h63;        memory[41925] <=  8'h61;        memory[41926] <=  8'h74;        memory[41927] <=  8'h72;        memory[41928] <=  8'h63;        memory[41929] <=  8'h61;        memory[41930] <=  8'h74;        memory[41931] <=  8'h63;        memory[41932] <=  8'h62;        memory[41933] <=  8'h61;        memory[41934] <=  8'h74;        memory[41935] <=  8'h62;        memory[41936] <=  8'h72;        memory[41937] <=  8'h63;        memory[41938] <=  8'h61;        memory[41939] <=  8'h74;        memory[41940] <=  8'h72;        memory[41941] <=  8'h6e;        memory[41942] <=  8'h62;        memory[41943] <=  8'h61;        memory[41944] <=  8'h63;        memory[41945] <=  8'h61;        memory[41946] <=  8'h74;        memory[41947] <=  8'h79;        memory[41948] <=  8'h73;        memory[41949] <=  8'h6e;        memory[41950] <=  8'h63;        memory[41951] <=  8'h74;        memory[41952] <=  8'h61;        memory[41953] <=  8'h6e;        memory[41954] <=  8'h62;        memory[41955] <=  8'h61;        memory[41956] <=  8'h63;        memory[41957] <=  8'h72;        memory[41958] <=  8'h6e;        memory[41959] <=  8'h74;        memory[41960] <=  8'h61;        memory[41961] <=  8'h62;        memory[41962] <=  8'h74;        memory[41963] <=  8'h6e;        memory[41964] <=  8'h61;        memory[41965] <=  8'h72;        memory[41966] <=  8'h62;        memory[41967] <=  8'h78;        memory[41968] <=  8'h74;        memory[41969] <=  8'h61;        memory[41970] <=  8'h72;        memory[41971] <=  8'h62;        memory[41972] <=  8'h61;        memory[41973] <=  8'h72;        memory[41974] <=  8'h74;        memory[41975] <=  8'h74;        memory[41976] <=  8'h62;        memory[41977] <=  8'h61;        memory[41978] <=  8'h72;        memory[41979] <=  8'h74;        memory[41980] <=  8'h78;        memory[41981] <=  8'h61;        memory[41982] <=  8'h74;        memory[41983] <=  8'h6b;        memory[41984] <=  8'h73;        memory[41985] <=  8'h68;        memory[41986] <=  8'h63;        memory[41987] <=  8'h66;        memory[41988] <=  8'h69;        memory[41989] <=  8'h77;        memory[41990] <=  8'h68;        memory[41991] <=  8'h61;        memory[41992] <=  8'h74;        memory[41993] <=  8'h61;        memory[41994] <=  8'h6e;        memory[41995] <=  8'h61;        memory[41996] <=  8'h62;        memory[41997] <=  8'h61;        memory[41998] <=  8'h63;        memory[41999] <=  8'h61;        memory[42000] <=  8'h74;        memory[42001] <=  8'h61;        memory[42002] <=  8'h62;        memory[42003] <=  8'h61;        memory[42004] <=  8'h72;        memory[42005] <=  8'h63;        memory[42006] <=  8'h61;        memory[42007] <=  8'h68;        memory[42008] <=  8'h64;        memory[42009] <=  8'h75;        memory[42010] <=  8'h63;        memory[42011] <=  8'h74;        memory[42012] <=  8'h61;        memory[42013] <=  8'h64;        memory[42014] <=  8'h61;        memory[42015] <=  8'h61;        memory[42016] <=  8'h63;        memory[42017] <=  8'h61;        memory[42018] <=  8'h72;        memory[42019] <=  8'h63;        memory[42020] <=  8'h74;        memory[42021] <=  8'h72;        memory[42022] <=  8'h63;        memory[42023] <=  8'h61;        memory[42024] <=  8'h74;        memory[42025] <=  8'h72;        memory[42026] <=  8'h63;        memory[42027] <=  8'h61;        memory[42028] <=  8'h74;        memory[42029] <=  8'h63;        memory[42030] <=  8'h62;        memory[42031] <=  8'h61;        memory[42032] <=  8'h74;        memory[42033] <=  8'h62;        memory[42034] <=  8'h72;        memory[42035] <=  8'h63;        memory[42036] <=  8'h61;        memory[42037] <=  8'h74;        memory[42038] <=  8'h72;        memory[42039] <=  8'h6e;        memory[42040] <=  8'h62;        memory[42041] <=  8'h61;        memory[42042] <=  8'h63;        memory[42043] <=  8'h61;        memory[42044] <=  8'h74;        memory[42045] <=  8'h79;        memory[42046] <=  8'h73;        memory[42047] <=  8'h6e;        memory[42048] <=  8'h63;        memory[42049] <=  8'h74;        memory[42050] <=  8'h61;        memory[42051] <=  8'h6e;        memory[42052] <=  8'h62;        memory[42053] <=  8'h61;        memory[42054] <=  8'h63;        memory[42055] <=  8'h72;        memory[42056] <=  8'h6e;        memory[42057] <=  8'h74;        memory[42058] <=  8'h61;        memory[42059] <=  8'h62;        memory[42060] <=  8'h74;        memory[42061] <=  8'h6e;        memory[42062] <=  8'h61;        memory[42063] <=  8'h72;        memory[42064] <=  8'h62;        memory[42065] <=  8'h78;        memory[42066] <=  8'h74;        memory[42067] <=  8'h61;        memory[42068] <=  8'h72;        memory[42069] <=  8'h5d;        memory[42070] <=  8'h5d;        memory[42071] <=  8'h65;        memory[42072] <=  8'h66;        memory[42073] <=  8'h77;        memory[42074] <=  8'h65;        memory[42075] <=  8'h5d;        memory[42076] <=  8'h65;        memory[42077] <=  8'h67;        memory[42078] <=  8'h73;        memory[42079] <=  8'h67;        memory[42080] <=  8'h66;        memory[42081] <=  8'h62;        memory[42082] <=  8'h61;        memory[42083] <=  8'h72;        memory[42084] <=  8'h74;        memory[42085] <=  8'h74;        memory[42086] <=  8'h62;        memory[42087] <=  8'h61;        memory[42088] <=  8'h72;        memory[42089] <=  8'h74;        memory[42090] <=  8'h78;        memory[42091] <=  8'h61;        memory[42092] <=  8'h74;        memory[42093] <=  8'h6b;        memory[42094] <=  8'h73;        memory[42095] <=  8'h68;        memory[42096] <=  8'h63;        memory[42097] <=  8'h66;        memory[42098] <=  8'h69;        memory[42099] <=  8'h77;        memory[42100] <=  8'h68;        memory[42101] <=  8'h61;        memory[42102] <=  8'h74;        memory[42103] <=  8'h61;        memory[42104] <=  8'h6e;        memory[42105] <=  8'h61;        memory[42106] <=  8'h62;        memory[42107] <=  8'h61;        memory[42108] <=  8'h63;        memory[42109] <=  8'h61;        memory[42110] <=  8'h74;        memory[42111] <=  8'h61;        memory[42112] <=  8'h62;        memory[42113] <=  8'h61;        memory[42114] <=  8'h72;        memory[42115] <=  8'h63;        memory[42116] <=  8'h61;        memory[42117] <=  8'h68;        memory[42118] <=  8'h64;        memory[42119] <=  8'h75;        memory[42120] <=  8'h63;        memory[42121] <=  8'h74;        memory[42122] <=  8'h61;        memory[42123] <=  8'h64;        memory[42124] <=  8'h61;        memory[42125] <=  8'h61;        memory[42126] <=  8'h63;        memory[42127] <=  8'h61;        memory[42128] <=  8'h72;        memory[42129] <=  8'h63;        memory[42130] <=  8'h74;        memory[42131] <=  8'h72;        memory[42132] <=  8'h63;        memory[42133] <=  8'h61;        memory[42134] <=  8'h74;        memory[42135] <=  8'h72;        memory[42136] <=  8'h63;        memory[42137] <=  8'h61;        memory[42138] <=  8'h74;        memory[42139] <=  8'h63;        memory[42140] <=  8'h62;        memory[42141] <=  8'h61;        memory[42142] <=  8'h74;        memory[42143] <=  8'h62;        memory[42144] <=  8'h72;        memory[42145] <=  8'h63;        memory[42146] <=  8'h61;        memory[42147] <=  8'h74;        memory[42148] <=  8'h72;        memory[42149] <=  8'h6e;        memory[42150] <=  8'h62;        memory[42151] <=  8'h61;        memory[42152] <=  8'h63;        memory[42153] <=  8'h61;        memory[42154] <=  8'h74;        memory[42155] <=  8'h79;        memory[42156] <=  8'h73;        memory[42157] <=  8'h6e;        memory[42158] <=  8'h63;        memory[42159] <=  8'h74;        memory[42160] <=  8'h61;        memory[42161] <=  8'h6e;        memory[42162] <=  8'h62;        memory[42163] <=  8'h61;        memory[42164] <=  8'h63;        memory[42165] <=  8'h72;        memory[42166] <=  8'h6e;        memory[42167] <=  8'h74;        memory[42168] <=  8'h61;        memory[42169] <=  8'h62;        memory[42170] <=  8'h74;        memory[42171] <=  8'h6e;        memory[42172] <=  8'h61;        memory[42173] <=  8'h72;        memory[42174] <=  8'h62;        memory[42175] <=  8'h78;        memory[42176] <=  8'h74;        memory[42177] <=  8'h61;        memory[42178] <=  8'h72;        memory[42179] <=  8'h62;        memory[42180] <=  8'h61;        memory[42181] <=  8'h72;        memory[42182] <=  8'h74;        memory[42183] <=  8'h74;        memory[42184] <=  8'h62;        memory[42185] <=  8'h61;        memory[42186] <=  8'h72;        memory[42187] <=  8'h74;        memory[42188] <=  8'h78;        memory[42189] <=  8'h61;        memory[42190] <=  8'h74;        memory[42191] <=  8'h6b;        memory[42192] <=  8'h73;        memory[42193] <=  8'h68;        memory[42194] <=  8'h63;        memory[42195] <=  8'h66;        memory[42196] <=  8'h69;        memory[42197] <=  8'h77;        memory[42198] <=  8'h68;        memory[42199] <=  8'h61;        memory[42200] <=  8'h74;        memory[42201] <=  8'h61;        memory[42202] <=  8'h6e;        memory[42203] <=  8'h61;        memory[42204] <=  8'h62;        memory[42205] <=  8'h61;        memory[42206] <=  8'h63;        memory[42207] <=  8'h61;        memory[42208] <=  8'h74;        memory[42209] <=  8'h61;        memory[42210] <=  8'h62;        memory[42211] <=  8'h61;        memory[42212] <=  8'h72;        memory[42213] <=  8'h63;        memory[42214] <=  8'h61;        memory[42215] <=  8'h68;        memory[42216] <=  8'h64;        memory[42217] <=  8'h75;        memory[42218] <=  8'h63;        memory[42219] <=  8'h74;        memory[42220] <=  8'h61;        memory[42221] <=  8'h64;        memory[42222] <=  8'h61;        memory[42223] <=  8'h61;        memory[42224] <=  8'h63;        memory[42225] <=  8'h61;        memory[42226] <=  8'h72;        memory[42227] <=  8'h63;        memory[42228] <=  8'h74;        memory[42229] <=  8'h72;        memory[42230] <=  8'h63;        memory[42231] <=  8'h61;        memory[42232] <=  8'h74;        memory[42233] <=  8'h72;        memory[42234] <=  8'h63;        memory[42235] <=  8'h61;        memory[42236] <=  8'h74;        memory[42237] <=  8'h63;        memory[42238] <=  8'h62;        memory[42239] <=  8'h61;        memory[42240] <=  8'h74;        memory[42241] <=  8'h62;        memory[42242] <=  8'h72;        memory[42243] <=  8'h63;        memory[42244] <=  8'h61;        memory[42245] <=  8'h74;        memory[42246] <=  8'h72;        memory[42247] <=  8'h6e;        memory[42248] <=  8'h62;        memory[42249] <=  8'h61;        memory[42250] <=  8'h63;        memory[42251] <=  8'h61;        memory[42252] <=  8'h74;        memory[42253] <=  8'h79;        memory[42254] <=  8'h73;        memory[42255] <=  8'h6e;        memory[42256] <=  8'h63;        memory[42257] <=  8'h74;        memory[42258] <=  8'h61;        memory[42259] <=  8'h6e;        memory[42260] <=  8'h62;        memory[42261] <=  8'h61;        memory[42262] <=  8'h63;        memory[42263] <=  8'h72;        memory[42264] <=  8'h6e;        memory[42265] <=  8'h74;        memory[42266] <=  8'h61;        memory[42267] <=  8'h62;        memory[42268] <=  8'h74;        memory[42269] <=  8'h6e;        memory[42270] <=  8'h61;        memory[42271] <=  8'h72;        memory[42272] <=  8'h62;        memory[42273] <=  8'h78;        memory[42274] <=  8'h74;        memory[42275] <=  8'h61;        memory[42276] <=  8'h72;        memory[42277] <=  8'h64;        memory[42278] <=  8'h66;        memory[42279] <=  8'h73;        memory[42280] <=  8'h67;        memory[42281] <=  8'h76;        memory[42282] <=  8'h68;        memory[42283] <=  8'h62;        memory[42284] <=  8'h6b;        memory[42285] <=  8'h6a;        memory[42286] <=  8'h6e;        memory[42287] <=  8'h6d;        memory[42288] <=  8'h62;        memory[42289] <=  8'h76;        memory[42290] <=  8'h78;        memory[42291] <=  8'h63;        memory[42292] <=  8'h73;        memory[42293] <=  8'h66;        memory[42294] <=  8'h72;        memory[42295] <=  8'h74;        memory[42296] <=  8'h79;        memory[42297] <=  8'h75;        memory[42298] <=  8'h6a;        memory[42299] <=  8'h6e;        memory[42300] <=  8'h62;        memory[42301] <=  8'h76;        memory[42302] <=  8'h63;        memory[42303] <=  8'h64;        memory[42304] <=  8'h74;        memory[42305] <=  8'h79;        memory[42306] <=  8'h75;        memory[42307] <=  8'h69;        memory[42308] <=  8'h6b;        memory[42309] <=  8'h6d;        memory[42310] <=  8'h6e;        memory[42311] <=  8'h62;        memory[42312] <=  8'h76;        memory[42313] <=  8'h63;        memory[42314] <=  8'h78;        memory[42315] <=  8'h73;        memory[42316] <=  8'h64;        memory[42317] <=  8'h72;        memory[42318] <=  8'h74;        memory[42319] <=  8'h79;        memory[42320] <=  8'h75;        memory[42321] <=  8'h69;        memory[42322] <=  8'h6b;        memory[42323] <=  8'h6d;        memory[42324] <=  8'h6e;        memory[42325] <=  8'h62;        memory[42326] <=  8'h76;        memory[42327] <=  8'h63;        memory[42328] <=  8'h73;        memory[42329] <=  8'h77;        memory[42330] <=  8'h33;        memory[42331] <=  8'h34;        memory[42332] <=  8'h35;        memory[42333] <=  8'h36;        memory[42334] <=  8'h37;        memory[42335] <=  8'h38;        memory[42336] <=  8'h69;        memory[42337] <=  8'h6b;        memory[42338] <=  8'h6d;        memory[42339] <=  8'h6e;        memory[42340] <=  8'h62;        memory[42341] <=  8'h76;        memory[42342] <=  8'h63;        memory[42343] <=  8'h64;        memory[42344] <=  8'h65;        memory[42345] <=  8'h72;        memory[42346] <=  8'h36;        memory[42347] <=  8'h37;        memory[42348] <=  8'h38;        memory[42349] <=  8'h69;        memory[42350] <=  8'h6f;        memory[42351] <=  8'h6b;        memory[42352] <=  8'h6a;        memory[42353] <=  8'h6e;        memory[42354] <=  8'h62;        memory[42355] <=  8'h76;        memory[42356] <=  8'h63;        memory[42357] <=  8'h64;        memory[42358] <=  8'h72;        memory[42359] <=  8'h74;        memory[42360] <=  8'h79;        memory[42361] <=  8'h75;        memory[42362] <=  8'h73;        memory[42363] <=  8'h6a;        memory[42364] <=  8'h63;        memory[42365] <=  8'h6e;        memory[42366] <=  8'h62;        memory[42367] <=  8'h64;        memory[42368] <=  8'h66;        memory[42369] <=  8'h73;        memory[42370] <=  8'h74;        memory[42371] <=  8'h79;        memory[42372] <=  8'h75;        memory[42373] <=  8'h61;        memory[42374] <=  8'h69;        memory[42375] <=  8'h6b;        memory[42376] <=  8'h78;        memory[42377] <=  8'h6d;        memory[42378] <=  8'h6e;        memory[42379] <=  8'h73;        memory[42380] <=  8'h6a;        memory[42381] <=  8'h6f;        memory[42382] <=  8'h64;        memory[42383] <=  8'h6c;        memory[42384] <=  8'h63;        memory[42385] <=  8'h78;        memory[42386] <=  8'h62;        memory[42387] <=  8'h61;        memory[42388] <=  8'h72;        memory[42389] <=  8'h74;        memory[42390] <=  8'h78;        memory[42391] <=  8'h61;        memory[42392] <=  8'h74;        memory[42393] <=  8'h6b;        memory[42394] <=  8'h73;        memory[42395] <=  8'h68;        memory[42396] <=  8'h63;        memory[42397] <=  8'h66;        memory[42398] <=  8'h69;        memory[42399] <=  8'h77;        memory[42400] <=  8'h68;        memory[42401] <=  8'h61;        memory[42402] <=  8'h74;        memory[42403] <=  8'h61;        memory[42404] <=  8'h6e;        memory[42405] <=  8'h61;        memory[42406] <=  8'h62;        memory[42407] <=  8'h61;        memory[42408] <=  8'h63;        memory[42409] <=  8'h61;        memory[42410] <=  8'h74;        memory[42411] <=  8'h61;        memory[42412] <=  8'h62;        memory[42413] <=  8'h61;        memory[42414] <=  8'h72;        memory[42415] <=  8'h63;        memory[42416] <=  8'h61;        memory[42417] <=  8'h68;        memory[42418] <=  8'h64;        memory[42419] <=  8'h75;        memory[42420] <=  8'h63;        memory[42421] <=  8'h74;        memory[42422] <=  8'h61;        memory[42423] <=  8'h64;        memory[42424] <=  8'h61;        memory[42425] <=  8'h61;        memory[42426] <=  8'h63;        memory[42427] <=  8'h61;        memory[42428] <=  8'h72;        memory[42429] <=  8'h62;        memory[42430] <=  8'h61;        memory[42431] <=  8'h72;        memory[42432] <=  8'h74;        memory[42433] <=  8'h78;        memory[42434] <=  8'h61;        memory[42435] <=  8'h74;        memory[42436] <=  8'h6b;        memory[42437] <=  8'h73;        memory[42438] <=  8'h68;        memory[42439] <=  8'h63;        memory[42440] <=  8'h66;        memory[42441] <=  8'h69;        memory[42442] <=  8'h77;        memory[42443] <=  8'h68;        memory[42444] <=  8'h61;        memory[42445] <=  8'h74;        memory[42446] <=  8'h61;        memory[42447] <=  8'h6e;        memory[42448] <=  8'h61;        memory[42449] <=  8'h62;        memory[42450] <=  8'h61;        memory[42451] <=  8'h63;        memory[42452] <=  8'h61;        memory[42453] <=  8'h74;        memory[42454] <=  8'h61;        memory[42455] <=  8'h62;        memory[42456] <=  8'h61;        memory[42457] <=  8'h72;        memory[42458] <=  8'h63;        memory[42459] <=  8'h61;        memory[42460] <=  8'h68;        memory[42461] <=  8'h64;        memory[42462] <=  8'h75;        memory[42463] <=  8'h63;        memory[42464] <=  8'h74;        memory[42465] <=  8'h61;        memory[42466] <=  8'h64;        memory[42467] <=  8'h61;        memory[42468] <=  8'h61;        memory[42469] <=  8'h63;        memory[42470] <=  8'h61;        memory[42471] <=  8'h72;        memory[42472] <=  8'h62;        memory[42473] <=  8'h61;        memory[42474] <=  8'h72;        memory[42475] <=  8'h74;        memory[42476] <=  8'h78;        memory[42477] <=  8'h61;        memory[42478] <=  8'h74;        memory[42479] <=  8'h6b;        memory[42480] <=  8'h73;        memory[42481] <=  8'h68;        memory[42482] <=  8'h63;        memory[42483] <=  8'h66;        memory[42484] <=  8'h69;        memory[42485] <=  8'h77;        memory[42486] <=  8'h68;        memory[42487] <=  8'h61;        memory[42488] <=  8'h74;        memory[42489] <=  8'h61;        memory[42490] <=  8'h6e;        memory[42491] <=  8'h61;        memory[42492] <=  8'h62;        memory[42493] <=  8'h61;        memory[42494] <=  8'h63;        memory[42495] <=  8'h61;        memory[42496] <=  8'h74;        memory[42497] <=  8'h61;        memory[42498] <=  8'h62;        memory[42499] <=  8'h61;        memory[42500] <=  8'h72;        memory[42501] <=  8'h63;        memory[42502] <=  8'h61;        memory[42503] <=  8'h68;        memory[42504] <=  8'h64;        memory[42505] <=  8'h75;        memory[42506] <=  8'h63;        memory[42507] <=  8'h74;        memory[42508] <=  8'h61;        memory[42509] <=  8'h64;        memory[42510] <=  8'h61;        memory[42511] <=  8'h61;        memory[42512] <=  8'h63;        memory[42513] <=  8'h61;        memory[42514] <=  8'h72;        memory[42515] <=  8'h62;        memory[42516] <=  8'h61;        memory[42517] <=  8'h72;        memory[42518] <=  8'h74;        memory[42519] <=  8'h78;        memory[42520] <=  8'h61;        memory[42521] <=  8'h74;        memory[42522] <=  8'h6b;        memory[42523] <=  8'h73;        memory[42524] <=  8'h68;        memory[42525] <=  8'h63;        memory[42526] <=  8'h66;        memory[42527] <=  8'h69;        memory[42528] <=  8'h77;        memory[42529] <=  8'h68;        memory[42530] <=  8'h61;        memory[42531] <=  8'h74;        memory[42532] <=  8'h61;        memory[42533] <=  8'h6e;        memory[42534] <=  8'h61;        memory[42535] <=  8'h62;        memory[42536] <=  8'h61;        memory[42537] <=  8'h63;        memory[42538] <=  8'h61;        memory[42539] <=  8'h74;        memory[42540] <=  8'h61;        memory[42541] <=  8'h62;        memory[42542] <=  8'h61;        memory[42543] <=  8'h72;        memory[42544] <=  8'h63;        memory[42545] <=  8'h61;        memory[42546] <=  8'h68;        memory[42547] <=  8'h64;        memory[42548] <=  8'h75;        memory[42549] <=  8'h63;        memory[42550] <=  8'h74;        memory[42551] <=  8'h61;        memory[42552] <=  8'h64;        memory[42553] <=  8'h61;        memory[42554] <=  8'h61;        memory[42555] <=  8'h63;        memory[42556] <=  8'h61;        memory[42557] <=  8'h72;        memory[42558] <=  8'h62;        memory[42559] <=  8'h61;        memory[42560] <=  8'h72;        memory[42561] <=  8'h74;        memory[42562] <=  8'h78;        memory[42563] <=  8'h61;        memory[42564] <=  8'h74;        memory[42565] <=  8'h6b;        memory[42566] <=  8'h73;        memory[42567] <=  8'h68;        memory[42568] <=  8'h63;        memory[42569] <=  8'h66;        memory[42570] <=  8'h69;        memory[42571] <=  8'h77;        memory[42572] <=  8'h68;        memory[42573] <=  8'h61;        memory[42574] <=  8'h74;        memory[42575] <=  8'h61;        memory[42576] <=  8'h6e;        memory[42577] <=  8'h61;        memory[42578] <=  8'h62;        memory[42579] <=  8'h61;        memory[42580] <=  8'h63;        memory[42581] <=  8'h61;        memory[42582] <=  8'h74;        memory[42583] <=  8'h61;        memory[42584] <=  8'h62;        memory[42585] <=  8'h61;        memory[42586] <=  8'h72;        memory[42587] <=  8'h63;        memory[42588] <=  8'h61;        memory[42589] <=  8'h68;        memory[42590] <=  8'h64;        memory[42591] <=  8'h75;        memory[42592] <=  8'h63;        memory[42593] <=  8'h74;        memory[42594] <=  8'h61;        memory[42595] <=  8'h64;        memory[42596] <=  8'h61;        memory[42597] <=  8'h61;        memory[42598] <=  8'h63;        memory[42599] <=  8'h61;        memory[42600] <=  8'h72;        memory[42601] <=  8'h62;        memory[42602] <=  8'h61;        memory[42603] <=  8'h72;        memory[42604] <=  8'h74;        memory[42605] <=  8'h78;        memory[42606] <=  8'h61;        memory[42607] <=  8'h74;        memory[42608] <=  8'h6b;        memory[42609] <=  8'h73;        memory[42610] <=  8'h68;        memory[42611] <=  8'h63;        memory[42612] <=  8'h66;        memory[42613] <=  8'h69;        memory[42614] <=  8'h77;        memory[42615] <=  8'h68;        memory[42616] <=  8'h61;        memory[42617] <=  8'h74;        memory[42618] <=  8'h61;        memory[42619] <=  8'h6e;        memory[42620] <=  8'h61;        memory[42621] <=  8'h62;        memory[42622] <=  8'h61;        memory[42623] <=  8'h63;        memory[42624] <=  8'h61;        memory[42625] <=  8'h74;        memory[42626] <=  8'h61;        memory[42627] <=  8'h62;        memory[42628] <=  8'h61;        memory[42629] <=  8'h72;        memory[42630] <=  8'h63;        memory[42631] <=  8'h61;        memory[42632] <=  8'h68;        memory[42633] <=  8'h64;        memory[42634] <=  8'h75;        memory[42635] <=  8'h63;        memory[42636] <=  8'h74;        memory[42637] <=  8'h61;        memory[42638] <=  8'h64;        memory[42639] <=  8'h61;        memory[42640] <=  8'h61;        memory[42641] <=  8'h63;        memory[42642] <=  8'h61;        memory[42643] <=  8'h72;        memory[42644] <=  8'h62;        memory[42645] <=  8'h61;        memory[42646] <=  8'h72;        memory[42647] <=  8'h74;        memory[42648] <=  8'h78;        memory[42649] <=  8'h61;        memory[42650] <=  8'h74;        memory[42651] <=  8'h6b;        memory[42652] <=  8'h73;        memory[42653] <=  8'h68;        memory[42654] <=  8'h63;        memory[42655] <=  8'h66;        memory[42656] <=  8'h69;        memory[42657] <=  8'h77;        memory[42658] <=  8'h68;        memory[42659] <=  8'h61;        memory[42660] <=  8'h74;        memory[42661] <=  8'h61;        memory[42662] <=  8'h6e;        memory[42663] <=  8'h61;        memory[42664] <=  8'h62;        memory[42665] <=  8'h61;        memory[42666] <=  8'h63;        memory[42667] <=  8'h61;        memory[42668] <=  8'h74;        memory[42669] <=  8'h61;        memory[42670] <=  8'h62;        memory[42671] <=  8'h61;        memory[42672] <=  8'h72;        memory[42673] <=  8'h63;        memory[42674] <=  8'h61;        memory[42675] <=  8'h68;        memory[42676] <=  8'h64;        memory[42677] <=  8'h75;        memory[42678] <=  8'h63;        memory[42679] <=  8'h74;        memory[42680] <=  8'h61;        memory[42681] <=  8'h64;        memory[42682] <=  8'h61;        memory[42683] <=  8'h61;        memory[42684] <=  8'h63;        memory[42685] <=  8'h61;        memory[42686] <=  8'h72;        memory[42687] <=  8'h62;        memory[42688] <=  8'h61;        memory[42689] <=  8'h72;        memory[42690] <=  8'h74;        memory[42691] <=  8'h78;        memory[42692] <=  8'h61;        memory[42693] <=  8'h74;        memory[42694] <=  8'h6b;        memory[42695] <=  8'h73;        memory[42696] <=  8'h68;        memory[42697] <=  8'h63;        memory[42698] <=  8'h66;        memory[42699] <=  8'h69;        memory[42700] <=  8'h77;        memory[42701] <=  8'h68;        memory[42702] <=  8'h61;        memory[42703] <=  8'h74;        memory[42704] <=  8'h61;        memory[42705] <=  8'h6e;        memory[42706] <=  8'h61;        memory[42707] <=  8'h62;        memory[42708] <=  8'h61;        memory[42709] <=  8'h63;        memory[42710] <=  8'h61;        memory[42711] <=  8'h74;        memory[42712] <=  8'h61;        memory[42713] <=  8'h62;        memory[42714] <=  8'h61;        memory[42715] <=  8'h72;        memory[42716] <=  8'h63;        memory[42717] <=  8'h61;        memory[42718] <=  8'h68;        memory[42719] <=  8'h64;        memory[42720] <=  8'h75;        memory[42721] <=  8'h63;        memory[42722] <=  8'h74;        memory[42723] <=  8'h61;        memory[42724] <=  8'h64;        memory[42725] <=  8'h61;        memory[42726] <=  8'h61;        memory[42727] <=  8'h63;        memory[42728] <=  8'h61;        memory[42729] <=  8'h72;        memory[42730] <=  8'h62;        memory[42731] <=  8'h61;        memory[42732] <=  8'h72;        memory[42733] <=  8'h74;        memory[42734] <=  8'h78;        memory[42735] <=  8'h61;        memory[42736] <=  8'h74;        memory[42737] <=  8'h6b;        memory[42738] <=  8'h73;        memory[42739] <=  8'h68;        memory[42740] <=  8'h63;        memory[42741] <=  8'h66;        memory[42742] <=  8'h69;        memory[42743] <=  8'h77;        memory[42744] <=  8'h68;        memory[42745] <=  8'h61;        memory[42746] <=  8'h74;        memory[42747] <=  8'h61;        memory[42748] <=  8'h6e;        memory[42749] <=  8'h61;        memory[42750] <=  8'h62;        memory[42751] <=  8'h61;        memory[42752] <=  8'h63;        memory[42753] <=  8'h61;        memory[42754] <=  8'h74;        memory[42755] <=  8'h61;        memory[42756] <=  8'h62;        memory[42757] <=  8'h61;        memory[42758] <=  8'h72;        memory[42759] <=  8'h63;        memory[42760] <=  8'h61;        memory[42761] <=  8'h68;        memory[42762] <=  8'h64;        memory[42763] <=  8'h75;        memory[42764] <=  8'h63;        memory[42765] <=  8'h74;        memory[42766] <=  8'h61;        memory[42767] <=  8'h64;        memory[42768] <=  8'h61;        memory[42769] <=  8'h61;        memory[42770] <=  8'h63;        memory[42771] <=  8'h61;        memory[42772] <=  8'h72;        memory[42773] <=  8'h62;        memory[42774] <=  8'h61;        memory[42775] <=  8'h72;        memory[42776] <=  8'h74;        memory[42777] <=  8'h74;        memory[42778] <=  8'h62;        memory[42779] <=  8'h61;        memory[42780] <=  8'h72;        memory[42781] <=  8'h74;        memory[42782] <=  8'h78;        memory[42783] <=  8'h61;        memory[42784] <=  8'h74;        memory[42785] <=  8'h6b;        memory[42786] <=  8'h73;        memory[42787] <=  8'h68;        memory[42788] <=  8'h63;        memory[42789] <=  8'h66;        memory[42790] <=  8'h69;        memory[42791] <=  8'h77;        memory[42792] <=  8'h68;        memory[42793] <=  8'h61;        memory[42794] <=  8'h74;        memory[42795] <=  8'h61;        memory[42796] <=  8'h6e;        memory[42797] <=  8'h61;        memory[42798] <=  8'h62;        memory[42799] <=  8'h61;        memory[42800] <=  8'h63;        memory[42801] <=  8'h61;        memory[42802] <=  8'h74;        memory[42803] <=  8'h61;        memory[42804] <=  8'h62;        memory[42805] <=  8'h61;        memory[42806] <=  8'h72;        memory[42807] <=  8'h63;        memory[42808] <=  8'h61;        memory[42809] <=  8'h68;        memory[42810] <=  8'h64;        memory[42811] <=  8'h75;        memory[42812] <=  8'h63;        memory[42813] <=  8'h74;        memory[42814] <=  8'h61;        memory[42815] <=  8'h64;        memory[42816] <=  8'h61;        memory[42817] <=  8'h61;        memory[42818] <=  8'h63;        memory[42819] <=  8'h61;        memory[42820] <=  8'h72;        memory[42821] <=  8'h63;        memory[42822] <=  8'h74;        memory[42823] <=  8'h72;        memory[42824] <=  8'h63;        memory[42825] <=  8'h61;        memory[42826] <=  8'h74;        memory[42827] <=  8'h72;        memory[42828] <=  8'h63;        memory[42829] <=  8'h61;        memory[42830] <=  8'h74;        memory[42831] <=  8'h63;        memory[42832] <=  8'h62;        memory[42833] <=  8'h61;        memory[42834] <=  8'h74;        memory[42835] <=  8'h62;        memory[42836] <=  8'h72;        memory[42837] <=  8'h63;        memory[42838] <=  8'h61;        memory[42839] <=  8'h72;        memory[42840] <=  8'h62;        memory[42841] <=  8'h78;        memory[42842] <=  8'h74;        memory[42843] <=  8'h61;        memory[42844] <=  8'h72;        memory[42845] <=  8'h64;        memory[42846] <=  8'h66;        memory[42847] <=  8'h73;        memory[42848] <=  8'h67;        memory[42849] <=  8'h76;        memory[42850] <=  8'h68;        memory[42851] <=  8'h62;        memory[42852] <=  8'h6b;        memory[42853] <=  8'h6a;        memory[42854] <=  8'h6e;        memory[42855] <=  8'h6d;        memory[42856] <=  8'h62;        memory[42857] <=  8'h76;        memory[42858] <=  8'h78;        memory[42859] <=  8'h63;        memory[42860] <=  8'h73;        memory[42861] <=  8'h66;        memory[42862] <=  8'h72;        memory[42863] <=  8'h74;        memory[42864] <=  8'h79;        memory[42865] <=  8'h75;        memory[42866] <=  8'h6a;        memory[42867] <=  8'h6e;        memory[42868] <=  8'h62;        memory[42869] <=  8'h76;        memory[42870] <=  8'h63;        memory[42871] <=  8'h64;        memory[42872] <=  8'h74;        memory[42873] <=  8'h79;        memory[42874] <=  8'h75;        memory[42875] <=  8'h69;        memory[42876] <=  8'h6b;        memory[42877] <=  8'h6d;        memory[42878] <=  8'h6e;        memory[42879] <=  8'h62;        memory[42880] <=  8'h76;        memory[42881] <=  8'h63;        memory[42882] <=  8'h78;        memory[42883] <=  8'h73;        memory[42884] <=  8'h64;        memory[42885] <=  8'h72;        memory[42886] <=  8'h74;        memory[42887] <=  8'h79;        memory[42888] <=  8'h75;        memory[42889] <=  8'h69;        memory[42890] <=  8'h6b;        memory[42891] <=  8'h6d;        memory[42892] <=  8'h6e;        memory[42893] <=  8'h62;        memory[42894] <=  8'h76;        memory[42895] <=  8'h63;        memory[42896] <=  8'h73;        memory[42897] <=  8'h77;        memory[42898] <=  8'h33;        memory[42899] <=  8'h34;        memory[42900] <=  8'h35;        memory[42901] <=  8'h36;        memory[42902] <=  8'h37;        memory[42903] <=  8'h38;        memory[42904] <=  8'h69;        memory[42905] <=  8'h6b;        memory[42906] <=  8'h6d;        memory[42907] <=  8'h6e;        memory[42908] <=  8'h62;        memory[42909] <=  8'h76;        memory[42910] <=  8'h63;        memory[42911] <=  8'h64;        memory[42912] <=  8'h65;        memory[42913] <=  8'h72;        memory[42914] <=  8'h36;        memory[42915] <=  8'h37;        memory[42916] <=  8'h38;        memory[42917] <=  8'h69;        memory[42918] <=  8'h6f;        memory[42919] <=  8'h6b;        memory[42920] <=  8'h6a;        memory[42921] <=  8'h6e;        memory[42922] <=  8'h62;        memory[42923] <=  8'h76;        memory[42924] <=  8'h63;        memory[42925] <=  8'h64;        memory[42926] <=  8'h72;        memory[42927] <=  8'h74;        memory[42928] <=  8'h79;        memory[42929] <=  8'h75;        memory[42930] <=  8'h73;        memory[42931] <=  8'h6a;        memory[42932] <=  8'h63;        memory[42933] <=  8'h6e;        memory[42934] <=  8'h62;        memory[42935] <=  8'h64;        memory[42936] <=  8'h66;        memory[42937] <=  8'h73;        memory[42938] <=  8'h74;        memory[42939] <=  8'h79;        memory[42940] <=  8'h75;        memory[42941] <=  8'h61;        memory[42942] <=  8'h69;        memory[42943] <=  8'h6b;        memory[42944] <=  8'h78;        memory[42945] <=  8'h6d;        memory[42946] <=  8'h6e;        memory[42947] <=  8'h73;        memory[42948] <=  8'h6a;        memory[42949] <=  8'h6f;        memory[42950] <=  8'h64;        memory[42951] <=  8'h6c;        memory[42952] <=  8'h63;        memory[42953] <=  8'h78;        memory[42954] <=  8'h2c;        memory[42955] <=  8'h6d;        memory[42956] <=  8'h73;        memory[42957] <=  8'h6b;        memory[42958] <=  8'h64;        memory[42959] <=  8'h6c;        memory[42960] <=  8'h70;        memory[42961] <=  8'h5b;        memory[42962] <=  8'h3b;        memory[42963] <=  8'h73;        memory[42964] <=  8'h6c;        memory[42965] <=  8'h64;        memory[42966] <=  8'h70;        memory[42967] <=  8'h76;        memory[42968] <=  8'h63;        memory[42969] <=  8'h5b;        memory[42970] <=  8'h78;        memory[42971] <=  8'h76;        memory[42972] <=  8'h63;        memory[42973] <=  8'h5b;        memory[42974] <=  8'h78;        memory[42975] <=  8'h70;        memory[42976] <=  8'h6f;        memory[42977] <=  8'h20;        memory[42978] <=  8'h62;        memory[42979] <=  8'h61;        memory[42980] <=  8'h72;        memory[42981] <=  8'h74;        memory[42982] <=  8'h74;        memory[42983] <=  8'h62;        memory[42984] <=  8'h61;        memory[42985] <=  8'h72;        memory[42986] <=  8'h74;        memory[42987] <=  8'h78;        memory[42988] <=  8'h61;        memory[42989] <=  8'h74;        memory[42990] <=  8'h6b;        memory[42991] <=  8'h73;        memory[42992] <=  8'h68;        memory[42993] <=  8'h63;        memory[42994] <=  8'h66;        memory[42995] <=  8'h69;        memory[42996] <=  8'h77;        memory[42997] <=  8'h68;        memory[42998] <=  8'h61;        memory[42999] <=  8'h69;        memory[43000] <=  8'h6a;        memory[43001] <=  8'h78;        memory[43002] <=  8'h5d;        memory[43003] <=  8'h65;        memory[43004] <=  8'h6b;        memory[43005] <=  8'h6f;        memory[43006] <=  8'h39;        memory[43007] <=  8'h64;        memory[43008] <=  8'h75;        memory[43009] <=  8'h38;        memory[43010] <=  8'h79;        memory[43011] <=  8'h20;        memory[43012] <=  8'h37;        memory[43013] <=  8'h63;        memory[43014] <=  8'h67;        memory[43015] <=  8'h78;        memory[43016] <=  8'h63;        memory[43017] <=  8'h75;        memory[43018] <=  8'h68;        memory[43019] <=  8'h69;        memory[43020] <=  8'h6a;        memory[43021] <=  8'h77;        memory[43022] <=  8'h69;        memory[43023] <=  8'h64;        memory[43024] <=  8'h66;        memory[43025] <=  8'h68;        memory[43026] <=  8'h75;        memory[43027] <=  8'h76;        memory[43028] <=  8'h64;        memory[43029] <=  8'h62;        memory[43030] <=  8'h66;        memory[43031] <=  8'h6a;        memory[43032] <=  8'h6e;        memory[43033] <=  8'h6b;        memory[43034] <=  8'h6a;        memory[43035] <=  8'h65;        memory[43036] <=  8'h38;        memory[43037] <=  8'h66;        memory[43038] <=  8'h37;        memory[43039] <=  8'h67;        memory[43040] <=  8'h79;        memory[43041] <=  8'h76;        memory[43042] <=  8'h63;        memory[43043] <=  8'h68;        memory[43044] <=  8'h69;        memory[43045] <=  8'h6a;        memory[43046] <=  8'h33;        memory[43047] <=  8'h65;        memory[43048] <=  8'h67;        memory[43049] <=  8'h79;        memory[43050] <=  8'h72;        memory[43051] <=  8'h64;        memory[43052] <=  8'h62;        memory[43053] <=  8'h6e;        memory[43054] <=  8'h63;        memory[43055] <=  8'h7a;        memory[43056] <=  8'h6a;        memory[43057] <=  8'h6f;        memory[43058] <=  8'h66;        memory[43059] <=  8'h78;        memory[43060] <=  8'h6a;        memory[43061] <=  8'h69;        memory[43062] <=  8'h63;        memory[43063] <=  8'h68;        memory[43064] <=  8'h62;        memory[43065] <=  8'h6e;        memory[43066] <=  8'h6d;        memory[43067] <=  8'h63;        memory[43068] <=  8'h73;        memory[43069] <=  8'h6c;        memory[43070] <=  8'h6b;        memory[43071] <=  8'h6a;        memory[43072] <=  8'h69;        memory[43073] <=  8'h68;        memory[43074] <=  8'h76;        memory[43075] <=  8'h75;        memory[43076] <=  8'h69;        memory[43077] <=  8'h64;        memory[43078] <=  8'h68;        memory[43079] <=  8'h75;        memory[43080] <=  8'h67;        memory[43081] <=  8'h79;        memory[43082] <=  8'h62;        memory[43083] <=  8'h68;        memory[43084] <=  8'h65;        memory[43085] <=  8'h6a;        memory[43086] <=  8'h72;        memory[43087] <=  8'h6b;        memory[43088] <=  8'h6a;        memory[43089] <=  8'h6f;        memory[43090] <=  8'h64;        memory[43091] <=  8'h67;        memory[43092] <=  8'h69;        memory[43093] <=  8'h75;        memory[43094] <=  8'h69;        memory[43095] <=  8'h67;        memory[43096] <=  8'h76;        memory[43097] <=  8'h79;        memory[43098] <=  8'h75;        memory[43099] <=  8'h67;        memory[43100] <=  8'h78;        memory[43101] <=  8'h68;        memory[43102] <=  8'h63;        memory[43103] <=  8'h20;        memory[43104] <=  8'h20;        memory[43105] <=  8'h20;        memory[43106] <=  8'h78;        memory[43107] <=  8'h76;        memory[43108] <=  8'h20;        memory[43109] <=  8'h63;        memory[43110] <=  8'h78;        memory[43111] <=  8'h67;        memory[43112] <=  8'h79;        memory[43113] <=  8'h63;        memory[43114] <=  8'h75;        memory[43115] <=  8'h68;        memory[43116] <=  8'h6a;        memory[43117] <=  8'h6b;        memory[43118] <=  8'h61;        memory[43119] <=  8'h6c;        memory[43120] <=  8'h78;        memory[43121] <=  8'h76;        memory[43122] <=  8'h70;        memory[43123] <=  8'h6f;        memory[43124] <=  8'h69;        memory[43125] <=  8'h6a;        memory[43126] <=  8'h69;        memory[43127] <=  8'h68;        memory[43128] <=  8'h6a;        memory[43129] <=  8'h62;        memory[43130] <=  8'h77;        memory[43131] <=  8'h65;        memory[43132] <=  8'h6e;        memory[43133] <=  8'h61;        memory[43134] <=  8'h66;        memory[43135] <=  8'h6d;        memory[43136] <=  8'h64;        memory[43137] <=  8'h6b;        memory[43138] <=  8'h6d;        memory[43139] <=  8'h76;        memory[43140] <=  8'h6c;        memory[43141] <=  8'h63;        memory[43142] <=  8'h6f;        memory[43143] <=  8'h64;        memory[43144] <=  8'h69;        memory[43145] <=  8'h75;        memory[43146] <=  8'h68;        memory[43147] <=  8'h73;        memory[43148] <=  8'h66;        memory[43149] <=  8'h65;        memory[43150] <=  8'h62;        memory[43151] <=  8'h6e;        memory[43152] <=  8'h64;        memory[43153] <=  8'h73;        memory[43154] <=  8'h63;        memory[43155] <=  8'h6b;        memory[43156] <=  8'h20;        memory[43157] <=  8'h78;        memory[43158] <=  8'h6a;        memory[43159] <=  8'h78;        memory[43160] <=  8'h63;        memory[43161] <=  8'h73;        memory[43162] <=  8'h64;        memory[43163] <=  8'h66;        memory[43164] <=  8'h6b;        memory[43165] <=  8'h64;        memory[43166] <=  8'h6e;        memory[43167] <=  8'h6d;        memory[43168] <=  8'h64;        memory[43169] <=  8'h73;        memory[43170] <=  8'h63;        memory[43171] <=  8'h6b;        memory[43172] <=  8'h78;        memory[43173] <=  8'h6c;        memory[43174] <=  8'h6f;        memory[43175] <=  8'h66;        memory[43176] <=  8'h6a;        memory[43177] <=  8'h69;        memory[43178] <=  8'h61;        memory[43179] <=  8'h62;        memory[43180] <=  8'h6e;        memory[43181] <=  8'h20;        memory[43182] <=  8'h78;        memory[43183] <=  8'h6b;        memory[43184] <=  8'h6d;        memory[43185] <=  8'h20;        memory[43186] <=  8'h6f;        memory[43187] <=  8'h63;        memory[43188] <=  8'h76;        memory[43189] <=  8'h73;        memory[43190] <=  8'h64;        memory[43191] <=  8'h69;        memory[43192] <=  8'h66;        memory[43193] <=  8'h68;        memory[43194] <=  8'h65;        memory[43195] <=  8'h71;        memory[43196] <=  8'h6a;        memory[43197] <=  8'h77;        memory[43198] <=  8'h62;        memory[43199] <=  8'h65;        memory[43200] <=  8'h6e;        memory[43201] <=  8'h20;        memory[43202] <=  8'h6d;        memory[43203] <=  8'h64;        memory[43204] <=  8'h73;        memory[43205] <=  8'h6c;        memory[43206] <=  8'h76;        memory[43207] <=  8'h6b;        memory[43208] <=  8'h63;        memory[43209] <=  8'h78;        memory[43210] <=  8'h20;        memory[43211] <=  8'h6f;        memory[43212] <=  8'h78;        memory[43213] <=  8'h69;        memory[43214] <=  8'h63;        memory[43215] <=  8'h6a;        memory[43216] <=  8'h76;        memory[43217] <=  8'h64;        memory[43218] <=  8'h66;        memory[43219] <=  8'h65;        memory[43220] <=  8'h71;        memory[43221] <=  8'h6e;        memory[43222] <=  8'h20;        memory[43223] <=  8'h64;        memory[43224] <=  8'h6d;        memory[43225] <=  8'h73;        memory[43226] <=  8'h6c;        memory[43227] <=  8'h63;        memory[43228] <=  8'h78;        memory[43229] <=  8'h6b;        memory[43230] <=  8'h20;        memory[43231] <=  8'h6f;        memory[43232] <=  8'h78;        memory[43233] <=  8'h63;        memory[43234] <=  8'h76;        memory[43235] <=  8'h6a;        memory[43236] <=  8'h64;        memory[43237] <=  8'h62;        memory[43238] <=  8'h71;        memory[43239] <=  8'h77;        memory[43240] <=  8'h65;        memory[43241] <=  8'h6e;        memory[43242] <=  8'h6d;        memory[43243] <=  8'h64;        memory[43244] <=  8'h6c;        memory[43245] <=  8'h73;        memory[43246] <=  8'h2c;        memory[43247] <=  8'h76;        memory[43248] <=  8'h63;        memory[43249] <=  8'h78;        memory[43250] <=  8'h20;        memory[43251] <=  8'h63;        memory[43252] <=  8'h6f;        memory[43253] <=  8'h69;        memory[43254] <=  8'h76;        memory[43255] <=  8'h68;        memory[43256] <=  8'h73;        memory[43257] <=  8'h64;        memory[43258] <=  8'h62;        memory[43259] <=  8'h71;        memory[43260] <=  8'h77;        memory[43261] <=  8'h65;        memory[43262] <=  8'h6e;        memory[43263] <=  8'h64;        memory[43264] <=  8'h6b;        memory[43265] <=  8'h73;        memory[43266] <=  8'h76;        memory[43267] <=  8'h6f;        memory[43268] <=  8'h63;        memory[43269] <=  8'h20;        memory[43270] <=  8'h76;        memory[43271] <=  8'h69;        memory[43272] <=  8'h75;        memory[43273] <=  8'h69;        memory[43274] <=  8'h68;        memory[43275] <=  8'h63;        memory[43276] <=  8'h78;        memory[43277] <=  8'h69;        memory[43278] <=  8'h6f;        memory[43279] <=  8'h76;        memory[43280] <=  8'h73;        memory[43281] <=  8'h64;        memory[43282] <=  8'h61;        memory[43283] <=  8'h64;        memory[43284] <=  8'h6e;        memory[43285] <=  8'h77;        memory[43286] <=  8'h71;        memory[43287] <=  8'h6b;        memory[43288] <=  8'h6c;        memory[43289] <=  8'h73;        memory[43290] <=  8'h76;        memory[43291] <=  8'h6e;        memory[43292] <=  8'h62;        memory[43293] <=  8'h20;        memory[43294] <=  8'h64;        memory[43295] <=  8'h66;        memory[43296] <=  8'h6a;        memory[43297] <=  8'h6b;        memory[43298] <=  8'h71;        memory[43299] <=  8'h64;        memory[43300] <=  8'h77;        memory[43301] <=  8'h65;        memory[43302] <=  8'h6e;        memory[43303] <=  8'h62;        memory[43304] <=  8'h20;        memory[43305] <=  8'h64;        memory[43306] <=  8'h73;        memory[43307] <=  8'h76;        memory[43308] <=  8'h68;        memory[43309] <=  8'h64;        memory[43310] <=  8'h61;        memory[43311] <=  8'h71;        memory[43312] <=  8'h77;        memory[43313] <=  8'h6a;        memory[43314] <=  8'h65;        memory[43315] <=  8'h6e;        memory[43316] <=  8'h64;        memory[43317] <=  8'h20;        memory[43318] <=  8'h61;        memory[43319] <=  8'h63;        memory[43320] <=  8'h62;        memory[43321] <=  8'h68;        memory[43322] <=  8'h64;        memory[43323] <=  8'h61;        memory[43324] <=  8'h77;        memory[43325] <=  8'h71;        memory[43326] <=  8'h6e;        memory[43327] <=  8'h20;        memory[43328] <=  8'h62;        memory[43329] <=  8'h73;        memory[43330] <=  8'h76;        memory[43331] <=  8'h61;        memory[43332] <=  8'h67;        memory[43333] <=  8'h76;        memory[43334] <=  8'h68;        memory[43335] <=  8'h67;        memory[43336] <=  8'h61;        memory[43337] <=  8'h73;        memory[43338] <=  8'h6a;        memory[43339] <=  8'h6b;        memory[43340] <=  8'h63;        memory[43341] <=  8'h78;        memory[43342] <=  8'h76;        memory[43343] <=  8'h6e;        memory[43344] <=  8'h73;        memory[43345] <=  8'h64;        memory[43346] <=  8'h20;        memory[43347] <=  8'h66;        memory[43348] <=  8'h62;        memory[43349] <=  8'h64;        memory[43350] <=  8'h61;        memory[43351] <=  8'h73;        memory[43352] <=  8'h76;        memory[43353] <=  8'h67;        memory[43354] <=  8'h63;        memory[43355] <=  8'h79;        memory[43356] <=  8'h7a;        memory[43357] <=  8'h78;        memory[43358] <=  8'h79;        memory[43359] <=  8'h75;        memory[43360] <=  8'h20;        memory[43361] <=  8'h69;        memory[43362] <=  8'h6a;        memory[43363] <=  8'h64;        memory[43364] <=  8'h66;        memory[43365] <=  8'h6b;        memory[43366] <=  8'h61;        memory[43367] <=  8'h64;        memory[43368] <=  8'h63;        memory[43369] <=  8'h78;        memory[43370] <=  8'h68;        memory[43371] <=  8'h20;        memory[43372] <=  8'h67;        memory[43373] <=  8'h61;        memory[43374] <=  8'h68;        memory[43375] <=  8'h75;        memory[43376] <=  8'h64;        memory[43377] <=  8'h73;        memory[43378] <=  8'h69;        memory[43379] <=  8'h6a;        memory[43380] <=  8'h61;        memory[43381] <=  8'h6b;        memory[43382] <=  8'h63;        memory[43383] <=  8'h62;        memory[43384] <=  8'h61;        memory[43385] <=  8'h72;        memory[43386] <=  8'h73;        memory[43387] <=  8'h68;        memory[43388] <=  8'h64;        memory[43389] <=  8'h66;        memory[43390] <=  8'h67;        memory[43391] <=  8'h73;        memory[43392] <=  8'h68;        memory[43393] <=  8'h64;        memory[43394] <=  8'h66;        memory[43395] <=  8'h68;        memory[43396] <=  8'h64;        memory[43397] <=  8'h6a;        memory[43398] <=  8'h68;        memory[43399] <=  8'h62;        memory[43400] <=  8'h67;        memory[43401] <=  8'h63;        memory[43402] <=  8'h61;        memory[43403] <=  8'h66;        memory[43404] <=  8'h73;        memory[43405] <=  8'h79;        memory[43406] <=  8'h67;        memory[43407] <=  8'h6b;        memory[43408] <=  8'h75;        memory[43409] <=  8'h64;        memory[43410] <=  8'h68;        memory[43411] <=  8'h62;        memory[43412] <=  8'h77;        memory[43413] <=  8'h76;        memory[43414] <=  8'h67;        memory[43415] <=  8'h61;        memory[43416] <=  8'h66;        memory[43417] <=  8'h64;        memory[43418] <=  8'h74;        memory[43419] <=  8'h75;        memory[43420] <=  8'h66;        memory[43421] <=  8'h79;        memory[43422] <=  8'h67;        memory[43423] <=  8'h69;        memory[43424] <=  8'h75;        memory[43425] <=  8'h68;        memory[43426] <=  8'h6c;        memory[43427] <=  8'h6a;        memory[43428] <=  8'h62;        memory[43429] <=  8'h6b;        memory[43430] <=  8'h68;        memory[43431] <=  8'h76;        memory[43432] <=  8'h67;        memory[43433] <=  8'h63;        memory[43434] <=  8'h66;        memory[43435] <=  8'h78;        memory[43436] <=  8'h64;        memory[43437] <=  8'h74;        memory[43438] <=  8'h75;        memory[43439] <=  8'h79;        memory[43440] <=  8'h69;        memory[43441] <=  8'h75;        memory[43442] <=  8'h68;        memory[43443] <=  8'h6c;        memory[43444] <=  8'h6a;        memory[43445] <=  8'h6b;        memory[43446] <=  8'h67;        memory[43447] <=  8'h6a;        memory[43448] <=  8'h63;        memory[43449] <=  8'h66;        memory[43450] <=  8'h68;        memory[43451] <=  8'h64;        memory[43452] <=  8'h67;        memory[43453] <=  8'h72;        memory[43454] <=  8'h79;        memory[43455] <=  8'h74;        memory[43456] <=  8'h66;        memory[43457] <=  8'h75;        memory[43458] <=  8'h79;        memory[43459] <=  8'h69;        memory[43460] <=  8'h68;        memory[43461] <=  8'h6c;        memory[43462] <=  8'h62;        memory[43463] <=  8'h6d;        memory[43464] <=  8'h76;        memory[43465] <=  8'h6e;        memory[43466] <=  8'h63;        memory[43467] <=  8'h66;        memory[43468] <=  8'h68;        memory[43469] <=  8'h64;        memory[43470] <=  8'h74;        memory[43471] <=  8'h75;        memory[43472] <=  8'h67;        memory[43473] <=  8'h79;        memory[43474] <=  8'h69;        memory[43475] <=  8'h68;        memory[43476] <=  8'h75;        memory[43477] <=  8'h6a;        memory[43478] <=  8'h6c;        memory[43479] <=  8'h62;        memory[43480] <=  8'h6d;        memory[43481] <=  8'h76;        memory[43482] <=  8'h6e;        memory[43483] <=  8'h63;        memory[43484] <=  8'h66;        memory[43485] <=  8'h68;        memory[43486] <=  8'h67;        memory[43487] <=  8'h79;        memory[43488] <=  8'h68;        memory[43489] <=  8'h75;        memory[43490] <=  8'h6a;        memory[43491] <=  8'h6e;        memory[43492] <=  8'h2c;        memory[43493] <=  8'h62;        memory[43494] <=  8'h6e;        memory[43495] <=  8'h6d;        memory[43496] <=  8'h76;        memory[43497] <=  8'h6e;        memory[43498] <=  8'h63;        memory[43499] <=  8'h66;        memory[43500] <=  8'h68;        memory[43501] <=  8'h74;        memory[43502] <=  8'h79;        memory[43503] <=  8'h69;        memory[43504] <=  8'h75;        memory[43505] <=  8'h6c;        memory[43506] <=  8'h6a;        memory[43507] <=  8'h62;        memory[43508] <=  8'h6d;        memory[43509] <=  8'h76;        memory[43510] <=  8'h6e;        memory[43511] <=  8'h63;        memory[43512] <=  8'h66;        memory[43513] <=  8'h74;        memory[43514] <=  8'h75;        memory[43515] <=  8'h79;        memory[43516] <=  8'h69;        memory[43517] <=  8'h68;        memory[43518] <=  8'h6b;        memory[43519] <=  8'h62;        memory[43520] <=  8'h76;        memory[43521] <=  8'h63;        memory[43522] <=  8'h66;        memory[43523] <=  8'h67;        memory[43524] <=  8'h74;        memory[43525] <=  8'h75;        memory[43526] <=  8'h79;        memory[43527] <=  8'h69;        memory[43528] <=  8'h75;        memory[43529] <=  8'h68;        memory[43530] <=  8'h6a;        memory[43531] <=  8'h6b;        memory[43532] <=  8'h62;        memory[43533] <=  8'h76;        memory[43534] <=  8'h63;        memory[43535] <=  8'h66;        memory[43536] <=  8'h74;        memory[43537] <=  8'h75;        memory[43538] <=  8'h79;        memory[43539] <=  8'h69;        memory[43540] <=  8'h75;        memory[43541] <=  8'h6a;        memory[43542] <=  8'h6b;        memory[43543] <=  8'h6e;        memory[43544] <=  8'h62;        memory[43545] <=  8'h76;        memory[43546] <=  8'h67;        memory[43547] <=  8'h66;        memory[43548] <=  8'h74;        memory[43549] <=  8'h79;        memory[43550] <=  8'h75;        memory[43551] <=  8'h75;        memory[43552] <=  8'h69;        memory[43553] <=  8'h6a;        memory[43554] <=  8'h6b;        memory[43555] <=  8'h68;        memory[43556] <=  8'h62;        memory[43557] <=  8'h6a;        memory[43558] <=  8'h67;        memory[43559] <=  8'h68;        memory[43560] <=  8'h66;        memory[43561] <=  8'h79;        memory[43562] <=  8'h74;        memory[43563] <=  8'h79;        memory[43564] <=  8'h69;        memory[43565] <=  8'h75;        memory[43566] <=  8'h64;        memory[43567] <=  8'h6a;        memory[43568] <=  8'h6b;        memory[43569] <=  8'h68;        memory[43570] <=  8'h63;        memory[43571] <=  8'h7a;        memory[43572] <=  8'h67;        memory[43573] <=  8'h68;        memory[43574] <=  8'h74;        memory[43575] <=  8'h75;        memory[43576] <=  8'h79;        memory[43577] <=  8'h69;        memory[43578] <=  8'h61;        memory[43579] <=  8'h73;        memory[43580] <=  8'h75;        memory[43581] <=  8'h6a;        memory[43582] <=  8'h6b;        memory[43583] <=  8'h62;        memory[43584] <=  8'h6e;        memory[43585] <=  8'h61;        memory[43586] <=  8'h76;        memory[43587] <=  8'h63;        memory[43588] <=  8'h66;        memory[43589] <=  8'h68;        memory[43590] <=  8'h75;        memory[43591] <=  8'h61;        memory[43592] <=  8'h73;        memory[43593] <=  8'h79;        memory[43594] <=  8'h64;        memory[43595] <=  8'h75;        memory[43596] <=  8'h69;        memory[43597] <=  8'h6a;        memory[43598] <=  8'h61;        memory[43599] <=  8'h6b;        memory[43600] <=  8'h62;        memory[43601] <=  8'h63;        memory[43602] <=  8'h78;        memory[43603] <=  8'h68;        memory[43604] <=  8'h67;        memory[43605] <=  8'h79;        memory[43606] <=  8'h75;        memory[43607] <=  8'h7a;        memory[43608] <=  8'h63;        memory[43609] <=  8'h61;        memory[43610] <=  8'h73;        memory[43611] <=  8'h69;        memory[43612] <=  8'h75;        memory[43613] <=  8'h6f;        memory[43614] <=  8'h69;        memory[43615] <=  8'h6a;        memory[43616] <=  8'h61;        memory[43617] <=  8'h6c;        memory[43618] <=  8'h63;        memory[43619] <=  8'h78;        memory[43620] <=  8'h62;        memory[43621] <=  8'h63;        memory[43622] <=  8'h20;        memory[43623] <=  8'h6e;        memory[43624] <=  8'h76;        memory[43625] <=  8'h63;        memory[43626] <=  8'h61;        memory[43627] <=  8'h64;        memory[43628] <=  8'h73;        memory[43629] <=  8'h67;        memory[43630] <=  8'h79;        memory[43631] <=  8'h68;        memory[43632] <=  8'h75;        memory[43633] <=  8'h61;        memory[43634] <=  8'h6a;        memory[43635] <=  8'h6b;        memory[43636] <=  8'h78;        memory[43637] <=  8'h62;        memory[43638] <=  8'h20;        memory[43639] <=  8'h6e;        memory[43640] <=  8'h76;        memory[43641] <=  8'h63;        memory[43642] <=  8'h61;        memory[43643] <=  8'h73;        memory[43644] <=  8'h67;        memory[43645] <=  8'h68;        memory[43646] <=  8'h75;        memory[43647] <=  8'h6a;        memory[43648] <=  8'h6c;        memory[43649] <=  8'h6b;        memory[43650] <=  8'h63;        memory[43651] <=  8'h78;        memory[43652] <=  8'h20;        memory[43653] <=  8'h6a;        memory[43654] <=  8'h6b;        memory[43655] <=  8'h68;        memory[43656] <=  8'h61;        memory[43657] <=  8'h73;        memory[43658] <=  8'h76;        memory[43659] <=  8'h64;        memory[43660] <=  8'h6e;        memory[43661] <=  8'h20;        memory[43662] <=  8'h62;        memory[43663] <=  8'h6e;        memory[43664] <=  8'h6d;        memory[43665] <=  8'h6b;        memory[43666] <=  8'h77;        memory[43667] <=  8'h64;        memory[43668] <=  8'h6f;        memory[43669] <=  8'h77;        memory[43670] <=  8'h69;        memory[43671] <=  8'h6f;        memory[43672] <=  8'h75;        memory[43673] <=  8'h69;        memory[43674] <=  8'h68;        memory[43675] <=  8'h62;        memory[43676] <=  8'h6e;        memory[43677] <=  8'h6b;        memory[43678] <=  8'h77;        memory[43679] <=  8'h69;        memory[43680] <=  8'h6f;        memory[43681] <=  8'h75;        memory[43682] <=  8'h71;        memory[43683] <=  8'h69;        memory[43684] <=  8'h79;        memory[43685] <=  8'h67;        memory[43686] <=  8'h6a;        memory[43687] <=  8'h64;        memory[43688] <=  8'h61;        memory[43689] <=  8'h76;        memory[43690] <=  8'h62;        memory[43691] <=  8'h6e;        memory[43692] <=  8'h6b;        memory[43693] <=  8'h6f;        memory[43694] <=  8'h70;        memory[43695] <=  8'h64;        memory[43696] <=  8'h76;        memory[43697] <=  8'h69;        memory[43698] <=  8'h6f;        memory[43699] <=  8'h75;        memory[43700] <=  8'h69;        memory[43701] <=  8'h48;        memory[43702] <=  8'h42;        memory[43703] <=  8'h6b;        memory[43704] <=  8'h64;        memory[43705] <=  8'h6e;        memory[43706] <=  8'h6c;        memory[43707] <=  8'h71;        memory[43708] <=  8'h6b;        memory[43709] <=  8'h6d;        memory[43710] <=  8'h6a;        memory[43711] <=  8'h70;        memory[43712] <=  8'h69;        memory[43713] <=  8'h6f;        memory[43714] <=  8'h68;        memory[43715] <=  8'h65;        memory[43716] <=  8'h66;        memory[43717] <=  8'h75;        memory[43718] <=  8'h67;        memory[43719] <=  8'h69;        memory[43720] <=  8'h73;        memory[43721] <=  8'h61;        memory[43722] <=  8'h62;        memory[43723] <=  8'h64;        memory[43724] <=  8'h6b;        memory[43725] <=  8'h6a;        memory[43726] <=  8'h6b;        memory[43727] <=  8'h6c;        memory[43728] <=  8'h6a;        memory[43729] <=  8'h69;        memory[43730] <=  8'h73;        memory[43731] <=  8'h6f;        memory[43732] <=  8'h71;        memory[43733] <=  8'h68;        memory[43734] <=  8'h77;        memory[43735] <=  8'h67;        memory[43736] <=  8'h69;        memory[43737] <=  8'h79;        memory[43738] <=  8'h6a;        memory[43739] <=  8'h64;        memory[43740] <=  8'h76;        memory[43741] <=  8'h62;        memory[43742] <=  8'h6e;        memory[43743] <=  8'h61;        memory[43744] <=  8'h73;        memory[43745] <=  8'h66;        memory[43746] <=  8'h6c;        memory[43747] <=  8'h6b;        memory[43748] <=  8'h64;        memory[43749] <=  8'h6a;        memory[43750] <=  8'h68;        memory[43751] <=  8'h63;        memory[43752] <=  8'h67;        memory[43753] <=  8'h6a;        memory[43754] <=  8'h76;        memory[43755] <=  8'h73;        memory[43756] <=  8'h64;        memory[43757] <=  8'h62;        memory[43758] <=  8'h62;        memory[43759] <=  8'h61;        memory[43760] <=  8'h72;        memory[43761] <=  8'h62;        memory[43762] <=  8'h62;        memory[43763] <=  8'h73;        memory[43764] <=  8'h62;        memory[43765] <=  8'h67;        memory[43766] <=  8'h73;        memory[43767] <=  8'h66;        memory[43768] <=  8'h67;        memory[43769] <=  8'h61;        memory[43770] <=  8'h68;        memory[43771] <=  8'h66;        memory[43772] <=  8'h73;        memory[43773] <=  8'h68;        memory[43774] <=  8'h61;        memory[43775] <=  8'h66;        memory[43776] <=  8'h73;        memory[43777] <=  8'h66;        memory[43778] <=  8'h68;        memory[43779] <=  8'h61;        memory[43780] <=  8'h69;        memory[43781] <=  8'h64;        memory[43782] <=  8'h75;        memory[43783] <=  8'h67;        memory[43784] <=  8'h64;        memory[43785] <=  8'h77;        memory[43786] <=  8'h62;        memory[43787] <=  8'h61;        memory[43788] <=  8'h62;        memory[43789] <=  8'h72;        memory[43790] <=  8'h62;        memory[43791] <=  8'h61;        memory[43792] <=  8'h62;        memory[43793] <=  8'h62;        memory[43794] <=  8'h74;        memory[43795] <=  8'h62;        memory[43796] <=  8'h62;        memory[43797] <=  8'h62;        memory[43798] <=  8'h62;        memory[43799] <=  8'h62;        memory[43800] <=  8'h62;        memory[43801] <=  8'h62;        memory[43802] <=  8'h62;        memory[43803] <=  8'h61;        memory[43804] <=  8'h62;        memory[43805] <=  8'h62;        memory[43806] <=  8'h72;        memory[43807] <=  8'h74;        memory[43808] <=  8'h62;        memory[43809] <=  8'h62;        memory[43810] <=  8'h61;        memory[43811] <=  8'h62;        memory[43812] <=  8'h72;        memory[43813] <=  8'h62;        memory[43814] <=  8'h74;        memory[43815] <=  8'h62;        memory[43816] <=  8'h62;        memory[43817] <=  8'h62;        memory[43818] <=  8'h63;        memory[43819] <=  8'h61;        memory[43820] <=  8'h72;        memory[43821] <=  8'h74;        memory[43822] <=  8'h73;        memory[43823] <=  8'h62;        memory[43824] <=  8'h61;        memory[43825] <=  8'h72;        memory[43826] <=  8'h74;        memory[43827] <=  8'h74;        memory[43828] <=  8'h62;        memory[43829] <=  8'h61;        memory[43830] <=  8'h72;        memory[43831] <=  8'h74;        memory[43832] <=  8'h78;        memory[43833] <=  8'h61;        memory[43834] <=  8'h74;        memory[43835] <=  8'h6b;        memory[43836] <=  8'h73;        memory[43837] <=  8'h68;        memory[43838] <=  8'h63;        memory[43839] <=  8'h66;        memory[43840] <=  8'h69;        memory[43841] <=  8'h77;        memory[43842] <=  8'h68;        memory[43843] <=  8'h61;        memory[43844] <=  8'h74;        memory[43845] <=  8'h61;        memory[43846] <=  8'h6e;        memory[43847] <=  8'h61;        memory[43848] <=  8'h62;        memory[43849] <=  8'h61;        memory[43850] <=  8'h63;        memory[43851] <=  8'h61;        memory[43852] <=  8'h74;        memory[43853] <=  8'h61;        memory[43854] <=  8'h62;        memory[43855] <=  8'h61;        memory[43856] <=  8'h72;        memory[43857] <=  8'h63;        memory[43858] <=  8'h61;        memory[43859] <=  8'h68;        memory[43860] <=  8'h64;        memory[43861] <=  8'h75;        memory[43862] <=  8'h63;        memory[43863] <=  8'h74;        memory[43864] <=  8'h61;        memory[43865] <=  8'h64;        memory[43866] <=  8'h61;        memory[43867] <=  8'h61;        memory[43868] <=  8'h63;        memory[43869] <=  8'h61;        memory[43870] <=  8'h72;        memory[43871] <=  8'h63;        memory[43872] <=  8'h74;        memory[43873] <=  8'h72;        memory[43874] <=  8'h63;        memory[43875] <=  8'h61;        memory[43876] <=  8'h74;        memory[43877] <=  8'h72;        memory[43878] <=  8'h63;        memory[43879] <=  8'h61;        memory[43880] <=  8'h74;        memory[43881] <=  8'h63;        memory[43882] <=  8'h62;        memory[43883] <=  8'h61;        memory[43884] <=  8'h74;        memory[43885] <=  8'h62;        memory[43886] <=  8'h72;        memory[43887] <=  8'h63;        memory[43888] <=  8'h61;        memory[43889] <=  8'h74;        memory[43890] <=  8'h72;        memory[43891] <=  8'h6e;        memory[43892] <=  8'h62;        memory[43893] <=  8'h61;        memory[43894] <=  8'h63;        memory[43895] <=  8'h61;        memory[43896] <=  8'h74;        memory[43897] <=  8'h79;        memory[43898] <=  8'h73;        memory[43899] <=  8'h6e;        memory[43900] <=  8'h63;        memory[43901] <=  8'h74;        memory[43902] <=  8'h61;        memory[43903] <=  8'h6e;        memory[43904] <=  8'h62;        memory[43905] <=  8'h61;        memory[43906] <=  8'h63;        memory[43907] <=  8'h72;        memory[43908] <=  8'h6e;        memory[43909] <=  8'h74;        memory[43910] <=  8'h61;        memory[43911] <=  8'h62;        memory[43912] <=  8'h74;        memory[43913] <=  8'h6e;        memory[43914] <=  8'h61;        memory[43915] <=  8'h72;        memory[43916] <=  8'h62;        memory[43917] <=  8'h78;        memory[43918] <=  8'h74;        memory[43919] <=  8'h61;        memory[43920] <=  8'h72;        memory[43921] <=  8'h62;        memory[43922] <=  8'h61;        memory[43923] <=  8'h72;        memory[43924] <=  8'h74;        memory[43925] <=  8'h74;        memory[43926] <=  8'h62;        memory[43927] <=  8'h61;        memory[43928] <=  8'h72;        memory[43929] <=  8'h74;        memory[43930] <=  8'h78;        memory[43931] <=  8'h61;        memory[43932] <=  8'h74;        memory[43933] <=  8'h6b;        memory[43934] <=  8'h73;        memory[43935] <=  8'h68;        memory[43936] <=  8'h63;        memory[43937] <=  8'h66;        memory[43938] <=  8'h69;        memory[43939] <=  8'h77;        memory[43940] <=  8'h68;        memory[43941] <=  8'h61;        memory[43942] <=  8'h74;        memory[43943] <=  8'h61;        memory[43944] <=  8'h6e;        memory[43945] <=  8'h61;        memory[43946] <=  8'h62;        memory[43947] <=  8'h61;        memory[43948] <=  8'h63;        memory[43949] <=  8'h61;        memory[43950] <=  8'h74;        memory[43951] <=  8'h61;        memory[43952] <=  8'h62;        memory[43953] <=  8'h61;        memory[43954] <=  8'h72;        memory[43955] <=  8'h63;        memory[43956] <=  8'h61;        memory[43957] <=  8'h68;        memory[43958] <=  8'h64;        memory[43959] <=  8'h75;        memory[43960] <=  8'h63;        memory[43961] <=  8'h74;        memory[43962] <=  8'h61;        memory[43963] <=  8'h64;        memory[43964] <=  8'h61;        memory[43965] <=  8'h61;        memory[43966] <=  8'h63;        memory[43967] <=  8'h61;        memory[43968] <=  8'h72;        memory[43969] <=  8'h63;        memory[43970] <=  8'h74;        memory[43971] <=  8'h72;        memory[43972] <=  8'h63;        memory[43973] <=  8'h61;        memory[43974] <=  8'h74;        memory[43975] <=  8'h72;        memory[43976] <=  8'h63;        memory[43977] <=  8'h61;        memory[43978] <=  8'h74;        memory[43979] <=  8'h63;        memory[43980] <=  8'h62;        memory[43981] <=  8'h61;        memory[43982] <=  8'h74;        memory[43983] <=  8'h62;        memory[43984] <=  8'h72;        memory[43985] <=  8'h63;        memory[43986] <=  8'h61;        memory[43987] <=  8'h74;        memory[43988] <=  8'h72;        memory[43989] <=  8'h6e;        memory[43990] <=  8'h62;        memory[43991] <=  8'h61;        memory[43992] <=  8'h63;        memory[43993] <=  8'h61;        memory[43994] <=  8'h74;        memory[43995] <=  8'h79;        memory[43996] <=  8'h73;        memory[43997] <=  8'h6e;        memory[43998] <=  8'h63;        memory[43999] <=  8'h74;        memory[44000] <=  8'h61;        memory[44001] <=  8'h6e;        memory[44002] <=  8'h62;        memory[44003] <=  8'h61;        memory[44004] <=  8'h63;        memory[44005] <=  8'h72;        memory[44006] <=  8'h6e;        memory[44007] <=  8'h74;        memory[44008] <=  8'h61;        memory[44009] <=  8'h62;        memory[44010] <=  8'h74;        memory[44011] <=  8'h6e;        memory[44012] <=  8'h61;        memory[44013] <=  8'h72;        memory[44014] <=  8'h62;        memory[44015] <=  8'h78;        memory[44016] <=  8'h74;        memory[44017] <=  8'h61;        memory[44018] <=  8'h72;        memory[44019] <=  8'h62;        memory[44020] <=  8'h61;        memory[44021] <=  8'h72;        memory[44022] <=  8'h74;        memory[44023] <=  8'h74;        memory[44024] <=  8'h62;        memory[44025] <=  8'h61;        memory[44026] <=  8'h72;        memory[44027] <=  8'h74;        memory[44028] <=  8'h78;        memory[44029] <=  8'h61;        memory[44030] <=  8'h74;        memory[44031] <=  8'h6b;        memory[44032] <=  8'h73;        memory[44033] <=  8'h68;        memory[44034] <=  8'h63;        memory[44035] <=  8'h66;        memory[44036] <=  8'h69;        memory[44037] <=  8'h77;        memory[44038] <=  8'h68;        memory[44039] <=  8'h61;        memory[44040] <=  8'h74;        memory[44041] <=  8'h61;        memory[44042] <=  8'h6e;        memory[44043] <=  8'h61;        memory[44044] <=  8'h62;        memory[44045] <=  8'h61;        memory[44046] <=  8'h63;        memory[44047] <=  8'h61;        memory[44048] <=  8'h74;        memory[44049] <=  8'h61;        memory[44050] <=  8'h62;        memory[44051] <=  8'h61;        memory[44052] <=  8'h72;        memory[44053] <=  8'h63;        memory[44054] <=  8'h61;        memory[44055] <=  8'h68;        memory[44056] <=  8'h64;        memory[44057] <=  8'h75;        memory[44058] <=  8'h63;        memory[44059] <=  8'h74;        memory[44060] <=  8'h61;        memory[44061] <=  8'h64;        memory[44062] <=  8'h61;        memory[44063] <=  8'h61;        memory[44064] <=  8'h63;        memory[44065] <=  8'h61;        memory[44066] <=  8'h72;        memory[44067] <=  8'h63;        memory[44068] <=  8'h74;        memory[44069] <=  8'h72;        memory[44070] <=  8'h63;        memory[44071] <=  8'h61;        memory[44072] <=  8'h74;        memory[44073] <=  8'h72;        memory[44074] <=  8'h63;        memory[44075] <=  8'h61;        memory[44076] <=  8'h74;        memory[44077] <=  8'h63;        memory[44078] <=  8'h62;        memory[44079] <=  8'h61;        memory[44080] <=  8'h74;        memory[44081] <=  8'h62;        memory[44082] <=  8'h72;        memory[44083] <=  8'h63;        memory[44084] <=  8'h61;        memory[44085] <=  8'h74;        memory[44086] <=  8'h72;        memory[44087] <=  8'h6e;        memory[44088] <=  8'h62;        memory[44089] <=  8'h61;        memory[44090] <=  8'h63;        memory[44091] <=  8'h61;        memory[44092] <=  8'h74;        memory[44093] <=  8'h79;        memory[44094] <=  8'h73;        memory[44095] <=  8'h6e;        memory[44096] <=  8'h63;        memory[44097] <=  8'h74;        memory[44098] <=  8'h61;        memory[44099] <=  8'h6e;        memory[44100] <=  8'h62;        memory[44101] <=  8'h61;        memory[44102] <=  8'h63;        memory[44103] <=  8'h72;        memory[44104] <=  8'h6e;        memory[44105] <=  8'h74;        memory[44106] <=  8'h61;        memory[44107] <=  8'h62;        memory[44108] <=  8'h74;        memory[44109] <=  8'h6e;        memory[44110] <=  8'h61;        memory[44111] <=  8'h72;        memory[44112] <=  8'h62;        memory[44113] <=  8'h78;        memory[44114] <=  8'h74;        memory[44115] <=  8'h61;        memory[44116] <=  8'h72;        memory[44117] <=  8'h5d;        memory[44118] <=  8'h5d;        memory[44119] <=  8'h65;        memory[44120] <=  8'h66;        memory[44121] <=  8'h77;        memory[44122] <=  8'h65;        memory[44123] <=  8'h5d;        memory[44124] <=  8'h65;        memory[44125] <=  8'h67;        memory[44126] <=  8'h73;        memory[44127] <=  8'h67;        memory[44128] <=  8'h66;        memory[44129] <=  8'h62;        memory[44130] <=  8'h61;        memory[44131] <=  8'h72;        memory[44132] <=  8'h74;        memory[44133] <=  8'h74;        memory[44134] <=  8'h62;        memory[44135] <=  8'h61;        memory[44136] <=  8'h72;        memory[44137] <=  8'h74;        memory[44138] <=  8'h78;        memory[44139] <=  8'h61;        memory[44140] <=  8'h74;        memory[44141] <=  8'h6b;        memory[44142] <=  8'h73;        memory[44143] <=  8'h68;        memory[44144] <=  8'h63;        memory[44145] <=  8'h66;        memory[44146] <=  8'h69;        memory[44147] <=  8'h77;        memory[44148] <=  8'h68;        memory[44149] <=  8'h61;        memory[44150] <=  8'h74;        memory[44151] <=  8'h61;        memory[44152] <=  8'h6e;        memory[44153] <=  8'h61;        memory[44154] <=  8'h62;        memory[44155] <=  8'h61;        memory[44156] <=  8'h63;        memory[44157] <=  8'h61;        memory[44158] <=  8'h74;        memory[44159] <=  8'h61;        memory[44160] <=  8'h62;        memory[44161] <=  8'h61;        memory[44162] <=  8'h72;        memory[44163] <=  8'h63;        memory[44164] <=  8'h61;        memory[44165] <=  8'h68;        memory[44166] <=  8'h64;        memory[44167] <=  8'h75;        memory[44168] <=  8'h63;        memory[44169] <=  8'h74;        memory[44170] <=  8'h61;        memory[44171] <=  8'h64;        memory[44172] <=  8'h61;        memory[44173] <=  8'h61;        memory[44174] <=  8'h63;        memory[44175] <=  8'h61;        memory[44176] <=  8'h72;        memory[44177] <=  8'h63;        memory[44178] <=  8'h74;        memory[44179] <=  8'h72;        memory[44180] <=  8'h63;        memory[44181] <=  8'h61;        memory[44182] <=  8'h74;        memory[44183] <=  8'h72;        memory[44184] <=  8'h63;        memory[44185] <=  8'h61;        memory[44186] <=  8'h74;        memory[44187] <=  8'h63;        memory[44188] <=  8'h62;        memory[44189] <=  8'h61;        memory[44190] <=  8'h74;        memory[44191] <=  8'h62;        memory[44192] <=  8'h72;        memory[44193] <=  8'h63;        memory[44194] <=  8'h61;        memory[44195] <=  8'h74;        memory[44196] <=  8'h72;        memory[44197] <=  8'h6e;        memory[44198] <=  8'h62;        memory[44199] <=  8'h61;        memory[44200] <=  8'h63;        memory[44201] <=  8'h61;        memory[44202] <=  8'h74;        memory[44203] <=  8'h79;        memory[44204] <=  8'h73;        memory[44205] <=  8'h6e;        memory[44206] <=  8'h63;        memory[44207] <=  8'h74;        memory[44208] <=  8'h61;        memory[44209] <=  8'h6e;        memory[44210] <=  8'h62;        memory[44211] <=  8'h61;        memory[44212] <=  8'h63;        memory[44213] <=  8'h72;        memory[44214] <=  8'h6e;        memory[44215] <=  8'h74;        memory[44216] <=  8'h61;        memory[44217] <=  8'h62;        memory[44218] <=  8'h74;        memory[44219] <=  8'h6e;        memory[44220] <=  8'h61;        memory[44221] <=  8'h72;        memory[44222] <=  8'h62;        memory[44223] <=  8'h78;        memory[44224] <=  8'h74;        memory[44225] <=  8'h61;        memory[44226] <=  8'h72;        memory[44227] <=  8'h62;        memory[44228] <=  8'h61;        memory[44229] <=  8'h72;        memory[44230] <=  8'h74;        memory[44231] <=  8'h74;        memory[44232] <=  8'h62;        memory[44233] <=  8'h61;        memory[44234] <=  8'h72;        memory[44235] <=  8'h74;        memory[44236] <=  8'h78;        memory[44237] <=  8'h61;        memory[44238] <=  8'h74;        memory[44239] <=  8'h6b;        memory[44240] <=  8'h73;        memory[44241] <=  8'h68;        memory[44242] <=  8'h63;        memory[44243] <=  8'h66;        memory[44244] <=  8'h69;        memory[44245] <=  8'h77;        memory[44246] <=  8'h68;        memory[44247] <=  8'h61;        memory[44248] <=  8'h74;        memory[44249] <=  8'h61;        memory[44250] <=  8'h6e;        memory[44251] <=  8'h61;        memory[44252] <=  8'h62;        memory[44253] <=  8'h61;        memory[44254] <=  8'h63;        memory[44255] <=  8'h61;        memory[44256] <=  8'h74;        memory[44257] <=  8'h61;        memory[44258] <=  8'h62;        memory[44259] <=  8'h61;        memory[44260] <=  8'h72;        memory[44261] <=  8'h63;        memory[44262] <=  8'h61;        memory[44263] <=  8'h68;        memory[44264] <=  8'h64;        memory[44265] <=  8'h75;        memory[44266] <=  8'h63;        memory[44267] <=  8'h74;        memory[44268] <=  8'h61;        memory[44269] <=  8'h64;        memory[44270] <=  8'h61;        memory[44271] <=  8'h61;        memory[44272] <=  8'h63;        memory[44273] <=  8'h61;        memory[44274] <=  8'h72;        memory[44275] <=  8'h63;        memory[44276] <=  8'h74;        memory[44277] <=  8'h72;        memory[44278] <=  8'h63;        memory[44279] <=  8'h61;        memory[44280] <=  8'h74;        memory[44281] <=  8'h72;        memory[44282] <=  8'h63;        memory[44283] <=  8'h61;        memory[44284] <=  8'h74;        memory[44285] <=  8'h63;        memory[44286] <=  8'h62;        memory[44287] <=  8'h61;        memory[44288] <=  8'h74;        memory[44289] <=  8'h62;        memory[44290] <=  8'h72;        memory[44291] <=  8'h63;        memory[44292] <=  8'h61;        memory[44293] <=  8'h74;        memory[44294] <=  8'h72;        memory[44295] <=  8'h6e;        memory[44296] <=  8'h62;        memory[44297] <=  8'h61;        memory[44298] <=  8'h63;        memory[44299] <=  8'h61;        memory[44300] <=  8'h74;        memory[44301] <=  8'h79;        memory[44302] <=  8'h73;        memory[44303] <=  8'h6e;        memory[44304] <=  8'h63;        memory[44305] <=  8'h74;        memory[44306] <=  8'h61;        memory[44307] <=  8'h6e;        memory[44308] <=  8'h62;        memory[44309] <=  8'h61;        memory[44310] <=  8'h63;        memory[44311] <=  8'h72;        memory[44312] <=  8'h6e;        memory[44313] <=  8'h74;        memory[44314] <=  8'h61;        memory[44315] <=  8'h62;        memory[44316] <=  8'h74;        memory[44317] <=  8'h6e;        memory[44318] <=  8'h61;        memory[44319] <=  8'h72;        memory[44320] <=  8'h62;        memory[44321] <=  8'h78;        memory[44322] <=  8'h74;        memory[44323] <=  8'h61;        memory[44324] <=  8'h72;        memory[44325] <=  8'h64;        memory[44326] <=  8'h66;        memory[44327] <=  8'h73;        memory[44328] <=  8'h67;        memory[44329] <=  8'h76;        memory[44330] <=  8'h68;        memory[44331] <=  8'h62;        memory[44332] <=  8'h6b;        memory[44333] <=  8'h6a;        memory[44334] <=  8'h6e;        memory[44335] <=  8'h6d;        memory[44336] <=  8'h62;        memory[44337] <=  8'h76;        memory[44338] <=  8'h78;        memory[44339] <=  8'h63;        memory[44340] <=  8'h73;        memory[44341] <=  8'h66;        memory[44342] <=  8'h72;        memory[44343] <=  8'h74;        memory[44344] <=  8'h79;        memory[44345] <=  8'h75;        memory[44346] <=  8'h6a;        memory[44347] <=  8'h6e;        memory[44348] <=  8'h62;        memory[44349] <=  8'h76;        memory[44350] <=  8'h63;        memory[44351] <=  8'h64;        memory[44352] <=  8'h74;        memory[44353] <=  8'h79;        memory[44354] <=  8'h75;        memory[44355] <=  8'h69;        memory[44356] <=  8'h6b;        memory[44357] <=  8'h6d;        memory[44358] <=  8'h6e;        memory[44359] <=  8'h62;        memory[44360] <=  8'h76;        memory[44361] <=  8'h63;        memory[44362] <=  8'h78;        memory[44363] <=  8'h73;        memory[44364] <=  8'h64;        memory[44365] <=  8'h72;        memory[44366] <=  8'h74;        memory[44367] <=  8'h79;        memory[44368] <=  8'h75;        memory[44369] <=  8'h69;        memory[44370] <=  8'h6b;        memory[44371] <=  8'h6d;        memory[44372] <=  8'h6e;        memory[44373] <=  8'h62;        memory[44374] <=  8'h76;        memory[44375] <=  8'h63;        memory[44376] <=  8'h73;        memory[44377] <=  8'h77;        memory[44378] <=  8'h33;        memory[44379] <=  8'h34;        memory[44380] <=  8'h35;        memory[44381] <=  8'h36;        memory[44382] <=  8'h37;        memory[44383] <=  8'h38;        memory[44384] <=  8'h69;        memory[44385] <=  8'h6b;        memory[44386] <=  8'h6d;        memory[44387] <=  8'h6e;        memory[44388] <=  8'h62;        memory[44389] <=  8'h76;        memory[44390] <=  8'h63;        memory[44391] <=  8'h64;        memory[44392] <=  8'h65;        memory[44393] <=  8'h72;        memory[44394] <=  8'h36;        memory[44395] <=  8'h37;        memory[44396] <=  8'h38;        memory[44397] <=  8'h69;        memory[44398] <=  8'h6f;        memory[44399] <=  8'h6b;        memory[44400] <=  8'h6a;        memory[44401] <=  8'h6e;        memory[44402] <=  8'h62;        memory[44403] <=  8'h76;        memory[44404] <=  8'h63;        memory[44405] <=  8'h64;        memory[44406] <=  8'h72;        memory[44407] <=  8'h74;        memory[44408] <=  8'h79;        memory[44409] <=  8'h75;        memory[44410] <=  8'h73;        memory[44411] <=  8'h6a;        memory[44412] <=  8'h63;        memory[44413] <=  8'h6e;        memory[44414] <=  8'h62;        memory[44415] <=  8'h64;        memory[44416] <=  8'h66;        memory[44417] <=  8'h73;        memory[44418] <=  8'h74;        memory[44419] <=  8'h79;        memory[44420] <=  8'h75;        memory[44421] <=  8'h61;        memory[44422] <=  8'h69;        memory[44423] <=  8'h6b;        memory[44424] <=  8'h78;        memory[44425] <=  8'h6d;        memory[44426] <=  8'h6e;        memory[44427] <=  8'h73;        memory[44428] <=  8'h6a;        memory[44429] <=  8'h6f;        memory[44430] <=  8'h64;        memory[44431] <=  8'h6c;        memory[44432] <=  8'h63;        memory[44433] <=  8'h78;        memory[44434] <=  8'h62;        memory[44435] <=  8'h61;        memory[44436] <=  8'h72;        memory[44437] <=  8'h74;        memory[44438] <=  8'h78;        memory[44439] <=  8'h61;        memory[44440] <=  8'h74;        memory[44441] <=  8'h6b;        memory[44442] <=  8'h73;        memory[44443] <=  8'h68;        memory[44444] <=  8'h63;        memory[44445] <=  8'h66;        memory[44446] <=  8'h69;        memory[44447] <=  8'h77;        memory[44448] <=  8'h68;        memory[44449] <=  8'h61;        memory[44450] <=  8'h74;        memory[44451] <=  8'h61;        memory[44452] <=  8'h6e;        memory[44453] <=  8'h61;        memory[44454] <=  8'h62;        memory[44455] <=  8'h61;        memory[44456] <=  8'h63;        memory[44457] <=  8'h61;        memory[44458] <=  8'h74;        memory[44459] <=  8'h61;        memory[44460] <=  8'h62;        memory[44461] <=  8'h61;        memory[44462] <=  8'h72;        memory[44463] <=  8'h63;        memory[44464] <=  8'h61;        memory[44465] <=  8'h68;        memory[44466] <=  8'h64;        memory[44467] <=  8'h75;        memory[44468] <=  8'h63;        memory[44469] <=  8'h74;        memory[44470] <=  8'h61;        memory[44471] <=  8'h64;        memory[44472] <=  8'h61;        memory[44473] <=  8'h61;        memory[44474] <=  8'h63;        memory[44475] <=  8'h61;        memory[44476] <=  8'h72;        memory[44477] <=  8'h62;        memory[44478] <=  8'h61;        memory[44479] <=  8'h72;        memory[44480] <=  8'h74;        memory[44481] <=  8'h78;        memory[44482] <=  8'h61;        memory[44483] <=  8'h74;        memory[44484] <=  8'h6b;        memory[44485] <=  8'h73;        memory[44486] <=  8'h68;        memory[44487] <=  8'h63;        memory[44488] <=  8'h66;        memory[44489] <=  8'h69;        memory[44490] <=  8'h77;        memory[44491] <=  8'h68;        memory[44492] <=  8'h61;        memory[44493] <=  8'h74;        memory[44494] <=  8'h61;        memory[44495] <=  8'h6e;        memory[44496] <=  8'h61;        memory[44497] <=  8'h62;        memory[44498] <=  8'h61;        memory[44499] <=  8'h63;        memory[44500] <=  8'h61;        memory[44501] <=  8'h74;        memory[44502] <=  8'h61;        memory[44503] <=  8'h62;        memory[44504] <=  8'h61;        memory[44505] <=  8'h72;        memory[44506] <=  8'h63;        memory[44507] <=  8'h61;        memory[44508] <=  8'h68;        memory[44509] <=  8'h64;        memory[44510] <=  8'h75;        memory[44511] <=  8'h63;        memory[44512] <=  8'h74;        memory[44513] <=  8'h61;        memory[44514] <=  8'h64;        memory[44515] <=  8'h61;        memory[44516] <=  8'h61;        memory[44517] <=  8'h63;        memory[44518] <=  8'h61;        memory[44519] <=  8'h72;        memory[44520] <=  8'h62;        memory[44521] <=  8'h61;        memory[44522] <=  8'h72;        memory[44523] <=  8'h74;        memory[44524] <=  8'h78;        memory[44525] <=  8'h61;        memory[44526] <=  8'h74;        memory[44527] <=  8'h6b;        memory[44528] <=  8'h73;        memory[44529] <=  8'h68;        memory[44530] <=  8'h63;        memory[44531] <=  8'h66;        memory[44532] <=  8'h69;        memory[44533] <=  8'h77;        memory[44534] <=  8'h68;        memory[44535] <=  8'h61;        memory[44536] <=  8'h74;        memory[44537] <=  8'h61;        memory[44538] <=  8'h6e;        memory[44539] <=  8'h61;        memory[44540] <=  8'h62;        memory[44541] <=  8'h61;        memory[44542] <=  8'h63;        memory[44543] <=  8'h61;        memory[44544] <=  8'h74;        memory[44545] <=  8'h61;        memory[44546] <=  8'h62;        memory[44547] <=  8'h61;        memory[44548] <=  8'h72;        memory[44549] <=  8'h63;        memory[44550] <=  8'h61;        memory[44551] <=  8'h68;        memory[44552] <=  8'h64;        memory[44553] <=  8'h75;        memory[44554] <=  8'h63;        memory[44555] <=  8'h74;        memory[44556] <=  8'h61;        memory[44557] <=  8'h64;        memory[44558] <=  8'h61;        memory[44559] <=  8'h61;        memory[44560] <=  8'h63;        memory[44561] <=  8'h61;        memory[44562] <=  8'h72;        memory[44563] <=  8'h62;        memory[44564] <=  8'h61;        memory[44565] <=  8'h72;        memory[44566] <=  8'h74;        memory[44567] <=  8'h78;        memory[44568] <=  8'h61;        memory[44569] <=  8'h74;        memory[44570] <=  8'h6b;        memory[44571] <=  8'h73;        memory[44572] <=  8'h68;        memory[44573] <=  8'h63;        memory[44574] <=  8'h66;        memory[44575] <=  8'h69;        memory[44576] <=  8'h77;        memory[44577] <=  8'h68;        memory[44578] <=  8'h61;        memory[44579] <=  8'h74;        memory[44580] <=  8'h61;        memory[44581] <=  8'h6e;        memory[44582] <=  8'h61;        memory[44583] <=  8'h62;        memory[44584] <=  8'h61;        memory[44585] <=  8'h63;        memory[44586] <=  8'h61;        memory[44587] <=  8'h74;        memory[44588] <=  8'h61;        memory[44589] <=  8'h62;        memory[44590] <=  8'h61;        memory[44591] <=  8'h72;        memory[44592] <=  8'h63;        memory[44593] <=  8'h61;        memory[44594] <=  8'h68;        memory[44595] <=  8'h64;        memory[44596] <=  8'h75;        memory[44597] <=  8'h63;        memory[44598] <=  8'h74;        memory[44599] <=  8'h61;        memory[44600] <=  8'h64;        memory[44601] <=  8'h61;        memory[44602] <=  8'h61;        memory[44603] <=  8'h63;        memory[44604] <=  8'h61;        memory[44605] <=  8'h72;        memory[44606] <=  8'h62;        memory[44607] <=  8'h61;        memory[44608] <=  8'h72;        memory[44609] <=  8'h74;        memory[44610] <=  8'h78;        memory[44611] <=  8'h61;        memory[44612] <=  8'h74;        memory[44613] <=  8'h6b;        memory[44614] <=  8'h73;        memory[44615] <=  8'h68;        memory[44616] <=  8'h63;        memory[44617] <=  8'h66;        memory[44618] <=  8'h69;        memory[44619] <=  8'h77;        memory[44620] <=  8'h68;        memory[44621] <=  8'h61;        memory[44622] <=  8'h74;        memory[44623] <=  8'h61;        memory[44624] <=  8'h6e;        memory[44625] <=  8'h61;        memory[44626] <=  8'h62;        memory[44627] <=  8'h61;        memory[44628] <=  8'h63;        memory[44629] <=  8'h61;        memory[44630] <=  8'h74;        memory[44631] <=  8'h61;        memory[44632] <=  8'h62;        memory[44633] <=  8'h61;        memory[44634] <=  8'h72;        memory[44635] <=  8'h63;        memory[44636] <=  8'h61;        memory[44637] <=  8'h68;        memory[44638] <=  8'h64;        memory[44639] <=  8'h75;        memory[44640] <=  8'h63;        memory[44641] <=  8'h74;        memory[44642] <=  8'h61;        memory[44643] <=  8'h64;        memory[44644] <=  8'h61;        memory[44645] <=  8'h61;        memory[44646] <=  8'h63;        memory[44647] <=  8'h61;        memory[44648] <=  8'h72;        memory[44649] <=  8'h62;        memory[44650] <=  8'h61;        memory[44651] <=  8'h72;        memory[44652] <=  8'h74;        memory[44653] <=  8'h78;        memory[44654] <=  8'h61;        memory[44655] <=  8'h74;        memory[44656] <=  8'h6b;        memory[44657] <=  8'h73;        memory[44658] <=  8'h68;        memory[44659] <=  8'h63;        memory[44660] <=  8'h66;        memory[44661] <=  8'h69;        memory[44662] <=  8'h77;        memory[44663] <=  8'h68;        memory[44664] <=  8'h61;        memory[44665] <=  8'h74;        memory[44666] <=  8'h61;        memory[44667] <=  8'h6e;        memory[44668] <=  8'h61;        memory[44669] <=  8'h62;        memory[44670] <=  8'h61;        memory[44671] <=  8'h63;        memory[44672] <=  8'h61;        memory[44673] <=  8'h74;        memory[44674] <=  8'h61;        memory[44675] <=  8'h62;        memory[44676] <=  8'h61;        memory[44677] <=  8'h72;        memory[44678] <=  8'h63;        memory[44679] <=  8'h61;        memory[44680] <=  8'h68;        memory[44681] <=  8'h64;        memory[44682] <=  8'h75;        memory[44683] <=  8'h63;        memory[44684] <=  8'h74;        memory[44685] <=  8'h61;        memory[44686] <=  8'h64;        memory[44687] <=  8'h61;        memory[44688] <=  8'h61;        memory[44689] <=  8'h63;        memory[44690] <=  8'h61;        memory[44691] <=  8'h72;        memory[44692] <=  8'h62;        memory[44693] <=  8'h61;        memory[44694] <=  8'h72;        memory[44695] <=  8'h74;        memory[44696] <=  8'h78;        memory[44697] <=  8'h61;        memory[44698] <=  8'h74;        memory[44699] <=  8'h6b;        memory[44700] <=  8'h73;        memory[44701] <=  8'h68;        memory[44702] <=  8'h63;        memory[44703] <=  8'h66;        memory[44704] <=  8'h69;        memory[44705] <=  8'h77;        memory[44706] <=  8'h68;        memory[44707] <=  8'h61;        memory[44708] <=  8'h74;        memory[44709] <=  8'h61;        memory[44710] <=  8'h6e;        memory[44711] <=  8'h61;        memory[44712] <=  8'h62;        memory[44713] <=  8'h61;        memory[44714] <=  8'h63;        memory[44715] <=  8'h61;        memory[44716] <=  8'h74;        memory[44717] <=  8'h61;        memory[44718] <=  8'h62;        memory[44719] <=  8'h61;        memory[44720] <=  8'h72;        memory[44721] <=  8'h63;        memory[44722] <=  8'h61;        memory[44723] <=  8'h68;        memory[44724] <=  8'h64;        memory[44725] <=  8'h75;        memory[44726] <=  8'h63;        memory[44727] <=  8'h74;        memory[44728] <=  8'h61;        memory[44729] <=  8'h64;        memory[44730] <=  8'h61;        memory[44731] <=  8'h61;        memory[44732] <=  8'h63;        memory[44733] <=  8'h61;        memory[44734] <=  8'h72;        memory[44735] <=  8'h62;        memory[44736] <=  8'h61;        memory[44737] <=  8'h72;        memory[44738] <=  8'h74;        memory[44739] <=  8'h78;        memory[44740] <=  8'h61;        memory[44741] <=  8'h74;        memory[44742] <=  8'h6b;        memory[44743] <=  8'h73;        memory[44744] <=  8'h68;        memory[44745] <=  8'h63;        memory[44746] <=  8'h66;        memory[44747] <=  8'h69;        memory[44748] <=  8'h77;        memory[44749] <=  8'h68;        memory[44750] <=  8'h61;        memory[44751] <=  8'h74;        memory[44752] <=  8'h61;        memory[44753] <=  8'h6e;        memory[44754] <=  8'h61;        memory[44755] <=  8'h62;        memory[44756] <=  8'h61;        memory[44757] <=  8'h63;        memory[44758] <=  8'h61;        memory[44759] <=  8'h74;        memory[44760] <=  8'h61;        memory[44761] <=  8'h62;        memory[44762] <=  8'h61;        memory[44763] <=  8'h72;        memory[44764] <=  8'h63;        memory[44765] <=  8'h61;        memory[44766] <=  8'h68;        memory[44767] <=  8'h64;        memory[44768] <=  8'h75;        memory[44769] <=  8'h63;        memory[44770] <=  8'h74;        memory[44771] <=  8'h61;        memory[44772] <=  8'h64;        memory[44773] <=  8'h61;        memory[44774] <=  8'h61;        memory[44775] <=  8'h63;        memory[44776] <=  8'h61;        memory[44777] <=  8'h72;        memory[44778] <=  8'h62;        memory[44779] <=  8'h61;        memory[44780] <=  8'h72;        memory[44781] <=  8'h74;        memory[44782] <=  8'h78;        memory[44783] <=  8'h61;        memory[44784] <=  8'h74;        memory[44785] <=  8'h6b;        memory[44786] <=  8'h73;        memory[44787] <=  8'h68;        memory[44788] <=  8'h63;        memory[44789] <=  8'h66;        memory[44790] <=  8'h69;        memory[44791] <=  8'h77;        memory[44792] <=  8'h68;        memory[44793] <=  8'h61;        memory[44794] <=  8'h74;        memory[44795] <=  8'h61;        memory[44796] <=  8'h6e;        memory[44797] <=  8'h61;        memory[44798] <=  8'h62;        memory[44799] <=  8'h61;        memory[44800] <=  8'h63;        memory[44801] <=  8'h61;        memory[44802] <=  8'h74;        memory[44803] <=  8'h61;        memory[44804] <=  8'h62;        memory[44805] <=  8'h61;        memory[44806] <=  8'h72;        memory[44807] <=  8'h63;        memory[44808] <=  8'h61;        memory[44809] <=  8'h68;        memory[44810] <=  8'h64;        memory[44811] <=  8'h75;        memory[44812] <=  8'h63;        memory[44813] <=  8'h74;        memory[44814] <=  8'h61;        memory[44815] <=  8'h64;        memory[44816] <=  8'h61;        memory[44817] <=  8'h61;        memory[44818] <=  8'h63;        memory[44819] <=  8'h61;        memory[44820] <=  8'h72;        memory[44821] <=  8'h62;        memory[44822] <=  8'h61;        memory[44823] <=  8'h72;        memory[44824] <=  8'h74;        memory[44825] <=  8'h74;        memory[44826] <=  8'h62;        memory[44827] <=  8'h61;        memory[44828] <=  8'h72;        memory[44829] <=  8'h74;        memory[44830] <=  8'h78;        memory[44831] <=  8'h61;        memory[44832] <=  8'h74;        memory[44833] <=  8'h6b;        memory[44834] <=  8'h73;        memory[44835] <=  8'h68;        memory[44836] <=  8'h63;        memory[44837] <=  8'h66;        memory[44838] <=  8'h69;        memory[44839] <=  8'h77;        memory[44840] <=  8'h68;        memory[44841] <=  8'h61;        memory[44842] <=  8'h74;        memory[44843] <=  8'h61;        memory[44844] <=  8'h6e;        memory[44845] <=  8'h61;        memory[44846] <=  8'h62;        memory[44847] <=  8'h61;        memory[44848] <=  8'h63;        memory[44849] <=  8'h61;        memory[44850] <=  8'h74;        memory[44851] <=  8'h61;        memory[44852] <=  8'h62;        memory[44853] <=  8'h61;        memory[44854] <=  8'h72;        memory[44855] <=  8'h63;        memory[44856] <=  8'h61;        memory[44857] <=  8'h68;        memory[44858] <=  8'h64;        memory[44859] <=  8'h75;        memory[44860] <=  8'h63;        memory[44861] <=  8'h74;        memory[44862] <=  8'h61;        memory[44863] <=  8'h64;        memory[44864] <=  8'h61;        memory[44865] <=  8'h61;        memory[44866] <=  8'h63;        memory[44867] <=  8'h61;        memory[44868] <=  8'h72;        memory[44869] <=  8'h63;        memory[44870] <=  8'h74;        memory[44871] <=  8'h72;        memory[44872] <=  8'h63;        memory[44873] <=  8'h61;        memory[44874] <=  8'h74;        memory[44875] <=  8'h72;        memory[44876] <=  8'h63;        memory[44877] <=  8'h61;        memory[44878] <=  8'h74;        memory[44879] <=  8'h63;        memory[44880] <=  8'h62;        memory[44881] <=  8'h61;        memory[44882] <=  8'h74;        memory[44883] <=  8'h62;        memory[44884] <=  8'h72;        memory[44885] <=  8'h63;        memory[44886] <=  8'h61;        memory[44887] <=  8'h72;        memory[44888] <=  8'h62;        memory[44889] <=  8'h78;        memory[44890] <=  8'h74;        memory[44891] <=  8'h61;        memory[44892] <=  8'h72;        memory[44893] <=  8'h64;        memory[44894] <=  8'h66;        memory[44895] <=  8'h73;        memory[44896] <=  8'h67;        memory[44897] <=  8'h76;        memory[44898] <=  8'h68;        memory[44899] <=  8'h62;        memory[44900] <=  8'h6b;        memory[44901] <=  8'h6a;        memory[44902] <=  8'h6e;        memory[44903] <=  8'h6d;        memory[44904] <=  8'h62;        memory[44905] <=  8'h76;        memory[44906] <=  8'h78;        memory[44907] <=  8'h63;        memory[44908] <=  8'h73;        memory[44909] <=  8'h66;        memory[44910] <=  8'h72;        memory[44911] <=  8'h74;        memory[44912] <=  8'h79;        memory[44913] <=  8'h75;        memory[44914] <=  8'h6a;        memory[44915] <=  8'h6e;        memory[44916] <=  8'h62;        memory[44917] <=  8'h76;        memory[44918] <=  8'h63;        memory[44919] <=  8'h64;        memory[44920] <=  8'h74;        memory[44921] <=  8'h79;        memory[44922] <=  8'h75;        memory[44923] <=  8'h69;        memory[44924] <=  8'h6b;        memory[44925] <=  8'h6d;        memory[44926] <=  8'h6e;        memory[44927] <=  8'h62;        memory[44928] <=  8'h76;        memory[44929] <=  8'h63;        memory[44930] <=  8'h78;        memory[44931] <=  8'h73;        memory[44932] <=  8'h64;        memory[44933] <=  8'h72;        memory[44934] <=  8'h74;        memory[44935] <=  8'h79;        memory[44936] <=  8'h75;        memory[44937] <=  8'h69;        memory[44938] <=  8'h6b;        memory[44939] <=  8'h6d;        memory[44940] <=  8'h6e;        memory[44941] <=  8'h62;        memory[44942] <=  8'h76;        memory[44943] <=  8'h63;        memory[44944] <=  8'h73;        memory[44945] <=  8'h77;        memory[44946] <=  8'h33;        memory[44947] <=  8'h34;        memory[44948] <=  8'h35;        memory[44949] <=  8'h36;        memory[44950] <=  8'h37;        memory[44951] <=  8'h38;        memory[44952] <=  8'h69;        memory[44953] <=  8'h6b;        memory[44954] <=  8'h6d;        memory[44955] <=  8'h6e;        memory[44956] <=  8'h62;        memory[44957] <=  8'h76;        memory[44958] <=  8'h63;        memory[44959] <=  8'h64;        memory[44960] <=  8'h65;        memory[44961] <=  8'h72;        memory[44962] <=  8'h36;        memory[44963] <=  8'h37;        memory[44964] <=  8'h38;        memory[44965] <=  8'h69;        memory[44966] <=  8'h6f;        memory[44967] <=  8'h6b;        memory[44968] <=  8'h6a;        memory[44969] <=  8'h6e;        memory[44970] <=  8'h62;        memory[44971] <=  8'h76;        memory[44972] <=  8'h63;        memory[44973] <=  8'h64;        memory[44974] <=  8'h72;        memory[44975] <=  8'h74;        memory[44976] <=  8'h79;        memory[44977] <=  8'h75;        memory[44978] <=  8'h73;        memory[44979] <=  8'h6a;        memory[44980] <=  8'h63;        memory[44981] <=  8'h6e;        memory[44982] <=  8'h62;        memory[44983] <=  8'h64;        memory[44984] <=  8'h66;        memory[44985] <=  8'h73;        memory[44986] <=  8'h74;        memory[44987] <=  8'h79;        memory[44988] <=  8'h75;        memory[44989] <=  8'h61;        memory[44990] <=  8'h69;        memory[44991] <=  8'h6b;        memory[44992] <=  8'h78;        memory[44993] <=  8'h6d;        memory[44994] <=  8'h6e;        memory[44995] <=  8'h73;        memory[44996] <=  8'h6a;        memory[44997] <=  8'h6f;        memory[44998] <=  8'h64;        memory[44999] <=  8'h6c;        memory[45000] <=  8'h63;        memory[45001] <=  8'h78;        memory[45002] <=  8'h2c;        memory[45003] <=  8'h6d;        memory[45004] <=  8'h73;        memory[45005] <=  8'h6b;        memory[45006] <=  8'h64;        memory[45007] <=  8'h6c;        memory[45008] <=  8'h70;        memory[45009] <=  8'h5b;        memory[45010] <=  8'h3b;        memory[45011] <=  8'h73;        memory[45012] <=  8'h6c;        memory[45013] <=  8'h64;        memory[45014] <=  8'h70;        memory[45015] <=  8'h76;        memory[45016] <=  8'h63;        memory[45017] <=  8'h5b;        memory[45018] <=  8'h78;        memory[45019] <=  8'h76;        memory[45020] <=  8'h63;        memory[45021] <=  8'h5b;        memory[45022] <=  8'h78;        memory[45023] <=  8'h70;        memory[45024] <=  8'h6f;        memory[45025] <=  8'h20;        memory[45026] <=  8'h62;        memory[45027] <=  8'h61;        memory[45028] <=  8'h72;        memory[45029] <=  8'h74;        memory[45030] <=  8'h74;        memory[45031] <=  8'h62;        memory[45032] <=  8'h61;        memory[45033] <=  8'h72;        memory[45034] <=  8'h74;        memory[45035] <=  8'h78;        memory[45036] <=  8'h61;        memory[45037] <=  8'h74;        memory[45038] <=  8'h6b;        memory[45039] <=  8'h73;        memory[45040] <=  8'h68;        memory[45041] <=  8'h63;        memory[45042] <=  8'h66;        memory[45043] <=  8'h69;        memory[45044] <=  8'h77;        memory[45045] <=  8'h68;        memory[45046] <=  8'h61;        memory[45047] <=  8'h69;        memory[45048] <=  8'h6a;        memory[45049] <=  8'h78;        memory[45050] <=  8'h5d;        memory[45051] <=  8'h65;        memory[45052] <=  8'h6b;        memory[45053] <=  8'h6f;        memory[45054] <=  8'h39;        memory[45055] <=  8'h64;        memory[45056] <=  8'h75;        memory[45057] <=  8'h38;        memory[45058] <=  8'h79;        memory[45059] <=  8'h20;        memory[45060] <=  8'h37;        memory[45061] <=  8'h63;        memory[45062] <=  8'h67;        memory[45063] <=  8'h78;        memory[45064] <=  8'h63;        memory[45065] <=  8'h75;        memory[45066] <=  8'h68;        memory[45067] <=  8'h69;        memory[45068] <=  8'h6a;        memory[45069] <=  8'h77;        memory[45070] <=  8'h69;        memory[45071] <=  8'h64;        memory[45072] <=  8'h66;        memory[45073] <=  8'h68;        memory[45074] <=  8'h75;        memory[45075] <=  8'h76;        memory[45076] <=  8'h64;        memory[45077] <=  8'h62;        memory[45078] <=  8'h66;        memory[45079] <=  8'h6a;        memory[45080] <=  8'h6e;        memory[45081] <=  8'h6b;        memory[45082] <=  8'h6a;        memory[45083] <=  8'h65;        memory[45084] <=  8'h38;        memory[45085] <=  8'h66;        memory[45086] <=  8'h37;        memory[45087] <=  8'h67;        memory[45088] <=  8'h79;        memory[45089] <=  8'h76;        memory[45090] <=  8'h63;        memory[45091] <=  8'h68;        memory[45092] <=  8'h69;        memory[45093] <=  8'h6a;        memory[45094] <=  8'h33;        memory[45095] <=  8'h65;        memory[45096] <=  8'h67;        memory[45097] <=  8'h79;        memory[45098] <=  8'h72;        memory[45099] <=  8'h64;        memory[45100] <=  8'h62;        memory[45101] <=  8'h6e;        memory[45102] <=  8'h63;        memory[45103] <=  8'h7a;        memory[45104] <=  8'h6a;        memory[45105] <=  8'h6f;        memory[45106] <=  8'h66;        memory[45107] <=  8'h78;        memory[45108] <=  8'h6a;        memory[45109] <=  8'h69;        memory[45110] <=  8'h63;        memory[45111] <=  8'h68;        memory[45112] <=  8'h62;        memory[45113] <=  8'h6e;        memory[45114] <=  8'h6d;        memory[45115] <=  8'h63;        memory[45116] <=  8'h73;        memory[45117] <=  8'h6c;        memory[45118] <=  8'h6b;        memory[45119] <=  8'h6a;        memory[45120] <=  8'h69;        memory[45121] <=  8'h68;        memory[45122] <=  8'h76;        memory[45123] <=  8'h75;        memory[45124] <=  8'h69;        memory[45125] <=  8'h64;        memory[45126] <=  8'h68;        memory[45127] <=  8'h75;        memory[45128] <=  8'h67;        memory[45129] <=  8'h79;        memory[45130] <=  8'h62;        memory[45131] <=  8'h68;        memory[45132] <=  8'h65;        memory[45133] <=  8'h6a;        memory[45134] <=  8'h72;        memory[45135] <=  8'h6b;        memory[45136] <=  8'h6a;        memory[45137] <=  8'h6f;        memory[45138] <=  8'h64;        memory[45139] <=  8'h67;        memory[45140] <=  8'h69;        memory[45141] <=  8'h75;        memory[45142] <=  8'h69;        memory[45143] <=  8'h67;        memory[45144] <=  8'h76;        memory[45145] <=  8'h79;        memory[45146] <=  8'h75;        memory[45147] <=  8'h67;        memory[45148] <=  8'h78;        memory[45149] <=  8'h68;        memory[45150] <=  8'h63;        memory[45151] <=  8'h20;        memory[45152] <=  8'h20;        memory[45153] <=  8'h20;        memory[45154] <=  8'h78;        memory[45155] <=  8'h76;        memory[45156] <=  8'h20;        memory[45157] <=  8'h63;        memory[45158] <=  8'h78;        memory[45159] <=  8'h67;        memory[45160] <=  8'h79;        memory[45161] <=  8'h63;        memory[45162] <=  8'h75;        memory[45163] <=  8'h68;        memory[45164] <=  8'h6a;        memory[45165] <=  8'h6b;        memory[45166] <=  8'h61;        memory[45167] <=  8'h6c;        memory[45168] <=  8'h78;        memory[45169] <=  8'h76;        memory[45170] <=  8'h70;        memory[45171] <=  8'h6f;        memory[45172] <=  8'h69;        memory[45173] <=  8'h6a;        memory[45174] <=  8'h69;        memory[45175] <=  8'h68;        memory[45176] <=  8'h6a;        memory[45177] <=  8'h62;        memory[45178] <=  8'h77;        memory[45179] <=  8'h65;        memory[45180] <=  8'h6e;        memory[45181] <=  8'h61;        memory[45182] <=  8'h66;        memory[45183] <=  8'h6d;        memory[45184] <=  8'h64;        memory[45185] <=  8'h6b;        memory[45186] <=  8'h6d;        memory[45187] <=  8'h76;        memory[45188] <=  8'h6c;        memory[45189] <=  8'h63;        memory[45190] <=  8'h6f;        memory[45191] <=  8'h64;        memory[45192] <=  8'h69;        memory[45193] <=  8'h75;        memory[45194] <=  8'h68;        memory[45195] <=  8'h73;        memory[45196] <=  8'h66;        memory[45197] <=  8'h65;        memory[45198] <=  8'h62;        memory[45199] <=  8'h6e;        memory[45200] <=  8'h64;        memory[45201] <=  8'h73;        memory[45202] <=  8'h63;        memory[45203] <=  8'h6b;        memory[45204] <=  8'h20;        memory[45205] <=  8'h78;        memory[45206] <=  8'h6a;        memory[45207] <=  8'h78;        memory[45208] <=  8'h63;        memory[45209] <=  8'h73;        memory[45210] <=  8'h64;        memory[45211] <=  8'h66;        memory[45212] <=  8'h6b;        memory[45213] <=  8'h64;        memory[45214] <=  8'h6e;        memory[45215] <=  8'h6d;        memory[45216] <=  8'h64;        memory[45217] <=  8'h73;        memory[45218] <=  8'h63;        memory[45219] <=  8'h6b;        memory[45220] <=  8'h78;        memory[45221] <=  8'h6c;        memory[45222] <=  8'h6f;        memory[45223] <=  8'h66;        memory[45224] <=  8'h6a;        memory[45225] <=  8'h69;        memory[45226] <=  8'h61;        memory[45227] <=  8'h62;        memory[45228] <=  8'h6e;        memory[45229] <=  8'h20;        memory[45230] <=  8'h78;        memory[45231] <=  8'h6b;        memory[45232] <=  8'h6d;        memory[45233] <=  8'h20;        memory[45234] <=  8'h6f;        memory[45235] <=  8'h63;        memory[45236] <=  8'h76;        memory[45237] <=  8'h73;        memory[45238] <=  8'h64;        memory[45239] <=  8'h69;        memory[45240] <=  8'h66;        memory[45241] <=  8'h68;        memory[45242] <=  8'h65;        memory[45243] <=  8'h71;        memory[45244] <=  8'h6a;        memory[45245] <=  8'h77;        memory[45246] <=  8'h62;        memory[45247] <=  8'h65;        memory[45248] <=  8'h6e;        memory[45249] <=  8'h20;        memory[45250] <=  8'h6d;        memory[45251] <=  8'h64;        memory[45252] <=  8'h73;        memory[45253] <=  8'h6c;        memory[45254] <=  8'h76;        memory[45255] <=  8'h6b;        memory[45256] <=  8'h63;        memory[45257] <=  8'h78;        memory[45258] <=  8'h20;        memory[45259] <=  8'h6f;        memory[45260] <=  8'h78;        memory[45261] <=  8'h69;        memory[45262] <=  8'h63;        memory[45263] <=  8'h6a;        memory[45264] <=  8'h76;        memory[45265] <=  8'h64;        memory[45266] <=  8'h66;        memory[45267] <=  8'h65;        memory[45268] <=  8'h71;        memory[45269] <=  8'h6e;        memory[45270] <=  8'h20;        memory[45271] <=  8'h64;        memory[45272] <=  8'h6d;        memory[45273] <=  8'h73;        memory[45274] <=  8'h6c;        memory[45275] <=  8'h63;        memory[45276] <=  8'h78;        memory[45277] <=  8'h6b;        memory[45278] <=  8'h20;        memory[45279] <=  8'h6f;        memory[45280] <=  8'h78;        memory[45281] <=  8'h63;        memory[45282] <=  8'h76;        memory[45283] <=  8'h6a;        memory[45284] <=  8'h64;        memory[45285] <=  8'h62;        memory[45286] <=  8'h71;        memory[45287] <=  8'h77;        memory[45288] <=  8'h65;        memory[45289] <=  8'h6e;        memory[45290] <=  8'h6d;        memory[45291] <=  8'h64;        memory[45292] <=  8'h6c;        memory[45293] <=  8'h73;        memory[45294] <=  8'h2c;        memory[45295] <=  8'h76;        memory[45296] <=  8'h63;        memory[45297] <=  8'h78;        memory[45298] <=  8'h20;        memory[45299] <=  8'h63;        memory[45300] <=  8'h6f;        memory[45301] <=  8'h69;        memory[45302] <=  8'h76;        memory[45303] <=  8'h68;        memory[45304] <=  8'h73;        memory[45305] <=  8'h64;        memory[45306] <=  8'h62;        memory[45307] <=  8'h71;        memory[45308] <=  8'h77;        memory[45309] <=  8'h65;        memory[45310] <=  8'h6e;        memory[45311] <=  8'h64;        memory[45312] <=  8'h6b;        memory[45313] <=  8'h73;        memory[45314] <=  8'h76;        memory[45315] <=  8'h6f;        memory[45316] <=  8'h63;        memory[45317] <=  8'h20;        memory[45318] <=  8'h76;        memory[45319] <=  8'h69;        memory[45320] <=  8'h75;        memory[45321] <=  8'h69;        memory[45322] <=  8'h68;        memory[45323] <=  8'h63;        memory[45324] <=  8'h78;        memory[45325] <=  8'h69;        memory[45326] <=  8'h6f;        memory[45327] <=  8'h76;        memory[45328] <=  8'h73;        memory[45329] <=  8'h64;        memory[45330] <=  8'h61;        memory[45331] <=  8'h64;        memory[45332] <=  8'h6e;        memory[45333] <=  8'h77;        memory[45334] <=  8'h71;        memory[45335] <=  8'h6b;        memory[45336] <=  8'h6c;        memory[45337] <=  8'h73;        memory[45338] <=  8'h76;        memory[45339] <=  8'h6e;        memory[45340] <=  8'h62;        memory[45341] <=  8'h20;        memory[45342] <=  8'h64;        memory[45343] <=  8'h66;        memory[45344] <=  8'h6a;        memory[45345] <=  8'h6b;        memory[45346] <=  8'h71;        memory[45347] <=  8'h64;        memory[45348] <=  8'h77;        memory[45349] <=  8'h65;        memory[45350] <=  8'h6e;        memory[45351] <=  8'h62;        memory[45352] <=  8'h20;        memory[45353] <=  8'h64;        memory[45354] <=  8'h73;        memory[45355] <=  8'h76;        memory[45356] <=  8'h68;        memory[45357] <=  8'h64;        memory[45358] <=  8'h61;        memory[45359] <=  8'h71;        memory[45360] <=  8'h77;        memory[45361] <=  8'h6a;        memory[45362] <=  8'h65;        memory[45363] <=  8'h6e;        memory[45364] <=  8'h64;        memory[45365] <=  8'h20;        memory[45366] <=  8'h61;        memory[45367] <=  8'h63;        memory[45368] <=  8'h62;        memory[45369] <=  8'h68;        memory[45370] <=  8'h64;        memory[45371] <=  8'h61;        memory[45372] <=  8'h77;        memory[45373] <=  8'h71;        memory[45374] <=  8'h6e;        memory[45375] <=  8'h20;        memory[45376] <=  8'h62;        memory[45377] <=  8'h73;        memory[45378] <=  8'h76;        memory[45379] <=  8'h61;        memory[45380] <=  8'h67;        memory[45381] <=  8'h76;        memory[45382] <=  8'h68;        memory[45383] <=  8'h67;        memory[45384] <=  8'h61;        memory[45385] <=  8'h73;        memory[45386] <=  8'h6a;        memory[45387] <=  8'h6b;        memory[45388] <=  8'h63;        memory[45389] <=  8'h78;        memory[45390] <=  8'h76;        memory[45391] <=  8'h6e;        memory[45392] <=  8'h73;        memory[45393] <=  8'h64;        memory[45394] <=  8'h20;        memory[45395] <=  8'h66;        memory[45396] <=  8'h62;        memory[45397] <=  8'h64;        memory[45398] <=  8'h61;        memory[45399] <=  8'h73;        memory[45400] <=  8'h76;        memory[45401] <=  8'h67;        memory[45402] <=  8'h63;        memory[45403] <=  8'h79;        memory[45404] <=  8'h7a;        memory[45405] <=  8'h78;        memory[45406] <=  8'h79;        memory[45407] <=  8'h75;        memory[45408] <=  8'h20;        memory[45409] <=  8'h69;        memory[45410] <=  8'h6a;        memory[45411] <=  8'h64;        memory[45412] <=  8'h66;        memory[45413] <=  8'h6b;        memory[45414] <=  8'h61;        memory[45415] <=  8'h64;        memory[45416] <=  8'h63;        memory[45417] <=  8'h78;        memory[45418] <=  8'h68;        memory[45419] <=  8'h20;        memory[45420] <=  8'h67;        memory[45421] <=  8'h61;        memory[45422] <=  8'h68;        memory[45423] <=  8'h75;        memory[45424] <=  8'h64;        memory[45425] <=  8'h73;        memory[45426] <=  8'h69;        memory[45427] <=  8'h6a;        memory[45428] <=  8'h61;        memory[45429] <=  8'h6b;        memory[45430] <=  8'h63;        memory[45431] <=  8'h62;        memory[45432] <=  8'h61;        memory[45433] <=  8'h72;        memory[45434] <=  8'h73;        memory[45435] <=  8'h68;        memory[45436] <=  8'h64;        memory[45437] <=  8'h66;        memory[45438] <=  8'h67;        memory[45439] <=  8'h73;        memory[45440] <=  8'h68;        memory[45441] <=  8'h64;        memory[45442] <=  8'h66;        memory[45443] <=  8'h68;        memory[45444] <=  8'h64;        memory[45445] <=  8'h6a;        memory[45446] <=  8'h68;        memory[45447] <=  8'h62;        memory[45448] <=  8'h67;        memory[45449] <=  8'h63;        memory[45450] <=  8'h61;        memory[45451] <=  8'h66;        memory[45452] <=  8'h73;        memory[45453] <=  8'h79;        memory[45454] <=  8'h67;        memory[45455] <=  8'h6b;        memory[45456] <=  8'h75;        memory[45457] <=  8'h64;        memory[45458] <=  8'h68;        memory[45459] <=  8'h62;        memory[45460] <=  8'h77;        memory[45461] <=  8'h76;        memory[45462] <=  8'h67;        memory[45463] <=  8'h61;        memory[45464] <=  8'h66;        memory[45465] <=  8'h64;        memory[45466] <=  8'h74;        memory[45467] <=  8'h75;        memory[45468] <=  8'h66;        memory[45469] <=  8'h79;        memory[45470] <=  8'h67;        memory[45471] <=  8'h69;        memory[45472] <=  8'h75;        memory[45473] <=  8'h68;        memory[45474] <=  8'h6c;        memory[45475] <=  8'h6a;        memory[45476] <=  8'h62;        memory[45477] <=  8'h6b;        memory[45478] <=  8'h68;        memory[45479] <=  8'h76;        memory[45480] <=  8'h67;        memory[45481] <=  8'h63;        memory[45482] <=  8'h66;        memory[45483] <=  8'h78;        memory[45484] <=  8'h64;        memory[45485] <=  8'h74;        memory[45486] <=  8'h75;        memory[45487] <=  8'h79;        memory[45488] <=  8'h69;        memory[45489] <=  8'h75;        memory[45490] <=  8'h68;        memory[45491] <=  8'h6c;        memory[45492] <=  8'h6a;        memory[45493] <=  8'h6b;        memory[45494] <=  8'h67;        memory[45495] <=  8'h6a;        memory[45496] <=  8'h63;        memory[45497] <=  8'h66;        memory[45498] <=  8'h68;        memory[45499] <=  8'h64;        memory[45500] <=  8'h67;        memory[45501] <=  8'h72;        memory[45502] <=  8'h79;        memory[45503] <=  8'h74;        memory[45504] <=  8'h66;        memory[45505] <=  8'h75;        memory[45506] <=  8'h79;        memory[45507] <=  8'h69;        memory[45508] <=  8'h68;        memory[45509] <=  8'h6c;        memory[45510] <=  8'h62;        memory[45511] <=  8'h6d;        memory[45512] <=  8'h76;        memory[45513] <=  8'h6e;        memory[45514] <=  8'h63;        memory[45515] <=  8'h66;        memory[45516] <=  8'h68;        memory[45517] <=  8'h64;        memory[45518] <=  8'h74;        memory[45519] <=  8'h75;        memory[45520] <=  8'h67;        memory[45521] <=  8'h79;        memory[45522] <=  8'h69;        memory[45523] <=  8'h68;        memory[45524] <=  8'h75;        memory[45525] <=  8'h6a;        memory[45526] <=  8'h6c;        memory[45527] <=  8'h62;        memory[45528] <=  8'h6d;        memory[45529] <=  8'h76;        memory[45530] <=  8'h6e;        memory[45531] <=  8'h63;        memory[45532] <=  8'h66;        memory[45533] <=  8'h68;        memory[45534] <=  8'h67;        memory[45535] <=  8'h79;        memory[45536] <=  8'h68;        memory[45537] <=  8'h75;        memory[45538] <=  8'h6a;        memory[45539] <=  8'h6e;        memory[45540] <=  8'h2c;        memory[45541] <=  8'h62;        memory[45542] <=  8'h6e;        memory[45543] <=  8'h6d;        memory[45544] <=  8'h76;        memory[45545] <=  8'h6e;        memory[45546] <=  8'h63;        memory[45547] <=  8'h66;        memory[45548] <=  8'h68;        memory[45549] <=  8'h74;        memory[45550] <=  8'h79;        memory[45551] <=  8'h69;        memory[45552] <=  8'h75;        memory[45553] <=  8'h6c;        memory[45554] <=  8'h6a;        memory[45555] <=  8'h62;        memory[45556] <=  8'h6d;        memory[45557] <=  8'h76;        memory[45558] <=  8'h6e;        memory[45559] <=  8'h63;        memory[45560] <=  8'h66;        memory[45561] <=  8'h74;        memory[45562] <=  8'h75;        memory[45563] <=  8'h79;        memory[45564] <=  8'h69;        memory[45565] <=  8'h68;        memory[45566] <=  8'h6b;        memory[45567] <=  8'h62;        memory[45568] <=  8'h76;        memory[45569] <=  8'h63;        memory[45570] <=  8'h66;        memory[45571] <=  8'h67;        memory[45572] <=  8'h74;        memory[45573] <=  8'h75;        memory[45574] <=  8'h79;        memory[45575] <=  8'h69;        memory[45576] <=  8'h75;        memory[45577] <=  8'h68;        memory[45578] <=  8'h6a;        memory[45579] <=  8'h6b;        memory[45580] <=  8'h62;        memory[45581] <=  8'h76;        memory[45582] <=  8'h63;        memory[45583] <=  8'h66;        memory[45584] <=  8'h74;        memory[45585] <=  8'h75;        memory[45586] <=  8'h79;        memory[45587] <=  8'h69;        memory[45588] <=  8'h75;        memory[45589] <=  8'h6a;        memory[45590] <=  8'h6b;        memory[45591] <=  8'h6e;        memory[45592] <=  8'h62;        memory[45593] <=  8'h76;        memory[45594] <=  8'h67;        memory[45595] <=  8'h66;        memory[45596] <=  8'h74;        memory[45597] <=  8'h79;        memory[45598] <=  8'h75;        memory[45599] <=  8'h75;        memory[45600] <=  8'h69;        memory[45601] <=  8'h6a;        memory[45602] <=  8'h6b;        memory[45603] <=  8'h68;        memory[45604] <=  8'h62;        memory[45605] <=  8'h6a;        memory[45606] <=  8'h67;        memory[45607] <=  8'h68;        memory[45608] <=  8'h66;        memory[45609] <=  8'h79;        memory[45610] <=  8'h74;        memory[45611] <=  8'h79;        memory[45612] <=  8'h69;        memory[45613] <=  8'h75;        memory[45614] <=  8'h64;        memory[45615] <=  8'h6a;        memory[45616] <=  8'h6b;        memory[45617] <=  8'h68;        memory[45618] <=  8'h63;        memory[45619] <=  8'h7a;        memory[45620] <=  8'h67;        memory[45621] <=  8'h68;        memory[45622] <=  8'h74;        memory[45623] <=  8'h75;        memory[45624] <=  8'h79;        memory[45625] <=  8'h69;        memory[45626] <=  8'h61;        memory[45627] <=  8'h73;        memory[45628] <=  8'h75;        memory[45629] <=  8'h6a;        memory[45630] <=  8'h6b;        memory[45631] <=  8'h62;        memory[45632] <=  8'h6e;        memory[45633] <=  8'h61;        memory[45634] <=  8'h76;        memory[45635] <=  8'h63;        memory[45636] <=  8'h66;        memory[45637] <=  8'h68;        memory[45638] <=  8'h75;        memory[45639] <=  8'h61;        memory[45640] <=  8'h73;        memory[45641] <=  8'h79;        memory[45642] <=  8'h64;        memory[45643] <=  8'h75;        memory[45644] <=  8'h69;        memory[45645] <=  8'h6a;        memory[45646] <=  8'h61;        memory[45647] <=  8'h6b;        memory[45648] <=  8'h62;        memory[45649] <=  8'h63;        memory[45650] <=  8'h78;        memory[45651] <=  8'h68;        memory[45652] <=  8'h67;        memory[45653] <=  8'h79;        memory[45654] <=  8'h75;        memory[45655] <=  8'h7a;        memory[45656] <=  8'h63;        memory[45657] <=  8'h61;        memory[45658] <=  8'h73;        memory[45659] <=  8'h69;        memory[45660] <=  8'h75;        memory[45661] <=  8'h6f;        memory[45662] <=  8'h69;        memory[45663] <=  8'h6a;        memory[45664] <=  8'h61;        memory[45665] <=  8'h6c;        memory[45666] <=  8'h63;        memory[45667] <=  8'h78;        memory[45668] <=  8'h62;        memory[45669] <=  8'h63;        memory[45670] <=  8'h20;        memory[45671] <=  8'h6e;        memory[45672] <=  8'h76;        memory[45673] <=  8'h63;        memory[45674] <=  8'h61;        memory[45675] <=  8'h64;        memory[45676] <=  8'h73;        memory[45677] <=  8'h67;        memory[45678] <=  8'h79;        memory[45679] <=  8'h68;        memory[45680] <=  8'h75;        memory[45681] <=  8'h61;        memory[45682] <=  8'h6a;        memory[45683] <=  8'h6b;        memory[45684] <=  8'h78;        memory[45685] <=  8'h62;        memory[45686] <=  8'h20;        memory[45687] <=  8'h6e;        memory[45688] <=  8'h76;        memory[45689] <=  8'h63;        memory[45690] <=  8'h61;        memory[45691] <=  8'h73;        memory[45692] <=  8'h67;        memory[45693] <=  8'h68;        memory[45694] <=  8'h75;        memory[45695] <=  8'h6a;        memory[45696] <=  8'h6c;        memory[45697] <=  8'h6b;        memory[45698] <=  8'h63;        memory[45699] <=  8'h78;        memory[45700] <=  8'h20;        memory[45701] <=  8'h6a;        memory[45702] <=  8'h6b;        memory[45703] <=  8'h68;        memory[45704] <=  8'h61;        memory[45705] <=  8'h73;        memory[45706] <=  8'h76;        memory[45707] <=  8'h64;        memory[45708] <=  8'h6e;        memory[45709] <=  8'h20;        memory[45710] <=  8'h62;        memory[45711] <=  8'h6e;        memory[45712] <=  8'h6d;        memory[45713] <=  8'h6b;        memory[45714] <=  8'h77;        memory[45715] <=  8'h64;        memory[45716] <=  8'h6f;        memory[45717] <=  8'h77;        memory[45718] <=  8'h69;        memory[45719] <=  8'h6f;        memory[45720] <=  8'h75;        memory[45721] <=  8'h69;        memory[45722] <=  8'h68;        memory[45723] <=  8'h62;        memory[45724] <=  8'h6e;        memory[45725] <=  8'h6b;        memory[45726] <=  8'h77;        memory[45727] <=  8'h69;        memory[45728] <=  8'h6f;        memory[45729] <=  8'h75;        memory[45730] <=  8'h71;        memory[45731] <=  8'h69;        memory[45732] <=  8'h79;        memory[45733] <=  8'h67;        memory[45734] <=  8'h6a;        memory[45735] <=  8'h64;        memory[45736] <=  8'h61;        memory[45737] <=  8'h76;        memory[45738] <=  8'h62;        memory[45739] <=  8'h6e;        memory[45740] <=  8'h6b;        memory[45741] <=  8'h6f;        memory[45742] <=  8'h70;        memory[45743] <=  8'h64;        memory[45744] <=  8'h76;        memory[45745] <=  8'h69;        memory[45746] <=  8'h6f;        memory[45747] <=  8'h75;        memory[45748] <=  8'h69;        memory[45749] <=  8'h48;        memory[45750] <=  8'h42;        memory[45751] <=  8'h6b;        memory[45752] <=  8'h64;        memory[45753] <=  8'h6e;        memory[45754] <=  8'h6c;        memory[45755] <=  8'h71;        memory[45756] <=  8'h6b;        memory[45757] <=  8'h6d;        memory[45758] <=  8'h6a;        memory[45759] <=  8'h70;        memory[45760] <=  8'h69;        memory[45761] <=  8'h6f;        memory[45762] <=  8'h68;        memory[45763] <=  8'h65;        memory[45764] <=  8'h66;        memory[45765] <=  8'h75;        memory[45766] <=  8'h67;        memory[45767] <=  8'h69;        memory[45768] <=  8'h73;        memory[45769] <=  8'h61;        memory[45770] <=  8'h62;        memory[45771] <=  8'h64;        memory[45772] <=  8'h6b;        memory[45773] <=  8'h6a;        memory[45774] <=  8'h6b;        memory[45775] <=  8'h6c;        memory[45776] <=  8'h6a;        memory[45777] <=  8'h69;        memory[45778] <=  8'h73;        memory[45779] <=  8'h6f;        memory[45780] <=  8'h71;        memory[45781] <=  8'h68;        memory[45782] <=  8'h77;        memory[45783] <=  8'h67;        memory[45784] <=  8'h69;        memory[45785] <=  8'h79;        memory[45786] <=  8'h6a;        memory[45787] <=  8'h64;        memory[45788] <=  8'h76;        memory[45789] <=  8'h62;        memory[45790] <=  8'h6e;        memory[45791] <=  8'h61;        memory[45792] <=  8'h73;        memory[45793] <=  8'h66;        memory[45794] <=  8'h6c;        memory[45795] <=  8'h6b;        memory[45796] <=  8'h64;        memory[45797] <=  8'h6a;        memory[45798] <=  8'h68;        memory[45799] <=  8'h63;        memory[45800] <=  8'h67;        memory[45801] <=  8'h6a;        memory[45802] <=  8'h76;        memory[45803] <=  8'h73;        memory[45804] <=  8'h64;        memory[45805] <=  8'h62;        memory[45806] <=  8'h62;        memory[45807] <=  8'h61;        memory[45808] <=  8'h72;        memory[45809] <=  8'h62;        memory[45810] <=  8'h62;        memory[45811] <=  8'h73;        memory[45812] <=  8'h62;        memory[45813] <=  8'h67;        memory[45814] <=  8'h73;        memory[45815] <=  8'h66;        memory[45816] <=  8'h67;        memory[45817] <=  8'h61;        memory[45818] <=  8'h68;        memory[45819] <=  8'h66;        memory[45820] <=  8'h73;        memory[45821] <=  8'h68;        memory[45822] <=  8'h61;        memory[45823] <=  8'h66;        memory[45824] <=  8'h73;        memory[45825] <=  8'h66;        memory[45826] <=  8'h68;        memory[45827] <=  8'h61;        memory[45828] <=  8'h69;        memory[45829] <=  8'h64;        memory[45830] <=  8'h75;        memory[45831] <=  8'h67;        memory[45832] <=  8'h64;        memory[45833] <=  8'h77;        memory[45834] <=  8'h62;        memory[45835] <=  8'h61;        memory[45836] <=  8'h62;        memory[45837] <=  8'h72;        memory[45838] <=  8'h62;        memory[45839] <=  8'h61;        memory[45840] <=  8'h62;        memory[45841] <=  8'h62;        memory[45842] <=  8'h74;        memory[45843] <=  8'h62;        memory[45844] <=  8'h62;        memory[45845] <=  8'h62;        memory[45846] <=  8'h62;        memory[45847] <=  8'h62;        memory[45848] <=  8'h62;        memory[45849] <=  8'h62;        memory[45850] <=  8'h62;        memory[45851] <=  8'h61;        memory[45852] <=  8'h62;        memory[45853] <=  8'h62;        memory[45854] <=  8'h72;        memory[45855] <=  8'h74;        memory[45856] <=  8'h62;        memory[45857] <=  8'h62;        memory[45858] <=  8'h61;        memory[45859] <=  8'h62;        memory[45860] <=  8'h72;        memory[45861] <=  8'h62;        memory[45862] <=  8'h74;        memory[45863] <=  8'h62;        memory[45864] <=  8'h62;        memory[45865] <=  8'h62;        memory[45866] <=  8'h63;        memory[45867] <=  8'h61;        memory[45868] <=  8'h72;        memory[45869] <=  8'h74;        memory[45870] <=  8'h73;        memory[45871] <=  8'h62;        memory[45872] <=  8'h61;        memory[45873] <=  8'h72;        memory[45874] <=  8'h74;        memory[45875] <=  8'h74;        memory[45876] <=  8'h62;        memory[45877] <=  8'h61;        memory[45878] <=  8'h72;        memory[45879] <=  8'h74;        memory[45880] <=  8'h78;        memory[45881] <=  8'h61;        memory[45882] <=  8'h74;        memory[45883] <=  8'h6b;        memory[45884] <=  8'h73;        memory[45885] <=  8'h68;        memory[45886] <=  8'h63;        memory[45887] <=  8'h66;        memory[45888] <=  8'h69;        memory[45889] <=  8'h77;        memory[45890] <=  8'h68;        memory[45891] <=  8'h61;        memory[45892] <=  8'h74;        memory[45893] <=  8'h61;        memory[45894] <=  8'h6e;        memory[45895] <=  8'h61;        memory[45896] <=  8'h62;        memory[45897] <=  8'h61;        memory[45898] <=  8'h63;        memory[45899] <=  8'h61;        memory[45900] <=  8'h74;        memory[45901] <=  8'h61;        memory[45902] <=  8'h62;        memory[45903] <=  8'h61;        memory[45904] <=  8'h72;        memory[45905] <=  8'h63;        memory[45906] <=  8'h61;        memory[45907] <=  8'h68;        memory[45908] <=  8'h64;        memory[45909] <=  8'h75;        memory[45910] <=  8'h63;        memory[45911] <=  8'h74;        memory[45912] <=  8'h61;        memory[45913] <=  8'h64;        memory[45914] <=  8'h61;        memory[45915] <=  8'h61;        memory[45916] <=  8'h63;        memory[45917] <=  8'h61;        memory[45918] <=  8'h72;        memory[45919] <=  8'h63;        memory[45920] <=  8'h74;        memory[45921] <=  8'h72;        memory[45922] <=  8'h63;        memory[45923] <=  8'h61;        memory[45924] <=  8'h74;        memory[45925] <=  8'h72;        memory[45926] <=  8'h63;        memory[45927] <=  8'h61;        memory[45928] <=  8'h74;        memory[45929] <=  8'h63;        memory[45930] <=  8'h62;        memory[45931] <=  8'h61;        memory[45932] <=  8'h74;        memory[45933] <=  8'h62;        memory[45934] <=  8'h72;        memory[45935] <=  8'h63;        memory[45936] <=  8'h61;        memory[45937] <=  8'h74;        memory[45938] <=  8'h72;        memory[45939] <=  8'h6e;        memory[45940] <=  8'h62;        memory[45941] <=  8'h61;        memory[45942] <=  8'h63;        memory[45943] <=  8'h61;        memory[45944] <=  8'h74;        memory[45945] <=  8'h79;        memory[45946] <=  8'h73;        memory[45947] <=  8'h6e;        memory[45948] <=  8'h63;        memory[45949] <=  8'h74;        memory[45950] <=  8'h61;        memory[45951] <=  8'h6e;        memory[45952] <=  8'h62;        memory[45953] <=  8'h61;        memory[45954] <=  8'h63;        memory[45955] <=  8'h72;        memory[45956] <=  8'h6e;        memory[45957] <=  8'h74;        memory[45958] <=  8'h61;        memory[45959] <=  8'h62;        memory[45960] <=  8'h74;        memory[45961] <=  8'h6e;        memory[45962] <=  8'h61;        memory[45963] <=  8'h72;        memory[45964] <=  8'h62;        memory[45965] <=  8'h78;        memory[45966] <=  8'h74;        memory[45967] <=  8'h61;        memory[45968] <=  8'h72;        memory[45969] <=  8'h62;        memory[45970] <=  8'h61;        memory[45971] <=  8'h72;        memory[45972] <=  8'h74;        memory[45973] <=  8'h74;        memory[45974] <=  8'h62;        memory[45975] <=  8'h61;        memory[45976] <=  8'h72;        memory[45977] <=  8'h74;        memory[45978] <=  8'h78;        memory[45979] <=  8'h61;        memory[45980] <=  8'h74;        memory[45981] <=  8'h6b;        memory[45982] <=  8'h73;        memory[45983] <=  8'h68;        memory[45984] <=  8'h63;        memory[45985] <=  8'h66;        memory[45986] <=  8'h69;        memory[45987] <=  8'h77;        memory[45988] <=  8'h68;        memory[45989] <=  8'h61;        memory[45990] <=  8'h74;        memory[45991] <=  8'h61;        memory[45992] <=  8'h6e;        memory[45993] <=  8'h61;        memory[45994] <=  8'h62;        memory[45995] <=  8'h61;        memory[45996] <=  8'h63;        memory[45997] <=  8'h61;        memory[45998] <=  8'h74;        memory[45999] <=  8'h61;        memory[46000] <=  8'h62;        memory[46001] <=  8'h61;        memory[46002] <=  8'h72;        memory[46003] <=  8'h63;        memory[46004] <=  8'h61;        memory[46005] <=  8'h68;        memory[46006] <=  8'h64;        memory[46007] <=  8'h75;        memory[46008] <=  8'h63;        memory[46009] <=  8'h74;        memory[46010] <=  8'h61;        memory[46011] <=  8'h64;        memory[46012] <=  8'h61;        memory[46013] <=  8'h61;        memory[46014] <=  8'h63;        memory[46015] <=  8'h61;        memory[46016] <=  8'h72;        memory[46017] <=  8'h63;        memory[46018] <=  8'h74;        memory[46019] <=  8'h72;        memory[46020] <=  8'h63;        memory[46021] <=  8'h61;        memory[46022] <=  8'h74;        memory[46023] <=  8'h72;        memory[46024] <=  8'h63;        memory[46025] <=  8'h61;        memory[46026] <=  8'h74;        memory[46027] <=  8'h63;        memory[46028] <=  8'h62;        memory[46029] <=  8'h61;        memory[46030] <=  8'h74;        memory[46031] <=  8'h62;        memory[46032] <=  8'h72;        memory[46033] <=  8'h63;        memory[46034] <=  8'h61;        memory[46035] <=  8'h74;        memory[46036] <=  8'h72;        memory[46037] <=  8'h6e;        memory[46038] <=  8'h62;        memory[46039] <=  8'h61;        memory[46040] <=  8'h63;        memory[46041] <=  8'h61;        memory[46042] <=  8'h74;        memory[46043] <=  8'h79;        memory[46044] <=  8'h73;        memory[46045] <=  8'h6e;        memory[46046] <=  8'h63;        memory[46047] <=  8'h74;        memory[46048] <=  8'h61;        memory[46049] <=  8'h6e;        memory[46050] <=  8'h62;        memory[46051] <=  8'h61;        memory[46052] <=  8'h63;        memory[46053] <=  8'h72;        memory[46054] <=  8'h6e;        memory[46055] <=  8'h74;        memory[46056] <=  8'h61;        memory[46057] <=  8'h62;        memory[46058] <=  8'h74;        memory[46059] <=  8'h6e;        memory[46060] <=  8'h61;        memory[46061] <=  8'h72;        memory[46062] <=  8'h62;        memory[46063] <=  8'h78;        memory[46064] <=  8'h74;        memory[46065] <=  8'h61;        memory[46066] <=  8'h72;        memory[46067] <=  8'h62;        memory[46068] <=  8'h61;        memory[46069] <=  8'h72;        memory[46070] <=  8'h74;        memory[46071] <=  8'h74;        memory[46072] <=  8'h62;        memory[46073] <=  8'h61;        memory[46074] <=  8'h72;        memory[46075] <=  8'h74;        memory[46076] <=  8'h78;        memory[46077] <=  8'h61;        memory[46078] <=  8'h74;        memory[46079] <=  8'h6b;        memory[46080] <=  8'h73;        memory[46081] <=  8'h68;        memory[46082] <=  8'h63;        memory[46083] <=  8'h66;        memory[46084] <=  8'h69;        memory[46085] <=  8'h77;        memory[46086] <=  8'h68;        memory[46087] <=  8'h61;        memory[46088] <=  8'h74;        memory[46089] <=  8'h61;        memory[46090] <=  8'h6e;        memory[46091] <=  8'h61;        memory[46092] <=  8'h62;        memory[46093] <=  8'h61;        memory[46094] <=  8'h63;        memory[46095] <=  8'h61;        memory[46096] <=  8'h74;        memory[46097] <=  8'h61;        memory[46098] <=  8'h62;        memory[46099] <=  8'h61;        memory[46100] <=  8'h72;        memory[46101] <=  8'h63;        memory[46102] <=  8'h61;        memory[46103] <=  8'h68;        memory[46104] <=  8'h64;        memory[46105] <=  8'h75;        memory[46106] <=  8'h63;        memory[46107] <=  8'h74;        memory[46108] <=  8'h61;        memory[46109] <=  8'h64;        memory[46110] <=  8'h61;        memory[46111] <=  8'h61;        memory[46112] <=  8'h63;        memory[46113] <=  8'h61;        memory[46114] <=  8'h72;        memory[46115] <=  8'h63;        memory[46116] <=  8'h74;        memory[46117] <=  8'h72;        memory[46118] <=  8'h63;        memory[46119] <=  8'h61;        memory[46120] <=  8'h74;        memory[46121] <=  8'h72;        memory[46122] <=  8'h63;        memory[46123] <=  8'h61;        memory[46124] <=  8'h74;        memory[46125] <=  8'h63;        memory[46126] <=  8'h62;        memory[46127] <=  8'h61;        memory[46128] <=  8'h74;        memory[46129] <=  8'h62;        memory[46130] <=  8'h72;        memory[46131] <=  8'h63;        memory[46132] <=  8'h61;        memory[46133] <=  8'h74;        memory[46134] <=  8'h72;        memory[46135] <=  8'h6e;        memory[46136] <=  8'h62;        memory[46137] <=  8'h61;        memory[46138] <=  8'h63;        memory[46139] <=  8'h61;        memory[46140] <=  8'h74;        memory[46141] <=  8'h79;        memory[46142] <=  8'h73;        memory[46143] <=  8'h6e;        memory[46144] <=  8'h63;        memory[46145] <=  8'h74;        memory[46146] <=  8'h61;        memory[46147] <=  8'h6e;        memory[46148] <=  8'h62;        memory[46149] <=  8'h61;        memory[46150] <=  8'h63;        memory[46151] <=  8'h72;        memory[46152] <=  8'h6e;        memory[46153] <=  8'h74;        memory[46154] <=  8'h61;        memory[46155] <=  8'h62;        memory[46156] <=  8'h74;        memory[46157] <=  8'h6e;        memory[46158] <=  8'h61;        memory[46159] <=  8'h72;        memory[46160] <=  8'h62;        memory[46161] <=  8'h78;        memory[46162] <=  8'h74;        memory[46163] <=  8'h61;        memory[46164] <=  8'h72;        memory[46165] <=  8'h5d;        memory[46166] <=  8'h5d;        memory[46167] <=  8'h65;        memory[46168] <=  8'h66;        memory[46169] <=  8'h77;        memory[46170] <=  8'h65;        memory[46171] <=  8'h5d;        memory[46172] <=  8'h65;        memory[46173] <=  8'h67;        memory[46174] <=  8'h73;        memory[46175] <=  8'h67;        memory[46176] <=  8'h66;        memory[46177] <=  8'h62;        memory[46178] <=  8'h61;        memory[46179] <=  8'h72;        memory[46180] <=  8'h74;        memory[46181] <=  8'h74;        memory[46182] <=  8'h62;        memory[46183] <=  8'h61;        memory[46184] <=  8'h72;        memory[46185] <=  8'h74;        memory[46186] <=  8'h78;        memory[46187] <=  8'h61;        memory[46188] <=  8'h74;        memory[46189] <=  8'h6b;        memory[46190] <=  8'h73;        memory[46191] <=  8'h68;        memory[46192] <=  8'h63;        memory[46193] <=  8'h66;        memory[46194] <=  8'h69;        memory[46195] <=  8'h77;        memory[46196] <=  8'h68;        memory[46197] <=  8'h61;        memory[46198] <=  8'h74;        memory[46199] <=  8'h61;        memory[46200] <=  8'h6e;        memory[46201] <=  8'h61;        memory[46202] <=  8'h62;        memory[46203] <=  8'h61;        memory[46204] <=  8'h63;        memory[46205] <=  8'h61;        memory[46206] <=  8'h74;        memory[46207] <=  8'h61;        memory[46208] <=  8'h62;        memory[46209] <=  8'h61;        memory[46210] <=  8'h72;        memory[46211] <=  8'h63;        memory[46212] <=  8'h61;        memory[46213] <=  8'h68;        memory[46214] <=  8'h64;        memory[46215] <=  8'h75;        memory[46216] <=  8'h63;        memory[46217] <=  8'h74;        memory[46218] <=  8'h61;        memory[46219] <=  8'h64;        memory[46220] <=  8'h61;        memory[46221] <=  8'h61;        memory[46222] <=  8'h63;        memory[46223] <=  8'h61;        memory[46224] <=  8'h72;        memory[46225] <=  8'h63;        memory[46226] <=  8'h74;        memory[46227] <=  8'h72;        memory[46228] <=  8'h63;        memory[46229] <=  8'h61;        memory[46230] <=  8'h74;        memory[46231] <=  8'h72;        memory[46232] <=  8'h63;        memory[46233] <=  8'h61;        memory[46234] <=  8'h74;        memory[46235] <=  8'h63;        memory[46236] <=  8'h62;        memory[46237] <=  8'h61;        memory[46238] <=  8'h74;        memory[46239] <=  8'h62;        memory[46240] <=  8'h72;        memory[46241] <=  8'h63;        memory[46242] <=  8'h61;        memory[46243] <=  8'h74;        memory[46244] <=  8'h72;        memory[46245] <=  8'h6e;        memory[46246] <=  8'h62;        memory[46247] <=  8'h61;        memory[46248] <=  8'h63;        memory[46249] <=  8'h61;        memory[46250] <=  8'h74;        memory[46251] <=  8'h79;        memory[46252] <=  8'h73;        memory[46253] <=  8'h6e;        memory[46254] <=  8'h63;        memory[46255] <=  8'h74;        memory[46256] <=  8'h61;        memory[46257] <=  8'h6e;        memory[46258] <=  8'h62;        memory[46259] <=  8'h61;        memory[46260] <=  8'h63;        memory[46261] <=  8'h72;        memory[46262] <=  8'h6e;        memory[46263] <=  8'h74;        memory[46264] <=  8'h61;        memory[46265] <=  8'h62;        memory[46266] <=  8'h74;        memory[46267] <=  8'h6e;        memory[46268] <=  8'h61;        memory[46269] <=  8'h72;        memory[46270] <=  8'h62;        memory[46271] <=  8'h78;        memory[46272] <=  8'h74;        memory[46273] <=  8'h61;        memory[46274] <=  8'h72;        memory[46275] <=  8'h62;        memory[46276] <=  8'h61;        memory[46277] <=  8'h72;        memory[46278] <=  8'h74;        memory[46279] <=  8'h74;        memory[46280] <=  8'h62;        memory[46281] <=  8'h61;        memory[46282] <=  8'h72;        memory[46283] <=  8'h74;        memory[46284] <=  8'h78;        memory[46285] <=  8'h61;        memory[46286] <=  8'h74;        memory[46287] <=  8'h6b;        memory[46288] <=  8'h73;        memory[46289] <=  8'h68;        memory[46290] <=  8'h63;        memory[46291] <=  8'h66;        memory[46292] <=  8'h69;        memory[46293] <=  8'h77;        memory[46294] <=  8'h68;        memory[46295] <=  8'h61;        memory[46296] <=  8'h74;        memory[46297] <=  8'h61;        memory[46298] <=  8'h6e;        memory[46299] <=  8'h61;        memory[46300] <=  8'h62;        memory[46301] <=  8'h61;        memory[46302] <=  8'h63;        memory[46303] <=  8'h61;        memory[46304] <=  8'h74;        memory[46305] <=  8'h61;        memory[46306] <=  8'h62;        memory[46307] <=  8'h61;        memory[46308] <=  8'h72;        memory[46309] <=  8'h63;        memory[46310] <=  8'h61;        memory[46311] <=  8'h68;        memory[46312] <=  8'h64;        memory[46313] <=  8'h75;        memory[46314] <=  8'h63;        memory[46315] <=  8'h74;        memory[46316] <=  8'h61;        memory[46317] <=  8'h64;        memory[46318] <=  8'h61;        memory[46319] <=  8'h61;        memory[46320] <=  8'h63;        memory[46321] <=  8'h61;        memory[46322] <=  8'h72;        memory[46323] <=  8'h63;        memory[46324] <=  8'h74;        memory[46325] <=  8'h72;        memory[46326] <=  8'h63;        memory[46327] <=  8'h61;        memory[46328] <=  8'h74;        memory[46329] <=  8'h72;        memory[46330] <=  8'h63;        memory[46331] <=  8'h61;        memory[46332] <=  8'h74;        memory[46333] <=  8'h63;        memory[46334] <=  8'h62;        memory[46335] <=  8'h61;        memory[46336] <=  8'h74;        memory[46337] <=  8'h62;        memory[46338] <=  8'h72;        memory[46339] <=  8'h63;        memory[46340] <=  8'h61;        memory[46341] <=  8'h74;        memory[46342] <=  8'h72;        memory[46343] <=  8'h6e;        memory[46344] <=  8'h62;        memory[46345] <=  8'h61;        memory[46346] <=  8'h63;        memory[46347] <=  8'h61;        memory[46348] <=  8'h74;        memory[46349] <=  8'h79;        memory[46350] <=  8'h73;        memory[46351] <=  8'h6e;        memory[46352] <=  8'h63;        memory[46353] <=  8'h74;        memory[46354] <=  8'h61;        memory[46355] <=  8'h6e;        memory[46356] <=  8'h62;        memory[46357] <=  8'h61;        memory[46358] <=  8'h63;        memory[46359] <=  8'h72;        memory[46360] <=  8'h6e;        memory[46361] <=  8'h74;        memory[46362] <=  8'h61;        memory[46363] <=  8'h62;        memory[46364] <=  8'h74;        memory[46365] <=  8'h6e;        memory[46366] <=  8'h61;        memory[46367] <=  8'h72;        memory[46368] <=  8'h62;        memory[46369] <=  8'h78;        memory[46370] <=  8'h74;        memory[46371] <=  8'h61;        memory[46372] <=  8'h72;        memory[46373] <=  8'h64;        memory[46374] <=  8'h66;        memory[46375] <=  8'h73;        memory[46376] <=  8'h67;        memory[46377] <=  8'h76;        memory[46378] <=  8'h68;        memory[46379] <=  8'h62;        memory[46380] <=  8'h6b;        memory[46381] <=  8'h6a;        memory[46382] <=  8'h6e;        memory[46383] <=  8'h6d;        memory[46384] <=  8'h62;        memory[46385] <=  8'h76;        memory[46386] <=  8'h78;        memory[46387] <=  8'h63;        memory[46388] <=  8'h73;        memory[46389] <=  8'h66;        memory[46390] <=  8'h72;        memory[46391] <=  8'h74;        memory[46392] <=  8'h79;        memory[46393] <=  8'h75;        memory[46394] <=  8'h6a;        memory[46395] <=  8'h6e;        memory[46396] <=  8'h62;        memory[46397] <=  8'h76;        memory[46398] <=  8'h63;        memory[46399] <=  8'h64;        memory[46400] <=  8'h74;        memory[46401] <=  8'h79;        memory[46402] <=  8'h75;        memory[46403] <=  8'h69;        memory[46404] <=  8'h6b;        memory[46405] <=  8'h6d;        memory[46406] <=  8'h6e;        memory[46407] <=  8'h62;        memory[46408] <=  8'h76;        memory[46409] <=  8'h63;        memory[46410] <=  8'h78;        memory[46411] <=  8'h73;        memory[46412] <=  8'h64;        memory[46413] <=  8'h72;        memory[46414] <=  8'h74;        memory[46415] <=  8'h79;        memory[46416] <=  8'h75;        memory[46417] <=  8'h69;        memory[46418] <=  8'h6b;        memory[46419] <=  8'h6d;        memory[46420] <=  8'h6e;        memory[46421] <=  8'h62;        memory[46422] <=  8'h76;        memory[46423] <=  8'h63;        memory[46424] <=  8'h73;        memory[46425] <=  8'h77;        memory[46426] <=  8'h33;        memory[46427] <=  8'h34;        memory[46428] <=  8'h35;        memory[46429] <=  8'h36;        memory[46430] <=  8'h37;        memory[46431] <=  8'h38;        memory[46432] <=  8'h69;        memory[46433] <=  8'h6b;        memory[46434] <=  8'h6d;        memory[46435] <=  8'h6e;        memory[46436] <=  8'h62;        memory[46437] <=  8'h76;        memory[46438] <=  8'h63;        memory[46439] <=  8'h64;        memory[46440] <=  8'h65;        memory[46441] <=  8'h72;        memory[46442] <=  8'h36;        memory[46443] <=  8'h37;        memory[46444] <=  8'h38;        memory[46445] <=  8'h69;        memory[46446] <=  8'h6f;        memory[46447] <=  8'h6b;        memory[46448] <=  8'h6a;        memory[46449] <=  8'h6e;        memory[46450] <=  8'h62;        memory[46451] <=  8'h76;        memory[46452] <=  8'h63;        memory[46453] <=  8'h64;        memory[46454] <=  8'h72;        memory[46455] <=  8'h74;        memory[46456] <=  8'h79;        memory[46457] <=  8'h75;        memory[46458] <=  8'h73;        memory[46459] <=  8'h6a;        memory[46460] <=  8'h63;        memory[46461] <=  8'h6e;        memory[46462] <=  8'h62;        memory[46463] <=  8'h64;        memory[46464] <=  8'h66;        memory[46465] <=  8'h73;        memory[46466] <=  8'h74;        memory[46467] <=  8'h79;        memory[46468] <=  8'h75;        memory[46469] <=  8'h61;        memory[46470] <=  8'h69;        memory[46471] <=  8'h6b;        memory[46472] <=  8'h78;        memory[46473] <=  8'h6d;        memory[46474] <=  8'h6e;        memory[46475] <=  8'h73;        memory[46476] <=  8'h6a;        memory[46477] <=  8'h6f;        memory[46478] <=  8'h64;        memory[46479] <=  8'h6c;        memory[46480] <=  8'h63;        memory[46481] <=  8'h78;        memory[46482] <=  8'h62;        memory[46483] <=  8'h61;        memory[46484] <=  8'h72;        memory[46485] <=  8'h74;        memory[46486] <=  8'h78;        memory[46487] <=  8'h61;        memory[46488] <=  8'h74;        memory[46489] <=  8'h6b;        memory[46490] <=  8'h73;        memory[46491] <=  8'h68;        memory[46492] <=  8'h63;        memory[46493] <=  8'h66;        memory[46494] <=  8'h69;        memory[46495] <=  8'h77;        memory[46496] <=  8'h68;        memory[46497] <=  8'h61;        memory[46498] <=  8'h74;        memory[46499] <=  8'h61;        memory[46500] <=  8'h6e;        memory[46501] <=  8'h61;        memory[46502] <=  8'h62;        memory[46503] <=  8'h61;        memory[46504] <=  8'h63;        memory[46505] <=  8'h61;        memory[46506] <=  8'h74;        memory[46507] <=  8'h61;        memory[46508] <=  8'h62;        memory[46509] <=  8'h61;        memory[46510] <=  8'h72;        memory[46511] <=  8'h63;        memory[46512] <=  8'h61;        memory[46513] <=  8'h68;        memory[46514] <=  8'h64;        memory[46515] <=  8'h75;        memory[46516] <=  8'h63;        memory[46517] <=  8'h74;        memory[46518] <=  8'h61;        memory[46519] <=  8'h64;        memory[46520] <=  8'h61;        memory[46521] <=  8'h61;        memory[46522] <=  8'h63;        memory[46523] <=  8'h61;        memory[46524] <=  8'h72;        memory[46525] <=  8'h62;        memory[46526] <=  8'h61;        memory[46527] <=  8'h72;        memory[46528] <=  8'h74;        memory[46529] <=  8'h78;        memory[46530] <=  8'h61;        memory[46531] <=  8'h74;        memory[46532] <=  8'h6b;        memory[46533] <=  8'h73;        memory[46534] <=  8'h68;        memory[46535] <=  8'h63;        memory[46536] <=  8'h66;        memory[46537] <=  8'h69;        memory[46538] <=  8'h77;        memory[46539] <=  8'h68;        memory[46540] <=  8'h61;        memory[46541] <=  8'h74;        memory[46542] <=  8'h61;        memory[46543] <=  8'h6e;        memory[46544] <=  8'h61;        memory[46545] <=  8'h62;        memory[46546] <=  8'h61;        memory[46547] <=  8'h63;        memory[46548] <=  8'h61;        memory[46549] <=  8'h74;        memory[46550] <=  8'h61;        memory[46551] <=  8'h62;        memory[46552] <=  8'h61;        memory[46553] <=  8'h72;        memory[46554] <=  8'h63;        memory[46555] <=  8'h61;        memory[46556] <=  8'h68;        memory[46557] <=  8'h64;        memory[46558] <=  8'h75;        memory[46559] <=  8'h63;        memory[46560] <=  8'h74;        memory[46561] <=  8'h61;        memory[46562] <=  8'h64;        memory[46563] <=  8'h61;        memory[46564] <=  8'h61;        memory[46565] <=  8'h63;        memory[46566] <=  8'h61;        memory[46567] <=  8'h72;        memory[46568] <=  8'h62;        memory[46569] <=  8'h61;        memory[46570] <=  8'h72;        memory[46571] <=  8'h74;        memory[46572] <=  8'h78;        memory[46573] <=  8'h61;        memory[46574] <=  8'h74;        memory[46575] <=  8'h6b;        memory[46576] <=  8'h73;        memory[46577] <=  8'h68;        memory[46578] <=  8'h63;        memory[46579] <=  8'h66;        memory[46580] <=  8'h69;        memory[46581] <=  8'h77;        memory[46582] <=  8'h68;        memory[46583] <=  8'h61;        memory[46584] <=  8'h74;        memory[46585] <=  8'h61;        memory[46586] <=  8'h6e;        memory[46587] <=  8'h61;        memory[46588] <=  8'h62;        memory[46589] <=  8'h61;        memory[46590] <=  8'h63;        memory[46591] <=  8'h61;        memory[46592] <=  8'h74;        memory[46593] <=  8'h61;        memory[46594] <=  8'h62;        memory[46595] <=  8'h61;        memory[46596] <=  8'h72;        memory[46597] <=  8'h63;        memory[46598] <=  8'h61;        memory[46599] <=  8'h68;        memory[46600] <=  8'h64;        memory[46601] <=  8'h75;        memory[46602] <=  8'h63;        memory[46603] <=  8'h74;        memory[46604] <=  8'h61;        memory[46605] <=  8'h64;        memory[46606] <=  8'h61;        memory[46607] <=  8'h61;        memory[46608] <=  8'h63;        memory[46609] <=  8'h61;        memory[46610] <=  8'h72;        memory[46611] <=  8'h62;        memory[46612] <=  8'h61;        memory[46613] <=  8'h72;        memory[46614] <=  8'h74;        memory[46615] <=  8'h78;        memory[46616] <=  8'h61;        memory[46617] <=  8'h74;        memory[46618] <=  8'h6b;        memory[46619] <=  8'h73;        memory[46620] <=  8'h68;        memory[46621] <=  8'h63;        memory[46622] <=  8'h66;        memory[46623] <=  8'h69;        memory[46624] <=  8'h77;        memory[46625] <=  8'h68;        memory[46626] <=  8'h61;        memory[46627] <=  8'h74;        memory[46628] <=  8'h61;        memory[46629] <=  8'h6e;        memory[46630] <=  8'h61;        memory[46631] <=  8'h62;        memory[46632] <=  8'h61;        memory[46633] <=  8'h63;        memory[46634] <=  8'h61;        memory[46635] <=  8'h74;        memory[46636] <=  8'h61;        memory[46637] <=  8'h62;        memory[46638] <=  8'h61;        memory[46639] <=  8'h72;        memory[46640] <=  8'h63;        memory[46641] <=  8'h61;        memory[46642] <=  8'h68;        memory[46643] <=  8'h64;        memory[46644] <=  8'h75;        memory[46645] <=  8'h63;        memory[46646] <=  8'h74;        memory[46647] <=  8'h61;        memory[46648] <=  8'h64;        memory[46649] <=  8'h61;        memory[46650] <=  8'h61;        memory[46651] <=  8'h63;        memory[46652] <=  8'h61;        memory[46653] <=  8'h72;        memory[46654] <=  8'h62;        memory[46655] <=  8'h61;        memory[46656] <=  8'h72;        memory[46657] <=  8'h74;        memory[46658] <=  8'h78;        memory[46659] <=  8'h61;        memory[46660] <=  8'h74;        memory[46661] <=  8'h6b;        memory[46662] <=  8'h73;        memory[46663] <=  8'h68;        memory[46664] <=  8'h63;        memory[46665] <=  8'h66;        memory[46666] <=  8'h69;        memory[46667] <=  8'h77;        memory[46668] <=  8'h68;        memory[46669] <=  8'h61;        memory[46670] <=  8'h74;        memory[46671] <=  8'h61;        memory[46672] <=  8'h6e;        memory[46673] <=  8'h61;        memory[46674] <=  8'h62;        memory[46675] <=  8'h61;        memory[46676] <=  8'h63;        memory[46677] <=  8'h61;        memory[46678] <=  8'h74;        memory[46679] <=  8'h61;        memory[46680] <=  8'h62;        memory[46681] <=  8'h61;        memory[46682] <=  8'h72;        memory[46683] <=  8'h63;        memory[46684] <=  8'h61;        memory[46685] <=  8'h68;        memory[46686] <=  8'h64;        memory[46687] <=  8'h75;        memory[46688] <=  8'h63;        memory[46689] <=  8'h74;        memory[46690] <=  8'h61;        memory[46691] <=  8'h64;        memory[46692] <=  8'h61;        memory[46693] <=  8'h61;        memory[46694] <=  8'h63;        memory[46695] <=  8'h61;        memory[46696] <=  8'h72;        memory[46697] <=  8'h62;        memory[46698] <=  8'h61;        memory[46699] <=  8'h72;        memory[46700] <=  8'h74;        memory[46701] <=  8'h78;        memory[46702] <=  8'h61;        memory[46703] <=  8'h74;        memory[46704] <=  8'h6b;        memory[46705] <=  8'h73;        memory[46706] <=  8'h68;        memory[46707] <=  8'h63;        memory[46708] <=  8'h66;        memory[46709] <=  8'h69;        memory[46710] <=  8'h77;        memory[46711] <=  8'h68;        memory[46712] <=  8'h61;        memory[46713] <=  8'h74;        memory[46714] <=  8'h61;        memory[46715] <=  8'h6e;        memory[46716] <=  8'h61;        memory[46717] <=  8'h62;        memory[46718] <=  8'h61;        memory[46719] <=  8'h63;        memory[46720] <=  8'h61;        memory[46721] <=  8'h74;        memory[46722] <=  8'h61;        memory[46723] <=  8'h62;        memory[46724] <=  8'h61;        memory[46725] <=  8'h72;        memory[46726] <=  8'h63;        memory[46727] <=  8'h61;        memory[46728] <=  8'h68;        memory[46729] <=  8'h64;        memory[46730] <=  8'h75;        memory[46731] <=  8'h63;        memory[46732] <=  8'h74;        memory[46733] <=  8'h61;        memory[46734] <=  8'h64;        memory[46735] <=  8'h61;        memory[46736] <=  8'h61;        memory[46737] <=  8'h63;        memory[46738] <=  8'h61;        memory[46739] <=  8'h72;        memory[46740] <=  8'h62;        memory[46741] <=  8'h61;        memory[46742] <=  8'h72;        memory[46743] <=  8'h74;        memory[46744] <=  8'h78;        memory[46745] <=  8'h61;        memory[46746] <=  8'h74;        memory[46747] <=  8'h6b;        memory[46748] <=  8'h73;        memory[46749] <=  8'h68;        memory[46750] <=  8'h63;        memory[46751] <=  8'h66;        memory[46752] <=  8'h69;        memory[46753] <=  8'h77;        memory[46754] <=  8'h68;        memory[46755] <=  8'h61;        memory[46756] <=  8'h74;        memory[46757] <=  8'h61;        memory[46758] <=  8'h6e;        memory[46759] <=  8'h61;        memory[46760] <=  8'h62;        memory[46761] <=  8'h61;        memory[46762] <=  8'h63;        memory[46763] <=  8'h61;        memory[46764] <=  8'h74;        memory[46765] <=  8'h61;        memory[46766] <=  8'h62;        memory[46767] <=  8'h61;        memory[46768] <=  8'h72;        memory[46769] <=  8'h63;        memory[46770] <=  8'h61;        memory[46771] <=  8'h68;        memory[46772] <=  8'h64;        memory[46773] <=  8'h75;        memory[46774] <=  8'h63;        memory[46775] <=  8'h74;        memory[46776] <=  8'h61;        memory[46777] <=  8'h64;        memory[46778] <=  8'h61;        memory[46779] <=  8'h61;        memory[46780] <=  8'h63;        memory[46781] <=  8'h61;        memory[46782] <=  8'h72;        memory[46783] <=  8'h62;        memory[46784] <=  8'h61;        memory[46785] <=  8'h72;        memory[46786] <=  8'h74;        memory[46787] <=  8'h78;        memory[46788] <=  8'h61;        memory[46789] <=  8'h74;        memory[46790] <=  8'h6b;        memory[46791] <=  8'h73;        memory[46792] <=  8'h68;        memory[46793] <=  8'h63;        memory[46794] <=  8'h66;        memory[46795] <=  8'h69;        memory[46796] <=  8'h77;        memory[46797] <=  8'h68;        memory[46798] <=  8'h61;        memory[46799] <=  8'h74;        memory[46800] <=  8'h61;        memory[46801] <=  8'h6e;        memory[46802] <=  8'h61;        memory[46803] <=  8'h62;        memory[46804] <=  8'h61;        memory[46805] <=  8'h63;        memory[46806] <=  8'h61;        memory[46807] <=  8'h74;        memory[46808] <=  8'h61;        memory[46809] <=  8'h62;        memory[46810] <=  8'h61;        memory[46811] <=  8'h72;        memory[46812] <=  8'h63;        memory[46813] <=  8'h61;        memory[46814] <=  8'h68;        memory[46815] <=  8'h64;        memory[46816] <=  8'h75;        memory[46817] <=  8'h63;        memory[46818] <=  8'h74;        memory[46819] <=  8'h61;        memory[46820] <=  8'h64;        memory[46821] <=  8'h61;        memory[46822] <=  8'h61;        memory[46823] <=  8'h63;        memory[46824] <=  8'h61;        memory[46825] <=  8'h72;        memory[46826] <=  8'h62;        memory[46827] <=  8'h61;        memory[46828] <=  8'h72;        memory[46829] <=  8'h74;        memory[46830] <=  8'h78;        memory[46831] <=  8'h61;        memory[46832] <=  8'h74;        memory[46833] <=  8'h6b;        memory[46834] <=  8'h73;        memory[46835] <=  8'h68;        memory[46836] <=  8'h63;        memory[46837] <=  8'h66;        memory[46838] <=  8'h69;        memory[46839] <=  8'h77;        memory[46840] <=  8'h68;        memory[46841] <=  8'h61;        memory[46842] <=  8'h74;        memory[46843] <=  8'h61;        memory[46844] <=  8'h6e;        memory[46845] <=  8'h61;        memory[46846] <=  8'h62;        memory[46847] <=  8'h61;        memory[46848] <=  8'h63;        memory[46849] <=  8'h61;        memory[46850] <=  8'h74;        memory[46851] <=  8'h61;        memory[46852] <=  8'h62;        memory[46853] <=  8'h61;        memory[46854] <=  8'h72;        memory[46855] <=  8'h63;        memory[46856] <=  8'h61;        memory[46857] <=  8'h68;        memory[46858] <=  8'h64;        memory[46859] <=  8'h75;        memory[46860] <=  8'h63;        memory[46861] <=  8'h74;        memory[46862] <=  8'h61;        memory[46863] <=  8'h64;        memory[46864] <=  8'h61;        memory[46865] <=  8'h61;        memory[46866] <=  8'h63;        memory[46867] <=  8'h61;        memory[46868] <=  8'h72;        memory[46869] <=  8'h62;        memory[46870] <=  8'h61;        memory[46871] <=  8'h72;        memory[46872] <=  8'h74;        memory[46873] <=  8'h74;        memory[46874] <=  8'h62;        memory[46875] <=  8'h61;        memory[46876] <=  8'h72;        memory[46877] <=  8'h74;        memory[46878] <=  8'h78;        memory[46879] <=  8'h61;        memory[46880] <=  8'h74;        memory[46881] <=  8'h6b;        memory[46882] <=  8'h73;        memory[46883] <=  8'h68;        memory[46884] <=  8'h63;        memory[46885] <=  8'h66;        memory[46886] <=  8'h69;        memory[46887] <=  8'h77;        memory[46888] <=  8'h68;        memory[46889] <=  8'h61;        memory[46890] <=  8'h74;        memory[46891] <=  8'h61;        memory[46892] <=  8'h6e;        memory[46893] <=  8'h61;        memory[46894] <=  8'h62;        memory[46895] <=  8'h61;        memory[46896] <=  8'h63;        memory[46897] <=  8'h61;        memory[46898] <=  8'h74;        memory[46899] <=  8'h61;        memory[46900] <=  8'h62;        memory[46901] <=  8'h61;        memory[46902] <=  8'h72;        memory[46903] <=  8'h63;        memory[46904] <=  8'h61;        memory[46905] <=  8'h68;        memory[46906] <=  8'h64;        memory[46907] <=  8'h75;        memory[46908] <=  8'h63;        memory[46909] <=  8'h74;        memory[46910] <=  8'h61;        memory[46911] <=  8'h64;        memory[46912] <=  8'h61;        memory[46913] <=  8'h61;        memory[46914] <=  8'h63;        memory[46915] <=  8'h61;        memory[46916] <=  8'h72;        memory[46917] <=  8'h63;        memory[46918] <=  8'h74;        memory[46919] <=  8'h72;        memory[46920] <=  8'h63;        memory[46921] <=  8'h61;        memory[46922] <=  8'h74;        memory[46923] <=  8'h72;        memory[46924] <=  8'h63;        memory[46925] <=  8'h61;        memory[46926] <=  8'h74;        memory[46927] <=  8'h63;        memory[46928] <=  8'h62;        memory[46929] <=  8'h61;        memory[46930] <=  8'h74;        memory[46931] <=  8'h62;        memory[46932] <=  8'h72;        memory[46933] <=  8'h63;        memory[46934] <=  8'h61;        memory[46935] <=  8'h72;        memory[46936] <=  8'h62;        memory[46937] <=  8'h78;        memory[46938] <=  8'h74;        memory[46939] <=  8'h61;        memory[46940] <=  8'h72;        memory[46941] <=  8'h64;        memory[46942] <=  8'h66;        memory[46943] <=  8'h73;        memory[46944] <=  8'h67;        memory[46945] <=  8'h76;        memory[46946] <=  8'h68;        memory[46947] <=  8'h62;        memory[46948] <=  8'h6b;        memory[46949] <=  8'h6a;        memory[46950] <=  8'h6e;        memory[46951] <=  8'h6d;        memory[46952] <=  8'h62;        memory[46953] <=  8'h76;        memory[46954] <=  8'h78;        memory[46955] <=  8'h63;        memory[46956] <=  8'h73;        memory[46957] <=  8'h66;        memory[46958] <=  8'h72;        memory[46959] <=  8'h74;        memory[46960] <=  8'h79;        memory[46961] <=  8'h75;        memory[46962] <=  8'h6a;        memory[46963] <=  8'h6e;        memory[46964] <=  8'h62;        memory[46965] <=  8'h76;        memory[46966] <=  8'h63;        memory[46967] <=  8'h64;        memory[46968] <=  8'h74;        memory[46969] <=  8'h79;        memory[46970] <=  8'h75;        memory[46971] <=  8'h69;        memory[46972] <=  8'h6b;        memory[46973] <=  8'h6d;        memory[46974] <=  8'h6e;        memory[46975] <=  8'h62;        memory[46976] <=  8'h76;        memory[46977] <=  8'h63;        memory[46978] <=  8'h78;        memory[46979] <=  8'h73;        memory[46980] <=  8'h64;        memory[46981] <=  8'h72;        memory[46982] <=  8'h74;        memory[46983] <=  8'h79;        memory[46984] <=  8'h75;        memory[46985] <=  8'h69;        memory[46986] <=  8'h6b;        memory[46987] <=  8'h6d;        memory[46988] <=  8'h6e;        memory[46989] <=  8'h62;        memory[46990] <=  8'h76;        memory[46991] <=  8'h63;        memory[46992] <=  8'h73;        memory[46993] <=  8'h77;        memory[46994] <=  8'h33;        memory[46995] <=  8'h34;        memory[46996] <=  8'h35;        memory[46997] <=  8'h36;        memory[46998] <=  8'h37;        memory[46999] <=  8'h38;        memory[47000] <=  8'h69;        memory[47001] <=  8'h6b;        memory[47002] <=  8'h6d;        memory[47003] <=  8'h6e;        memory[47004] <=  8'h62;        memory[47005] <=  8'h76;        memory[47006] <=  8'h63;        memory[47007] <=  8'h64;        memory[47008] <=  8'h65;        memory[47009] <=  8'h72;        memory[47010] <=  8'h36;        memory[47011] <=  8'h37;        memory[47012] <=  8'h38;        memory[47013] <=  8'h69;        memory[47014] <=  8'h6f;        memory[47015] <=  8'h6b;        memory[47016] <=  8'h6a;        memory[47017] <=  8'h6e;        memory[47018] <=  8'h62;        memory[47019] <=  8'h76;        memory[47020] <=  8'h63;        memory[47021] <=  8'h64;        memory[47022] <=  8'h72;        memory[47023] <=  8'h74;        memory[47024] <=  8'h79;        memory[47025] <=  8'h75;        memory[47026] <=  8'h73;        memory[47027] <=  8'h6a;        memory[47028] <=  8'h63;        memory[47029] <=  8'h6e;        memory[47030] <=  8'h62;        memory[47031] <=  8'h64;        memory[47032] <=  8'h66;        memory[47033] <=  8'h73;        memory[47034] <=  8'h74;        memory[47035] <=  8'h79;        memory[47036] <=  8'h75;        memory[47037] <=  8'h61;        memory[47038] <=  8'h69;        memory[47039] <=  8'h6b;        memory[47040] <=  8'h78;        memory[47041] <=  8'h6d;        memory[47042] <=  8'h6e;        memory[47043] <=  8'h73;        memory[47044] <=  8'h6a;        memory[47045] <=  8'h6f;        memory[47046] <=  8'h64;        memory[47047] <=  8'h6c;        memory[47048] <=  8'h63;        memory[47049] <=  8'h78;        memory[47050] <=  8'h2c;        memory[47051] <=  8'h6d;        memory[47052] <=  8'h73;        memory[47053] <=  8'h6b;        memory[47054] <=  8'h64;        memory[47055] <=  8'h6c;        memory[47056] <=  8'h70;        memory[47057] <=  8'h5b;        memory[47058] <=  8'h3b;        memory[47059] <=  8'h73;        memory[47060] <=  8'h6c;        memory[47061] <=  8'h64;        memory[47062] <=  8'h70;        memory[47063] <=  8'h76;        memory[47064] <=  8'h63;        memory[47065] <=  8'h5b;        memory[47066] <=  8'h78;        memory[47067] <=  8'h76;        memory[47068] <=  8'h63;        memory[47069] <=  8'h5b;        memory[47070] <=  8'h78;        memory[47071] <=  8'h70;        memory[47072] <=  8'h6f;        memory[47073] <=  8'h20;        memory[47074] <=  8'h62;        memory[47075] <=  8'h61;        memory[47076] <=  8'h72;        memory[47077] <=  8'h74;        memory[47078] <=  8'h74;        memory[47079] <=  8'h62;        memory[47080] <=  8'h61;        memory[47081] <=  8'h72;        memory[47082] <=  8'h74;        memory[47083] <=  8'h78;        memory[47084] <=  8'h61;        memory[47085] <=  8'h74;        memory[47086] <=  8'h6b;        memory[47087] <=  8'h73;        memory[47088] <=  8'h68;        memory[47089] <=  8'h63;        memory[47090] <=  8'h66;        memory[47091] <=  8'h69;        memory[47092] <=  8'h77;        memory[47093] <=  8'h68;        memory[47094] <=  8'h61;        memory[47095] <=  8'h69;        memory[47096] <=  8'h6a;        memory[47097] <=  8'h78;        memory[47098] <=  8'h5d;        memory[47099] <=  8'h65;        memory[47100] <=  8'h6b;        memory[47101] <=  8'h6f;        memory[47102] <=  8'h39;        memory[47103] <=  8'h64;        memory[47104] <=  8'h75;        memory[47105] <=  8'h38;        memory[47106] <=  8'h79;        memory[47107] <=  8'h20;        memory[47108] <=  8'h37;        memory[47109] <=  8'h63;        memory[47110] <=  8'h67;        memory[47111] <=  8'h78;        memory[47112] <=  8'h63;        memory[47113] <=  8'h75;        memory[47114] <=  8'h68;        memory[47115] <=  8'h69;        memory[47116] <=  8'h6a;        memory[47117] <=  8'h77;        memory[47118] <=  8'h69;        memory[47119] <=  8'h64;        memory[47120] <=  8'h66;        memory[47121] <=  8'h68;        memory[47122] <=  8'h75;        memory[47123] <=  8'h76;        memory[47124] <=  8'h64;        memory[47125] <=  8'h62;        memory[47126] <=  8'h66;        memory[47127] <=  8'h6a;        memory[47128] <=  8'h6e;        memory[47129] <=  8'h6b;        memory[47130] <=  8'h6a;        memory[47131] <=  8'h65;        memory[47132] <=  8'h38;        memory[47133] <=  8'h66;        memory[47134] <=  8'h37;        memory[47135] <=  8'h67;        memory[47136] <=  8'h79;        memory[47137] <=  8'h76;        memory[47138] <=  8'h63;        memory[47139] <=  8'h68;        memory[47140] <=  8'h69;        memory[47141] <=  8'h6a;        memory[47142] <=  8'h33;        memory[47143] <=  8'h65;        memory[47144] <=  8'h67;        memory[47145] <=  8'h79;        memory[47146] <=  8'h72;        memory[47147] <=  8'h64;        memory[47148] <=  8'h62;        memory[47149] <=  8'h6e;        memory[47150] <=  8'h63;        memory[47151] <=  8'h7a;        memory[47152] <=  8'h6a;        memory[47153] <=  8'h6f;        memory[47154] <=  8'h66;        memory[47155] <=  8'h78;        memory[47156] <=  8'h6a;        memory[47157] <=  8'h69;        memory[47158] <=  8'h63;        memory[47159] <=  8'h68;        memory[47160] <=  8'h62;        memory[47161] <=  8'h6e;        memory[47162] <=  8'h6d;        memory[47163] <=  8'h63;        memory[47164] <=  8'h73;        memory[47165] <=  8'h6c;        memory[47166] <=  8'h6b;        memory[47167] <=  8'h6a;        memory[47168] <=  8'h69;        memory[47169] <=  8'h68;        memory[47170] <=  8'h76;        memory[47171] <=  8'h75;        memory[47172] <=  8'h69;        memory[47173] <=  8'h64;        memory[47174] <=  8'h68;        memory[47175] <=  8'h75;        memory[47176] <=  8'h67;        memory[47177] <=  8'h79;        memory[47178] <=  8'h62;        memory[47179] <=  8'h68;        memory[47180] <=  8'h65;        memory[47181] <=  8'h6a;        memory[47182] <=  8'h72;        memory[47183] <=  8'h6b;        memory[47184] <=  8'h6a;        memory[47185] <=  8'h6f;        memory[47186] <=  8'h64;        memory[47187] <=  8'h67;        memory[47188] <=  8'h69;        memory[47189] <=  8'h75;        memory[47190] <=  8'h69;        memory[47191] <=  8'h67;        memory[47192] <=  8'h76;        memory[47193] <=  8'h79;        memory[47194] <=  8'h75;        memory[47195] <=  8'h67;        memory[47196] <=  8'h78;        memory[47197] <=  8'h68;        memory[47198] <=  8'h63;        memory[47199] <=  8'h20;        memory[47200] <=  8'h20;        memory[47201] <=  8'h20;        memory[47202] <=  8'h78;        memory[47203] <=  8'h76;        memory[47204] <=  8'h20;        memory[47205] <=  8'h63;        memory[47206] <=  8'h78;        memory[47207] <=  8'h67;        memory[47208] <=  8'h79;        memory[47209] <=  8'h63;        memory[47210] <=  8'h75;        memory[47211] <=  8'h68;        memory[47212] <=  8'h6a;        memory[47213] <=  8'h6b;        memory[47214] <=  8'h61;        memory[47215] <=  8'h6c;        memory[47216] <=  8'h78;        memory[47217] <=  8'h76;        memory[47218] <=  8'h70;        memory[47219] <=  8'h6f;        memory[47220] <=  8'h69;        memory[47221] <=  8'h6a;        memory[47222] <=  8'h69;        memory[47223] <=  8'h68;        memory[47224] <=  8'h6a;        memory[47225] <=  8'h62;        memory[47226] <=  8'h77;        memory[47227] <=  8'h65;        memory[47228] <=  8'h6e;        memory[47229] <=  8'h61;        memory[47230] <=  8'h66;        memory[47231] <=  8'h6d;        memory[47232] <=  8'h64;        memory[47233] <=  8'h6b;        memory[47234] <=  8'h6d;        memory[47235] <=  8'h76;        memory[47236] <=  8'h6c;        memory[47237] <=  8'h63;        memory[47238] <=  8'h6f;        memory[47239] <=  8'h64;        memory[47240] <=  8'h69;        memory[47241] <=  8'h75;        memory[47242] <=  8'h68;        memory[47243] <=  8'h73;        memory[47244] <=  8'h66;        memory[47245] <=  8'h65;        memory[47246] <=  8'h62;        memory[47247] <=  8'h6e;        memory[47248] <=  8'h64;        memory[47249] <=  8'h73;        memory[47250] <=  8'h63;        memory[47251] <=  8'h6b;        memory[47252] <=  8'h20;        memory[47253] <=  8'h78;        memory[47254] <=  8'h6a;        memory[47255] <=  8'h78;        memory[47256] <=  8'h63;        memory[47257] <=  8'h73;        memory[47258] <=  8'h64;        memory[47259] <=  8'h66;        memory[47260] <=  8'h6b;        memory[47261] <=  8'h64;        memory[47262] <=  8'h6e;        memory[47263] <=  8'h6d;        memory[47264] <=  8'h64;        memory[47265] <=  8'h73;        memory[47266] <=  8'h63;        memory[47267] <=  8'h6b;        memory[47268] <=  8'h78;        memory[47269] <=  8'h6c;        memory[47270] <=  8'h6f;        memory[47271] <=  8'h66;        memory[47272] <=  8'h6a;        memory[47273] <=  8'h69;        memory[47274] <=  8'h61;        memory[47275] <=  8'h62;        memory[47276] <=  8'h6e;        memory[47277] <=  8'h20;        memory[47278] <=  8'h78;        memory[47279] <=  8'h6b;        memory[47280] <=  8'h6d;        memory[47281] <=  8'h20;        memory[47282] <=  8'h6f;        memory[47283] <=  8'h63;        memory[47284] <=  8'h76;        memory[47285] <=  8'h73;        memory[47286] <=  8'h64;        memory[47287] <=  8'h69;        memory[47288] <=  8'h66;        memory[47289] <=  8'h68;        memory[47290] <=  8'h65;        memory[47291] <=  8'h71;        memory[47292] <=  8'h6a;        memory[47293] <=  8'h77;        memory[47294] <=  8'h62;        memory[47295] <=  8'h65;        memory[47296] <=  8'h6e;        memory[47297] <=  8'h20;        memory[47298] <=  8'h6d;        memory[47299] <=  8'h64;        memory[47300] <=  8'h73;        memory[47301] <=  8'h6c;        memory[47302] <=  8'h76;        memory[47303] <=  8'h6b;        memory[47304] <=  8'h63;        memory[47305] <=  8'h78;        memory[47306] <=  8'h20;        memory[47307] <=  8'h6f;        memory[47308] <=  8'h78;        memory[47309] <=  8'h69;        memory[47310] <=  8'h63;        memory[47311] <=  8'h6a;        memory[47312] <=  8'h76;        memory[47313] <=  8'h64;        memory[47314] <=  8'h66;        memory[47315] <=  8'h65;        memory[47316] <=  8'h71;        memory[47317] <=  8'h6e;        memory[47318] <=  8'h20;        memory[47319] <=  8'h64;        memory[47320] <=  8'h6d;        memory[47321] <=  8'h73;        memory[47322] <=  8'h6c;        memory[47323] <=  8'h63;        memory[47324] <=  8'h78;        memory[47325] <=  8'h6b;        memory[47326] <=  8'h20;        memory[47327] <=  8'h6f;        memory[47328] <=  8'h78;        memory[47329] <=  8'h63;        memory[47330] <=  8'h76;        memory[47331] <=  8'h6a;        memory[47332] <=  8'h64;        memory[47333] <=  8'h62;        memory[47334] <=  8'h71;        memory[47335] <=  8'h77;        memory[47336] <=  8'h65;        memory[47337] <=  8'h6e;        memory[47338] <=  8'h6d;        memory[47339] <=  8'h64;        memory[47340] <=  8'h6c;        memory[47341] <=  8'h73;        memory[47342] <=  8'h2c;        memory[47343] <=  8'h76;        memory[47344] <=  8'h63;        memory[47345] <=  8'h78;        memory[47346] <=  8'h20;        memory[47347] <=  8'h63;        memory[47348] <=  8'h6f;        memory[47349] <=  8'h69;        memory[47350] <=  8'h76;        memory[47351] <=  8'h68;        memory[47352] <=  8'h73;        memory[47353] <=  8'h64;        memory[47354] <=  8'h62;        memory[47355] <=  8'h71;        memory[47356] <=  8'h77;        memory[47357] <=  8'h65;        memory[47358] <=  8'h6e;        memory[47359] <=  8'h64;        memory[47360] <=  8'h6b;        memory[47361] <=  8'h73;        memory[47362] <=  8'h76;        memory[47363] <=  8'h6f;        memory[47364] <=  8'h63;        memory[47365] <=  8'h20;        memory[47366] <=  8'h76;        memory[47367] <=  8'h69;        memory[47368] <=  8'h75;        memory[47369] <=  8'h69;        memory[47370] <=  8'h68;        memory[47371] <=  8'h63;        memory[47372] <=  8'h78;        memory[47373] <=  8'h69;        memory[47374] <=  8'h6f;        memory[47375] <=  8'h76;        memory[47376] <=  8'h73;        memory[47377] <=  8'h64;        memory[47378] <=  8'h61;        memory[47379] <=  8'h64;        memory[47380] <=  8'h6e;        memory[47381] <=  8'h77;        memory[47382] <=  8'h71;        memory[47383] <=  8'h6b;        memory[47384] <=  8'h6c;        memory[47385] <=  8'h73;        memory[47386] <=  8'h76;        memory[47387] <=  8'h6e;        memory[47388] <=  8'h62;        memory[47389] <=  8'h20;        memory[47390] <=  8'h64;        memory[47391] <=  8'h66;        memory[47392] <=  8'h6a;        memory[47393] <=  8'h6b;        memory[47394] <=  8'h71;        memory[47395] <=  8'h64;        memory[47396] <=  8'h77;        memory[47397] <=  8'h65;        memory[47398] <=  8'h6e;        memory[47399] <=  8'h62;        memory[47400] <=  8'h20;        memory[47401] <=  8'h64;        memory[47402] <=  8'h73;        memory[47403] <=  8'h76;        memory[47404] <=  8'h68;        memory[47405] <=  8'h64;        memory[47406] <=  8'h61;        memory[47407] <=  8'h71;        memory[47408] <=  8'h77;        memory[47409] <=  8'h6a;        memory[47410] <=  8'h65;        memory[47411] <=  8'h6e;        memory[47412] <=  8'h64;        memory[47413] <=  8'h20;        memory[47414] <=  8'h61;        memory[47415] <=  8'h63;        memory[47416] <=  8'h62;        memory[47417] <=  8'h68;        memory[47418] <=  8'h64;        memory[47419] <=  8'h61;        memory[47420] <=  8'h77;        memory[47421] <=  8'h71;        memory[47422] <=  8'h6e;        memory[47423] <=  8'h20;        memory[47424] <=  8'h62;        memory[47425] <=  8'h73;        memory[47426] <=  8'h76;        memory[47427] <=  8'h61;        memory[47428] <=  8'h67;        memory[47429] <=  8'h76;        memory[47430] <=  8'h68;        memory[47431] <=  8'h67;        memory[47432] <=  8'h61;        memory[47433] <=  8'h73;        memory[47434] <=  8'h6a;        memory[47435] <=  8'h6b;        memory[47436] <=  8'h63;        memory[47437] <=  8'h78;        memory[47438] <=  8'h76;        memory[47439] <=  8'h6e;        memory[47440] <=  8'h73;        memory[47441] <=  8'h64;        memory[47442] <=  8'h20;        memory[47443] <=  8'h66;        memory[47444] <=  8'h62;        memory[47445] <=  8'h64;        memory[47446] <=  8'h61;        memory[47447] <=  8'h73;        memory[47448] <=  8'h76;        memory[47449] <=  8'h67;        memory[47450] <=  8'h63;        memory[47451] <=  8'h79;        memory[47452] <=  8'h7a;        memory[47453] <=  8'h78;        memory[47454] <=  8'h79;        memory[47455] <=  8'h75;        memory[47456] <=  8'h20;        memory[47457] <=  8'h69;        memory[47458] <=  8'h6a;        memory[47459] <=  8'h64;        memory[47460] <=  8'h66;        memory[47461] <=  8'h6b;        memory[47462] <=  8'h61;        memory[47463] <=  8'h64;        memory[47464] <=  8'h63;        memory[47465] <=  8'h78;        memory[47466] <=  8'h68;        memory[47467] <=  8'h20;        memory[47468] <=  8'h67;        memory[47469] <=  8'h61;        memory[47470] <=  8'h68;        memory[47471] <=  8'h75;        memory[47472] <=  8'h64;        memory[47473] <=  8'h73;        memory[47474] <=  8'h69;        memory[47475] <=  8'h6a;        memory[47476] <=  8'h61;        memory[47477] <=  8'h6b;        memory[47478] <=  8'h63;        memory[47479] <=  8'h62;        memory[47480] <=  8'h61;        memory[47481] <=  8'h72;        memory[47482] <=  8'h73;        memory[47483] <=  8'h68;        memory[47484] <=  8'h64;        memory[47485] <=  8'h66;        memory[47486] <=  8'h67;        memory[47487] <=  8'h73;        memory[47488] <=  8'h68;        memory[47489] <=  8'h64;        memory[47490] <=  8'h66;        memory[47491] <=  8'h68;        memory[47492] <=  8'h64;        memory[47493] <=  8'h6a;        memory[47494] <=  8'h68;        memory[47495] <=  8'h62;        memory[47496] <=  8'h67;        memory[47497] <=  8'h63;        memory[47498] <=  8'h61;        memory[47499] <=  8'h66;        memory[47500] <=  8'h73;        memory[47501] <=  8'h79;        memory[47502] <=  8'h67;        memory[47503] <=  8'h6b;        memory[47504] <=  8'h75;        memory[47505] <=  8'h64;        memory[47506] <=  8'h68;        memory[47507] <=  8'h62;        memory[47508] <=  8'h77;        memory[47509] <=  8'h76;        memory[47510] <=  8'h67;        memory[47511] <=  8'h61;        memory[47512] <=  8'h66;        memory[47513] <=  8'h64;        memory[47514] <=  8'h74;        memory[47515] <=  8'h75;        memory[47516] <=  8'h66;        memory[47517] <=  8'h79;        memory[47518] <=  8'h67;        memory[47519] <=  8'h69;        memory[47520] <=  8'h75;        memory[47521] <=  8'h68;        memory[47522] <=  8'h6c;        memory[47523] <=  8'h6a;        memory[47524] <=  8'h62;        memory[47525] <=  8'h6b;        memory[47526] <=  8'h68;        memory[47527] <=  8'h76;        memory[47528] <=  8'h67;        memory[47529] <=  8'h63;        memory[47530] <=  8'h66;        memory[47531] <=  8'h78;        memory[47532] <=  8'h64;        memory[47533] <=  8'h74;        memory[47534] <=  8'h75;        memory[47535] <=  8'h79;        memory[47536] <=  8'h69;        memory[47537] <=  8'h75;        memory[47538] <=  8'h68;        memory[47539] <=  8'h6c;        memory[47540] <=  8'h6a;        memory[47541] <=  8'h6b;        memory[47542] <=  8'h67;        memory[47543] <=  8'h6a;        memory[47544] <=  8'h63;        memory[47545] <=  8'h66;        memory[47546] <=  8'h68;        memory[47547] <=  8'h64;        memory[47548] <=  8'h67;        memory[47549] <=  8'h72;        memory[47550] <=  8'h79;        memory[47551] <=  8'h74;        memory[47552] <=  8'h66;        memory[47553] <=  8'h75;        memory[47554] <=  8'h79;        memory[47555] <=  8'h69;        memory[47556] <=  8'h68;        memory[47557] <=  8'h6c;        memory[47558] <=  8'h62;        memory[47559] <=  8'h6d;        memory[47560] <=  8'h76;        memory[47561] <=  8'h6e;        memory[47562] <=  8'h63;        memory[47563] <=  8'h66;        memory[47564] <=  8'h68;        memory[47565] <=  8'h64;        memory[47566] <=  8'h74;        memory[47567] <=  8'h75;        memory[47568] <=  8'h67;        memory[47569] <=  8'h79;        memory[47570] <=  8'h69;        memory[47571] <=  8'h68;        memory[47572] <=  8'h75;        memory[47573] <=  8'h6a;        memory[47574] <=  8'h6c;        memory[47575] <=  8'h62;        memory[47576] <=  8'h6d;        memory[47577] <=  8'h76;        memory[47578] <=  8'h6e;        memory[47579] <=  8'h63;        memory[47580] <=  8'h66;        memory[47581] <=  8'h68;        memory[47582] <=  8'h67;        memory[47583] <=  8'h79;        memory[47584] <=  8'h68;        memory[47585] <=  8'h75;        memory[47586] <=  8'h6a;        memory[47587] <=  8'h6e;        memory[47588] <=  8'h2c;        memory[47589] <=  8'h62;        memory[47590] <=  8'h6e;        memory[47591] <=  8'h6d;        memory[47592] <=  8'h76;        memory[47593] <=  8'h6e;        memory[47594] <=  8'h63;        memory[47595] <=  8'h66;        memory[47596] <=  8'h68;        memory[47597] <=  8'h74;        memory[47598] <=  8'h79;        memory[47599] <=  8'h69;        memory[47600] <=  8'h75;        memory[47601] <=  8'h6c;        memory[47602] <=  8'h6a;        memory[47603] <=  8'h62;        memory[47604] <=  8'h6d;        memory[47605] <=  8'h76;        memory[47606] <=  8'h6e;        memory[47607] <=  8'h63;        memory[47608] <=  8'h66;        memory[47609] <=  8'h74;        memory[47610] <=  8'h75;        memory[47611] <=  8'h79;        memory[47612] <=  8'h69;        memory[47613] <=  8'h68;        memory[47614] <=  8'h6b;        memory[47615] <=  8'h62;        memory[47616] <=  8'h76;        memory[47617] <=  8'h63;        memory[47618] <=  8'h66;        memory[47619] <=  8'h67;        memory[47620] <=  8'h74;        memory[47621] <=  8'h75;        memory[47622] <=  8'h79;        memory[47623] <=  8'h69;        memory[47624] <=  8'h75;        memory[47625] <=  8'h68;        memory[47626] <=  8'h6a;        memory[47627] <=  8'h6b;        memory[47628] <=  8'h62;        memory[47629] <=  8'h76;        memory[47630] <=  8'h63;        memory[47631] <=  8'h66;        memory[47632] <=  8'h74;        memory[47633] <=  8'h75;        memory[47634] <=  8'h79;        memory[47635] <=  8'h69;        memory[47636] <=  8'h75;        memory[47637] <=  8'h6a;        memory[47638] <=  8'h6b;        memory[47639] <=  8'h6e;        memory[47640] <=  8'h62;        memory[47641] <=  8'h76;        memory[47642] <=  8'h67;        memory[47643] <=  8'h66;        memory[47644] <=  8'h74;        memory[47645] <=  8'h79;        memory[47646] <=  8'h75;        memory[47647] <=  8'h75;        memory[47648] <=  8'h69;        memory[47649] <=  8'h6a;        memory[47650] <=  8'h6b;        memory[47651] <=  8'h68;        memory[47652] <=  8'h62;        memory[47653] <=  8'h6a;        memory[47654] <=  8'h67;        memory[47655] <=  8'h68;        memory[47656] <=  8'h66;        memory[47657] <=  8'h79;        memory[47658] <=  8'h74;        memory[47659] <=  8'h79;        memory[47660] <=  8'h69;        memory[47661] <=  8'h75;        memory[47662] <=  8'h64;        memory[47663] <=  8'h6a;        memory[47664] <=  8'h6b;        memory[47665] <=  8'h68;        memory[47666] <=  8'h63;        memory[47667] <=  8'h7a;        memory[47668] <=  8'h67;        memory[47669] <=  8'h68;        memory[47670] <=  8'h74;        memory[47671] <=  8'h75;        memory[47672] <=  8'h79;        memory[47673] <=  8'h69;        memory[47674] <=  8'h61;        memory[47675] <=  8'h73;        memory[47676] <=  8'h75;        memory[47677] <=  8'h6a;        memory[47678] <=  8'h6b;        memory[47679] <=  8'h62;        memory[47680] <=  8'h6e;        memory[47681] <=  8'h61;        memory[47682] <=  8'h76;        memory[47683] <=  8'h63;        memory[47684] <=  8'h66;        memory[47685] <=  8'h68;        memory[47686] <=  8'h75;        memory[47687] <=  8'h61;        memory[47688] <=  8'h73;        memory[47689] <=  8'h79;        memory[47690] <=  8'h64;        memory[47691] <=  8'h75;        memory[47692] <=  8'h69;        memory[47693] <=  8'h6a;        memory[47694] <=  8'h61;        memory[47695] <=  8'h6b;        memory[47696] <=  8'h62;        memory[47697] <=  8'h63;        memory[47698] <=  8'h78;        memory[47699] <=  8'h68;        memory[47700] <=  8'h67;        memory[47701] <=  8'h79;        memory[47702] <=  8'h75;        memory[47703] <=  8'h7a;        memory[47704] <=  8'h63;        memory[47705] <=  8'h61;        memory[47706] <=  8'h73;        memory[47707] <=  8'h69;        memory[47708] <=  8'h75;        memory[47709] <=  8'h6f;        memory[47710] <=  8'h69;        memory[47711] <=  8'h6a;        memory[47712] <=  8'h61;        memory[47713] <=  8'h6c;        memory[47714] <=  8'h63;        memory[47715] <=  8'h78;        memory[47716] <=  8'h62;        memory[47717] <=  8'h63;        memory[47718] <=  8'h20;        memory[47719] <=  8'h6e;        memory[47720] <=  8'h76;        memory[47721] <=  8'h63;        memory[47722] <=  8'h61;        memory[47723] <=  8'h64;        memory[47724] <=  8'h73;        memory[47725] <=  8'h67;        memory[47726] <=  8'h79;        memory[47727] <=  8'h68;        memory[47728] <=  8'h75;        memory[47729] <=  8'h61;        memory[47730] <=  8'h6a;        memory[47731] <=  8'h6b;        memory[47732] <=  8'h78;        memory[47733] <=  8'h62;        memory[47734] <=  8'h20;        memory[47735] <=  8'h6e;        memory[47736] <=  8'h76;        memory[47737] <=  8'h63;        memory[47738] <=  8'h61;        memory[47739] <=  8'h73;        memory[47740] <=  8'h67;        memory[47741] <=  8'h68;        memory[47742] <=  8'h75;        memory[47743] <=  8'h6a;        memory[47744] <=  8'h6c;        memory[47745] <=  8'h6b;        memory[47746] <=  8'h63;        memory[47747] <=  8'h78;        memory[47748] <=  8'h20;        memory[47749] <=  8'h6a;        memory[47750] <=  8'h6b;        memory[47751] <=  8'h68;        memory[47752] <=  8'h61;        memory[47753] <=  8'h73;        memory[47754] <=  8'h76;        memory[47755] <=  8'h64;        memory[47756] <=  8'h6e;        memory[47757] <=  8'h20;        memory[47758] <=  8'h62;        memory[47759] <=  8'h6e;        memory[47760] <=  8'h6d;        memory[47761] <=  8'h6b;        memory[47762] <=  8'h77;        memory[47763] <=  8'h64;        memory[47764] <=  8'h6f;        memory[47765] <=  8'h77;        memory[47766] <=  8'h69;        memory[47767] <=  8'h6f;        memory[47768] <=  8'h75;        memory[47769] <=  8'h69;        memory[47770] <=  8'h68;        memory[47771] <=  8'h62;        memory[47772] <=  8'h6e;        memory[47773] <=  8'h6b;        memory[47774] <=  8'h77;        memory[47775] <=  8'h69;        memory[47776] <=  8'h6f;        memory[47777] <=  8'h75;        memory[47778] <=  8'h71;        memory[47779] <=  8'h69;        memory[47780] <=  8'h79;        memory[47781] <=  8'h67;        memory[47782] <=  8'h6a;        memory[47783] <=  8'h64;        memory[47784] <=  8'h61;        memory[47785] <=  8'h76;        memory[47786] <=  8'h62;        memory[47787] <=  8'h6e;        memory[47788] <=  8'h6b;        memory[47789] <=  8'h6f;        memory[47790] <=  8'h70;        memory[47791] <=  8'h64;        memory[47792] <=  8'h76;        memory[47793] <=  8'h69;        memory[47794] <=  8'h6f;        memory[47795] <=  8'h75;        memory[47796] <=  8'h69;        memory[47797] <=  8'h48;        memory[47798] <=  8'h42;        memory[47799] <=  8'h6b;        memory[47800] <=  8'h64;        memory[47801] <=  8'h6e;        memory[47802] <=  8'h6c;        memory[47803] <=  8'h71;        memory[47804] <=  8'h6b;        memory[47805] <=  8'h6d;        memory[47806] <=  8'h6a;        memory[47807] <=  8'h70;        memory[47808] <=  8'h69;        memory[47809] <=  8'h6f;        memory[47810] <=  8'h68;        memory[47811] <=  8'h65;        memory[47812] <=  8'h66;        memory[47813] <=  8'h75;        memory[47814] <=  8'h67;        memory[47815] <=  8'h69;        memory[47816] <=  8'h73;        memory[47817] <=  8'h61;        memory[47818] <=  8'h62;        memory[47819] <=  8'h64;        memory[47820] <=  8'h6b;        memory[47821] <=  8'h6a;        memory[47822] <=  8'h6b;        memory[47823] <=  8'h6c;        memory[47824] <=  8'h6a;        memory[47825] <=  8'h69;        memory[47826] <=  8'h73;        memory[47827] <=  8'h6f;        memory[47828] <=  8'h71;        memory[47829] <=  8'h68;        memory[47830] <=  8'h77;        memory[47831] <=  8'h67;        memory[47832] <=  8'h69;        memory[47833] <=  8'h79;        memory[47834] <=  8'h6a;        memory[47835] <=  8'h64;        memory[47836] <=  8'h76;        memory[47837] <=  8'h62;        memory[47838] <=  8'h6e;        memory[47839] <=  8'h61;        memory[47840] <=  8'h73;        memory[47841] <=  8'h66;        memory[47842] <=  8'h6c;        memory[47843] <=  8'h6b;        memory[47844] <=  8'h64;        memory[47845] <=  8'h6a;        memory[47846] <=  8'h68;        memory[47847] <=  8'h63;        memory[47848] <=  8'h67;        memory[47849] <=  8'h6a;        memory[47850] <=  8'h76;        memory[47851] <=  8'h73;        memory[47852] <=  8'h64;        memory[47853] <=  8'h62;        memory[47854] <=  8'h62;        memory[47855] <=  8'h61;        memory[47856] <=  8'h72;        memory[47857] <=  8'h62;        memory[47858] <=  8'h62;        memory[47859] <=  8'h73;        memory[47860] <=  8'h62;        memory[47861] <=  8'h67;        memory[47862] <=  8'h73;        memory[47863] <=  8'h66;        memory[47864] <=  8'h67;        memory[47865] <=  8'h61;        memory[47866] <=  8'h68;        memory[47867] <=  8'h66;        memory[47868] <=  8'h73;        memory[47869] <=  8'h68;        memory[47870] <=  8'h61;        memory[47871] <=  8'h66;        memory[47872] <=  8'h73;        memory[47873] <=  8'h66;        memory[47874] <=  8'h68;        memory[47875] <=  8'h61;        memory[47876] <=  8'h69;        memory[47877] <=  8'h64;        memory[47878] <=  8'h75;        memory[47879] <=  8'h67;        memory[47880] <=  8'h64;        memory[47881] <=  8'h77;        memory[47882] <=  8'h62;        memory[47883] <=  8'h61;        memory[47884] <=  8'h62;        memory[47885] <=  8'h72;        memory[47886] <=  8'h62;        memory[47887] <=  8'h61;        memory[47888] <=  8'h62;        memory[47889] <=  8'h62;        memory[47890] <=  8'h74;        memory[47891] <=  8'h62;        memory[47892] <=  8'h62;        memory[47893] <=  8'h62;        memory[47894] <=  8'h62;        memory[47895] <=  8'h62;        memory[47896] <=  8'h62;        memory[47897] <=  8'h62;        memory[47898] <=  8'h62;        memory[47899] <=  8'h61;        memory[47900] <=  8'h62;        memory[47901] <=  8'h62;        memory[47902] <=  8'h72;        memory[47903] <=  8'h74;        memory[47904] <=  8'h62;        memory[47905] <=  8'h62;        memory[47906] <=  8'h61;        memory[47907] <=  8'h62;        memory[47908] <=  8'h72;        memory[47909] <=  8'h62;        memory[47910] <=  8'h74;        memory[47911] <=  8'h62;        memory[47912] <=  8'h62;        memory[47913] <=  8'h62;        memory[47914] <=  8'h63;        memory[47915] <=  8'h61;        memory[47916] <=  8'h72;        memory[47917] <=  8'h74;        memory[47918] <=  8'h73;        memory[47919] <=  8'h62;        memory[47920] <=  8'h61;        memory[47921] <=  8'h72;        memory[47922] <=  8'h74;        memory[47923] <=  8'h74;        memory[47924] <=  8'h62;        memory[47925] <=  8'h61;        memory[47926] <=  8'h72;        memory[47927] <=  8'h74;        memory[47928] <=  8'h78;        memory[47929] <=  8'h61;        memory[47930] <=  8'h74;        memory[47931] <=  8'h6b;        memory[47932] <=  8'h73;        memory[47933] <=  8'h68;        memory[47934] <=  8'h63;        memory[47935] <=  8'h66;        memory[47936] <=  8'h69;        memory[47937] <=  8'h77;        memory[47938] <=  8'h68;        memory[47939] <=  8'h61;        memory[47940] <=  8'h74;        memory[47941] <=  8'h61;        memory[47942] <=  8'h6e;        memory[47943] <=  8'h61;        memory[47944] <=  8'h62;        memory[47945] <=  8'h61;        memory[47946] <=  8'h63;        memory[47947] <=  8'h61;        memory[47948] <=  8'h74;        memory[47949] <=  8'h61;        memory[47950] <=  8'h62;        memory[47951] <=  8'h61;        memory[47952] <=  8'h72;        memory[47953] <=  8'h63;        memory[47954] <=  8'h61;        memory[47955] <=  8'h68;        memory[47956] <=  8'h64;        memory[47957] <=  8'h75;        memory[47958] <=  8'h63;        memory[47959] <=  8'h74;        memory[47960] <=  8'h61;        memory[47961] <=  8'h64;        memory[47962] <=  8'h61;        memory[47963] <=  8'h61;        memory[47964] <=  8'h63;        memory[47965] <=  8'h61;        memory[47966] <=  8'h72;        memory[47967] <=  8'h63;        memory[47968] <=  8'h74;        memory[47969] <=  8'h72;        memory[47970] <=  8'h63;        memory[47971] <=  8'h61;        memory[47972] <=  8'h74;        memory[47973] <=  8'h72;        memory[47974] <=  8'h63;        memory[47975] <=  8'h61;        memory[47976] <=  8'h74;        memory[47977] <=  8'h63;        memory[47978] <=  8'h62;        memory[47979] <=  8'h61;        memory[47980] <=  8'h74;        memory[47981] <=  8'h62;        memory[47982] <=  8'h72;        memory[47983] <=  8'h63;        memory[47984] <=  8'h61;        memory[47985] <=  8'h74;        memory[47986] <=  8'h72;        memory[47987] <=  8'h6e;        memory[47988] <=  8'h62;        memory[47989] <=  8'h61;        memory[47990] <=  8'h63;        memory[47991] <=  8'h61;        memory[47992] <=  8'h74;        memory[47993] <=  8'h79;        memory[47994] <=  8'h73;        memory[47995] <=  8'h6e;        memory[47996] <=  8'h63;        memory[47997] <=  8'h74;        memory[47998] <=  8'h61;        memory[47999] <=  8'h6e;        memory[48000] <=  8'h62;        memory[48001] <=  8'h61;        memory[48002] <=  8'h63;        memory[48003] <=  8'h72;        memory[48004] <=  8'h6e;        memory[48005] <=  8'h74;        memory[48006] <=  8'h61;        memory[48007] <=  8'h62;        memory[48008] <=  8'h74;        memory[48009] <=  8'h6e;        memory[48010] <=  8'h61;        memory[48011] <=  8'h72;        memory[48012] <=  8'h62;        memory[48013] <=  8'h78;        memory[48014] <=  8'h74;        memory[48015] <=  8'h61;        memory[48016] <=  8'h72;        memory[48017] <=  8'h62;        memory[48018] <=  8'h61;        memory[48019] <=  8'h72;        memory[48020] <=  8'h74;        memory[48021] <=  8'h74;        memory[48022] <=  8'h62;        memory[48023] <=  8'h61;        memory[48024] <=  8'h72;        memory[48025] <=  8'h74;        memory[48026] <=  8'h78;        memory[48027] <=  8'h61;        memory[48028] <=  8'h74;        memory[48029] <=  8'h6b;        memory[48030] <=  8'h73;        memory[48031] <=  8'h68;        memory[48032] <=  8'h63;        memory[48033] <=  8'h66;        memory[48034] <=  8'h69;        memory[48035] <=  8'h77;        memory[48036] <=  8'h68;        memory[48037] <=  8'h61;        memory[48038] <=  8'h74;        memory[48039] <=  8'h61;        memory[48040] <=  8'h6e;        memory[48041] <=  8'h61;        memory[48042] <=  8'h62;        memory[48043] <=  8'h61;        memory[48044] <=  8'h63;        memory[48045] <=  8'h61;        memory[48046] <=  8'h74;        memory[48047] <=  8'h61;        memory[48048] <=  8'h62;        memory[48049] <=  8'h61;        memory[48050] <=  8'h72;        memory[48051] <=  8'h63;        memory[48052] <=  8'h61;        memory[48053] <=  8'h68;        memory[48054] <=  8'h64;        memory[48055] <=  8'h75;        memory[48056] <=  8'h63;        memory[48057] <=  8'h74;        memory[48058] <=  8'h61;        memory[48059] <=  8'h64;        memory[48060] <=  8'h61;        memory[48061] <=  8'h61;        memory[48062] <=  8'h63;        memory[48063] <=  8'h61;        memory[48064] <=  8'h72;        memory[48065] <=  8'h63;        memory[48066] <=  8'h74;        memory[48067] <=  8'h72;        memory[48068] <=  8'h63;        memory[48069] <=  8'h61;        memory[48070] <=  8'h74;        memory[48071] <=  8'h72;        memory[48072] <=  8'h63;        memory[48073] <=  8'h61;        memory[48074] <=  8'h74;        memory[48075] <=  8'h63;        memory[48076] <=  8'h62;        memory[48077] <=  8'h61;        memory[48078] <=  8'h74;        memory[48079] <=  8'h62;        memory[48080] <=  8'h72;        memory[48081] <=  8'h63;        memory[48082] <=  8'h61;        memory[48083] <=  8'h74;        memory[48084] <=  8'h72;        memory[48085] <=  8'h6e;        memory[48086] <=  8'h62;        memory[48087] <=  8'h61;        memory[48088] <=  8'h63;        memory[48089] <=  8'h61;        memory[48090] <=  8'h74;        memory[48091] <=  8'h79;        memory[48092] <=  8'h73;        memory[48093] <=  8'h6e;        memory[48094] <=  8'h63;        memory[48095] <=  8'h74;        memory[48096] <=  8'h61;        memory[48097] <=  8'h6e;        memory[48098] <=  8'h62;        memory[48099] <=  8'h61;        memory[48100] <=  8'h63;        memory[48101] <=  8'h72;        memory[48102] <=  8'h6e;        memory[48103] <=  8'h74;        memory[48104] <=  8'h61;        memory[48105] <=  8'h62;        memory[48106] <=  8'h74;        memory[48107] <=  8'h6e;        memory[48108] <=  8'h61;        memory[48109] <=  8'h72;        memory[48110] <=  8'h62;        memory[48111] <=  8'h78;        memory[48112] <=  8'h74;        memory[48113] <=  8'h61;        memory[48114] <=  8'h72;        memory[48115] <=  8'h62;        memory[48116] <=  8'h61;        memory[48117] <=  8'h72;        memory[48118] <=  8'h74;        memory[48119] <=  8'h74;        memory[48120] <=  8'h62;        memory[48121] <=  8'h61;        memory[48122] <=  8'h72;        memory[48123] <=  8'h74;        memory[48124] <=  8'h78;        memory[48125] <=  8'h61;        memory[48126] <=  8'h74;        memory[48127] <=  8'h6b;        memory[48128] <=  8'h73;        memory[48129] <=  8'h68;        memory[48130] <=  8'h63;        memory[48131] <=  8'h66;        memory[48132] <=  8'h69;        memory[48133] <=  8'h77;        memory[48134] <=  8'h68;        memory[48135] <=  8'h61;        memory[48136] <=  8'h74;        memory[48137] <=  8'h61;        memory[48138] <=  8'h6e;        memory[48139] <=  8'h61;        memory[48140] <=  8'h62;        memory[48141] <=  8'h61;        memory[48142] <=  8'h63;        memory[48143] <=  8'h61;        memory[48144] <=  8'h74;        memory[48145] <=  8'h61;        memory[48146] <=  8'h62;        memory[48147] <=  8'h61;        memory[48148] <=  8'h72;        memory[48149] <=  8'h63;        memory[48150] <=  8'h61;        memory[48151] <=  8'h68;        memory[48152] <=  8'h64;        memory[48153] <=  8'h75;        memory[48154] <=  8'h63;        memory[48155] <=  8'h74;        memory[48156] <=  8'h61;        memory[48157] <=  8'h64;        memory[48158] <=  8'h61;        memory[48159] <=  8'h61;        memory[48160] <=  8'h63;        memory[48161] <=  8'h61;        memory[48162] <=  8'h72;        memory[48163] <=  8'h63;        memory[48164] <=  8'h74;        memory[48165] <=  8'h72;        memory[48166] <=  8'h63;        memory[48167] <=  8'h61;        memory[48168] <=  8'h74;        memory[48169] <=  8'h72;        memory[48170] <=  8'h63;        memory[48171] <=  8'h61;        memory[48172] <=  8'h74;        memory[48173] <=  8'h63;        memory[48174] <=  8'h62;        memory[48175] <=  8'h61;        memory[48176] <=  8'h74;        memory[48177] <=  8'h62;        memory[48178] <=  8'h72;        memory[48179] <=  8'h63;        memory[48180] <=  8'h61;        memory[48181] <=  8'h74;        memory[48182] <=  8'h72;        memory[48183] <=  8'h6e;        memory[48184] <=  8'h62;        memory[48185] <=  8'h61;        memory[48186] <=  8'h63;        memory[48187] <=  8'h61;        memory[48188] <=  8'h74;        memory[48189] <=  8'h79;        memory[48190] <=  8'h73;        memory[48191] <=  8'h6e;        memory[48192] <=  8'h63;        memory[48193] <=  8'h74;        memory[48194] <=  8'h61;        memory[48195] <=  8'h6e;        memory[48196] <=  8'h62;        memory[48197] <=  8'h61;        memory[48198] <=  8'h63;        memory[48199] <=  8'h72;        memory[48200] <=  8'h6e;        memory[48201] <=  8'h74;        memory[48202] <=  8'h61;        memory[48203] <=  8'h62;        memory[48204] <=  8'h74;        memory[48205] <=  8'h6e;        memory[48206] <=  8'h61;        memory[48207] <=  8'h72;        memory[48208] <=  8'h62;        memory[48209] <=  8'h78;        memory[48210] <=  8'h74;        memory[48211] <=  8'h61;        memory[48212] <=  8'h72;        memory[48213] <=  8'h5d;        memory[48214] <=  8'h5d;        memory[48215] <=  8'h65;        memory[48216] <=  8'h66;        memory[48217] <=  8'h77;        memory[48218] <=  8'h65;        memory[48219] <=  8'h5d;        memory[48220] <=  8'h65;        memory[48221] <=  8'h67;        memory[48222] <=  8'h73;        memory[48223] <=  8'h67;        memory[48224] <=  8'h66;        memory[48225] <=  8'h62;        memory[48226] <=  8'h61;        memory[48227] <=  8'h72;        memory[48228] <=  8'h74;        memory[48229] <=  8'h74;        memory[48230] <=  8'h62;        memory[48231] <=  8'h61;        memory[48232] <=  8'h72;        memory[48233] <=  8'h74;        memory[48234] <=  8'h78;        memory[48235] <=  8'h61;        memory[48236] <=  8'h74;        memory[48237] <=  8'h6b;        memory[48238] <=  8'h73;        memory[48239] <=  8'h68;        memory[48240] <=  8'h63;        memory[48241] <=  8'h66;        memory[48242] <=  8'h69;        memory[48243] <=  8'h77;        memory[48244] <=  8'h68;        memory[48245] <=  8'h61;        memory[48246] <=  8'h74;        memory[48247] <=  8'h61;        memory[48248] <=  8'h6e;        memory[48249] <=  8'h61;        memory[48250] <=  8'h62;        memory[48251] <=  8'h61;        memory[48252] <=  8'h63;        memory[48253] <=  8'h61;        memory[48254] <=  8'h74;        memory[48255] <=  8'h61;        memory[48256] <=  8'h62;        memory[48257] <=  8'h61;        memory[48258] <=  8'h72;        memory[48259] <=  8'h63;        memory[48260] <=  8'h61;        memory[48261] <=  8'h68;        memory[48262] <=  8'h64;        memory[48263] <=  8'h75;        memory[48264] <=  8'h63;        memory[48265] <=  8'h74;        memory[48266] <=  8'h61;        memory[48267] <=  8'h64;        memory[48268] <=  8'h61;        memory[48269] <=  8'h61;        memory[48270] <=  8'h63;        memory[48271] <=  8'h61;        memory[48272] <=  8'h72;        memory[48273] <=  8'h63;        memory[48274] <=  8'h74;        memory[48275] <=  8'h72;        memory[48276] <=  8'h63;        memory[48277] <=  8'h61;        memory[48278] <=  8'h74;        memory[48279] <=  8'h72;        memory[48280] <=  8'h63;        memory[48281] <=  8'h61;        memory[48282] <=  8'h74;        memory[48283] <=  8'h63;        memory[48284] <=  8'h62;        memory[48285] <=  8'h61;        memory[48286] <=  8'h74;        memory[48287] <=  8'h62;        memory[48288] <=  8'h72;        memory[48289] <=  8'h63;        memory[48290] <=  8'h61;        memory[48291] <=  8'h74;        memory[48292] <=  8'h72;        memory[48293] <=  8'h6e;        memory[48294] <=  8'h62;        memory[48295] <=  8'h61;        memory[48296] <=  8'h63;        memory[48297] <=  8'h61;        memory[48298] <=  8'h74;        memory[48299] <=  8'h79;        memory[48300] <=  8'h73;        memory[48301] <=  8'h6e;        memory[48302] <=  8'h63;        memory[48303] <=  8'h74;        memory[48304] <=  8'h61;        memory[48305] <=  8'h6e;        memory[48306] <=  8'h62;        memory[48307] <=  8'h61;        memory[48308] <=  8'h63;        memory[48309] <=  8'h72;        memory[48310] <=  8'h6e;        memory[48311] <=  8'h74;        memory[48312] <=  8'h61;        memory[48313] <=  8'h62;        memory[48314] <=  8'h74;        memory[48315] <=  8'h6e;        memory[48316] <=  8'h61;        memory[48317] <=  8'h72;        memory[48318] <=  8'h62;        memory[48319] <=  8'h78;        memory[48320] <=  8'h74;        memory[48321] <=  8'h61;        memory[48322] <=  8'h72;        memory[48323] <=  8'h62;        memory[48324] <=  8'h61;        memory[48325] <=  8'h72;        memory[48326] <=  8'h74;        memory[48327] <=  8'h74;        memory[48328] <=  8'h62;        memory[48329] <=  8'h61;        memory[48330] <=  8'h72;        memory[48331] <=  8'h74;        memory[48332] <=  8'h78;        memory[48333] <=  8'h61;        memory[48334] <=  8'h74;        memory[48335] <=  8'h6b;        memory[48336] <=  8'h73;        memory[48337] <=  8'h68;        memory[48338] <=  8'h63;        memory[48339] <=  8'h66;        memory[48340] <=  8'h69;        memory[48341] <=  8'h77;        memory[48342] <=  8'h68;        memory[48343] <=  8'h61;        memory[48344] <=  8'h74;        memory[48345] <=  8'h61;        memory[48346] <=  8'h6e;        memory[48347] <=  8'h61;        memory[48348] <=  8'h62;        memory[48349] <=  8'h61;        memory[48350] <=  8'h63;        memory[48351] <=  8'h61;        memory[48352] <=  8'h74;        memory[48353] <=  8'h61;        memory[48354] <=  8'h62;        memory[48355] <=  8'h61;        memory[48356] <=  8'h72;        memory[48357] <=  8'h63;        memory[48358] <=  8'h61;        memory[48359] <=  8'h68;        memory[48360] <=  8'h64;        memory[48361] <=  8'h75;        memory[48362] <=  8'h63;        memory[48363] <=  8'h74;        memory[48364] <=  8'h61;        memory[48365] <=  8'h64;        memory[48366] <=  8'h61;        memory[48367] <=  8'h61;        memory[48368] <=  8'h63;        memory[48369] <=  8'h61;        memory[48370] <=  8'h72;        memory[48371] <=  8'h63;        memory[48372] <=  8'h74;        memory[48373] <=  8'h72;        memory[48374] <=  8'h63;        memory[48375] <=  8'h61;        memory[48376] <=  8'h74;        memory[48377] <=  8'h72;        memory[48378] <=  8'h63;        memory[48379] <=  8'h61;        memory[48380] <=  8'h74;        memory[48381] <=  8'h63;        memory[48382] <=  8'h62;        memory[48383] <=  8'h61;        memory[48384] <=  8'h74;        memory[48385] <=  8'h62;        memory[48386] <=  8'h72;        memory[48387] <=  8'h63;        memory[48388] <=  8'h61;        memory[48389] <=  8'h74;        memory[48390] <=  8'h72;        memory[48391] <=  8'h6e;        memory[48392] <=  8'h62;        memory[48393] <=  8'h61;        memory[48394] <=  8'h63;        memory[48395] <=  8'h61;        memory[48396] <=  8'h74;        memory[48397] <=  8'h79;        memory[48398] <=  8'h73;        memory[48399] <=  8'h6e;        memory[48400] <=  8'h63;        memory[48401] <=  8'h74;        memory[48402] <=  8'h61;        memory[48403] <=  8'h6e;        memory[48404] <=  8'h62;        memory[48405] <=  8'h61;        memory[48406] <=  8'h63;        memory[48407] <=  8'h72;        memory[48408] <=  8'h6e;        memory[48409] <=  8'h74;        memory[48410] <=  8'h61;        memory[48411] <=  8'h62;        memory[48412] <=  8'h74;        memory[48413] <=  8'h6e;        memory[48414] <=  8'h61;        memory[48415] <=  8'h72;        memory[48416] <=  8'h62;        memory[48417] <=  8'h78;        memory[48418] <=  8'h74;        memory[48419] <=  8'h61;        memory[48420] <=  8'h72;        memory[48421] <=  8'h64;        memory[48422] <=  8'h66;        memory[48423] <=  8'h73;        memory[48424] <=  8'h67;        memory[48425] <=  8'h76;        memory[48426] <=  8'h68;        memory[48427] <=  8'h62;        memory[48428] <=  8'h6b;        memory[48429] <=  8'h6a;        memory[48430] <=  8'h6e;        memory[48431] <=  8'h6d;        memory[48432] <=  8'h62;        memory[48433] <=  8'h76;        memory[48434] <=  8'h78;        memory[48435] <=  8'h63;        memory[48436] <=  8'h73;        memory[48437] <=  8'h66;        memory[48438] <=  8'h72;        memory[48439] <=  8'h74;        memory[48440] <=  8'h79;        memory[48441] <=  8'h75;        memory[48442] <=  8'h6a;        memory[48443] <=  8'h6e;        memory[48444] <=  8'h62;        memory[48445] <=  8'h76;        memory[48446] <=  8'h63;        memory[48447] <=  8'h64;        memory[48448] <=  8'h74;        memory[48449] <=  8'h79;        memory[48450] <=  8'h75;        memory[48451] <=  8'h69;        memory[48452] <=  8'h6b;        memory[48453] <=  8'h6d;        memory[48454] <=  8'h6e;        memory[48455] <=  8'h62;        memory[48456] <=  8'h76;        memory[48457] <=  8'h63;        memory[48458] <=  8'h78;        memory[48459] <=  8'h73;        memory[48460] <=  8'h64;        memory[48461] <=  8'h72;        memory[48462] <=  8'h74;        memory[48463] <=  8'h79;        memory[48464] <=  8'h75;        memory[48465] <=  8'h69;        memory[48466] <=  8'h6b;        memory[48467] <=  8'h6d;        memory[48468] <=  8'h6e;        memory[48469] <=  8'h62;        memory[48470] <=  8'h76;        memory[48471] <=  8'h63;        memory[48472] <=  8'h73;        memory[48473] <=  8'h77;        memory[48474] <=  8'h33;        memory[48475] <=  8'h34;        memory[48476] <=  8'h35;        memory[48477] <=  8'h36;        memory[48478] <=  8'h37;        memory[48479] <=  8'h38;        memory[48480] <=  8'h69;        memory[48481] <=  8'h6b;        memory[48482] <=  8'h6d;        memory[48483] <=  8'h6e;        memory[48484] <=  8'h62;        memory[48485] <=  8'h76;        memory[48486] <=  8'h63;        memory[48487] <=  8'h64;        memory[48488] <=  8'h65;        memory[48489] <=  8'h72;        memory[48490] <=  8'h36;        memory[48491] <=  8'h37;        memory[48492] <=  8'h38;        memory[48493] <=  8'h69;        memory[48494] <=  8'h6f;        memory[48495] <=  8'h6b;        memory[48496] <=  8'h6a;        memory[48497] <=  8'h6e;        memory[48498] <=  8'h62;        memory[48499] <=  8'h76;        memory[48500] <=  8'h63;        memory[48501] <=  8'h64;        memory[48502] <=  8'h72;        memory[48503] <=  8'h74;        memory[48504] <=  8'h79;        memory[48505] <=  8'h75;        memory[48506] <=  8'h73;        memory[48507] <=  8'h6a;        memory[48508] <=  8'h63;        memory[48509] <=  8'h6e;        memory[48510] <=  8'h62;        memory[48511] <=  8'h64;        memory[48512] <=  8'h66;        memory[48513] <=  8'h73;        memory[48514] <=  8'h74;        memory[48515] <=  8'h79;        memory[48516] <=  8'h75;        memory[48517] <=  8'h61;        memory[48518] <=  8'h69;        memory[48519] <=  8'h6b;        memory[48520] <=  8'h78;        memory[48521] <=  8'h6d;        memory[48522] <=  8'h6e;        memory[48523] <=  8'h73;        memory[48524] <=  8'h6a;        memory[48525] <=  8'h6f;        memory[48526] <=  8'h64;        memory[48527] <=  8'h6c;        memory[48528] <=  8'h63;        memory[48529] <=  8'h78;        memory[48530] <=  8'h62;        memory[48531] <=  8'h61;        memory[48532] <=  8'h72;        memory[48533] <=  8'h74;        memory[48534] <=  8'h78;        memory[48535] <=  8'h61;        memory[48536] <=  8'h74;        memory[48537] <=  8'h6b;        memory[48538] <=  8'h73;        memory[48539] <=  8'h68;        memory[48540] <=  8'h63;        memory[48541] <=  8'h66;        memory[48542] <=  8'h69;        memory[48543] <=  8'h77;        memory[48544] <=  8'h68;        memory[48545] <=  8'h61;        memory[48546] <=  8'h74;        memory[48547] <=  8'h61;        memory[48548] <=  8'h6e;        memory[48549] <=  8'h61;        memory[48550] <=  8'h62;        memory[48551] <=  8'h61;        memory[48552] <=  8'h63;        memory[48553] <=  8'h61;        memory[48554] <=  8'h74;        memory[48555] <=  8'h61;        memory[48556] <=  8'h62;        memory[48557] <=  8'h61;        memory[48558] <=  8'h72;        memory[48559] <=  8'h63;        memory[48560] <=  8'h61;        memory[48561] <=  8'h68;        memory[48562] <=  8'h64;        memory[48563] <=  8'h75;        memory[48564] <=  8'h63;        memory[48565] <=  8'h74;        memory[48566] <=  8'h61;        memory[48567] <=  8'h64;        memory[48568] <=  8'h61;        memory[48569] <=  8'h61;        memory[48570] <=  8'h63;        memory[48571] <=  8'h61;        memory[48572] <=  8'h72;        memory[48573] <=  8'h62;        memory[48574] <=  8'h61;        memory[48575] <=  8'h72;        memory[48576] <=  8'h74;        memory[48577] <=  8'h78;        memory[48578] <=  8'h61;        memory[48579] <=  8'h74;        memory[48580] <=  8'h6b;        memory[48581] <=  8'h73;        memory[48582] <=  8'h68;        memory[48583] <=  8'h63;        memory[48584] <=  8'h66;        memory[48585] <=  8'h69;        memory[48586] <=  8'h77;        memory[48587] <=  8'h68;        memory[48588] <=  8'h61;        memory[48589] <=  8'h74;        memory[48590] <=  8'h61;        memory[48591] <=  8'h6e;        memory[48592] <=  8'h61;        memory[48593] <=  8'h62;        memory[48594] <=  8'h61;        memory[48595] <=  8'h63;        memory[48596] <=  8'h61;        memory[48597] <=  8'h74;        memory[48598] <=  8'h61;        memory[48599] <=  8'h62;        memory[48600] <=  8'h61;        memory[48601] <=  8'h72;        memory[48602] <=  8'h63;        memory[48603] <=  8'h61;        memory[48604] <=  8'h68;        memory[48605] <=  8'h64;        memory[48606] <=  8'h75;        memory[48607] <=  8'h63;        memory[48608] <=  8'h74;        memory[48609] <=  8'h61;        memory[48610] <=  8'h64;        memory[48611] <=  8'h61;        memory[48612] <=  8'h61;        memory[48613] <=  8'h63;        memory[48614] <=  8'h61;        memory[48615] <=  8'h72;        memory[48616] <=  8'h62;        memory[48617] <=  8'h61;        memory[48618] <=  8'h72;        memory[48619] <=  8'h74;        memory[48620] <=  8'h78;        memory[48621] <=  8'h61;        memory[48622] <=  8'h74;        memory[48623] <=  8'h6b;        memory[48624] <=  8'h73;        memory[48625] <=  8'h68;        memory[48626] <=  8'h63;        memory[48627] <=  8'h66;        memory[48628] <=  8'h69;        memory[48629] <=  8'h77;        memory[48630] <=  8'h68;        memory[48631] <=  8'h61;        memory[48632] <=  8'h74;        memory[48633] <=  8'h61;        memory[48634] <=  8'h6e;        memory[48635] <=  8'h61;        memory[48636] <=  8'h62;        memory[48637] <=  8'h61;        memory[48638] <=  8'h63;        memory[48639] <=  8'h61;        memory[48640] <=  8'h74;        memory[48641] <=  8'h61;        memory[48642] <=  8'h62;        memory[48643] <=  8'h61;        memory[48644] <=  8'h72;        memory[48645] <=  8'h63;        memory[48646] <=  8'h61;        memory[48647] <=  8'h68;        memory[48648] <=  8'h64;        memory[48649] <=  8'h75;        memory[48650] <=  8'h63;        memory[48651] <=  8'h74;        memory[48652] <=  8'h61;        memory[48653] <=  8'h64;        memory[48654] <=  8'h61;        memory[48655] <=  8'h61;        memory[48656] <=  8'h63;        memory[48657] <=  8'h61;        memory[48658] <=  8'h72;        memory[48659] <=  8'h62;        memory[48660] <=  8'h61;        memory[48661] <=  8'h72;        memory[48662] <=  8'h74;        memory[48663] <=  8'h78;        memory[48664] <=  8'h61;        memory[48665] <=  8'h74;        memory[48666] <=  8'h6b;        memory[48667] <=  8'h73;        memory[48668] <=  8'h68;        memory[48669] <=  8'h63;        memory[48670] <=  8'h66;        memory[48671] <=  8'h69;        memory[48672] <=  8'h77;        memory[48673] <=  8'h68;        memory[48674] <=  8'h61;        memory[48675] <=  8'h74;        memory[48676] <=  8'h61;        memory[48677] <=  8'h6e;        memory[48678] <=  8'h61;        memory[48679] <=  8'h62;        memory[48680] <=  8'h61;        memory[48681] <=  8'h63;        memory[48682] <=  8'h61;        memory[48683] <=  8'h74;        memory[48684] <=  8'h61;        memory[48685] <=  8'h62;        memory[48686] <=  8'h61;        memory[48687] <=  8'h72;        memory[48688] <=  8'h63;        memory[48689] <=  8'h61;        memory[48690] <=  8'h68;        memory[48691] <=  8'h64;        memory[48692] <=  8'h75;        memory[48693] <=  8'h63;        memory[48694] <=  8'h74;        memory[48695] <=  8'h61;        memory[48696] <=  8'h64;        memory[48697] <=  8'h61;        memory[48698] <=  8'h61;        memory[48699] <=  8'h63;        memory[48700] <=  8'h61;        memory[48701] <=  8'h72;        memory[48702] <=  8'h62;        memory[48703] <=  8'h61;        memory[48704] <=  8'h72;        memory[48705] <=  8'h74;        memory[48706] <=  8'h78;        memory[48707] <=  8'h61;        memory[48708] <=  8'h74;        memory[48709] <=  8'h6b;        memory[48710] <=  8'h73;        memory[48711] <=  8'h68;        memory[48712] <=  8'h63;        memory[48713] <=  8'h66;        memory[48714] <=  8'h69;        memory[48715] <=  8'h77;        memory[48716] <=  8'h68;        memory[48717] <=  8'h61;        memory[48718] <=  8'h74;        memory[48719] <=  8'h61;        memory[48720] <=  8'h6e;        memory[48721] <=  8'h61;        memory[48722] <=  8'h62;        memory[48723] <=  8'h61;        memory[48724] <=  8'h63;        memory[48725] <=  8'h61;        memory[48726] <=  8'h74;        memory[48727] <=  8'h61;        memory[48728] <=  8'h62;        memory[48729] <=  8'h61;        memory[48730] <=  8'h72;        memory[48731] <=  8'h63;        memory[48732] <=  8'h61;        memory[48733] <=  8'h68;        memory[48734] <=  8'h64;        memory[48735] <=  8'h75;        memory[48736] <=  8'h63;        memory[48737] <=  8'h74;        memory[48738] <=  8'h61;        memory[48739] <=  8'h64;        memory[48740] <=  8'h61;        memory[48741] <=  8'h61;        memory[48742] <=  8'h63;        memory[48743] <=  8'h61;        memory[48744] <=  8'h72;        memory[48745] <=  8'h62;        memory[48746] <=  8'h61;        memory[48747] <=  8'h72;        memory[48748] <=  8'h74;        memory[48749] <=  8'h78;        memory[48750] <=  8'h61;        memory[48751] <=  8'h74;        memory[48752] <=  8'h6b;        memory[48753] <=  8'h73;        memory[48754] <=  8'h68;        memory[48755] <=  8'h63;        memory[48756] <=  8'h66;        memory[48757] <=  8'h69;        memory[48758] <=  8'h77;        memory[48759] <=  8'h68;        memory[48760] <=  8'h61;        memory[48761] <=  8'h74;        memory[48762] <=  8'h61;        memory[48763] <=  8'h6e;        memory[48764] <=  8'h61;        memory[48765] <=  8'h62;        memory[48766] <=  8'h61;        memory[48767] <=  8'h63;        memory[48768] <=  8'h61;        memory[48769] <=  8'h74;        memory[48770] <=  8'h61;        memory[48771] <=  8'h62;        memory[48772] <=  8'h61;        memory[48773] <=  8'h72;        memory[48774] <=  8'h63;        memory[48775] <=  8'h61;        memory[48776] <=  8'h68;        memory[48777] <=  8'h64;        memory[48778] <=  8'h75;        memory[48779] <=  8'h63;        memory[48780] <=  8'h74;        memory[48781] <=  8'h61;        memory[48782] <=  8'h64;        memory[48783] <=  8'h61;        memory[48784] <=  8'h61;        memory[48785] <=  8'h63;        memory[48786] <=  8'h61;        memory[48787] <=  8'h72;        memory[48788] <=  8'h62;        memory[48789] <=  8'h61;        memory[48790] <=  8'h72;        memory[48791] <=  8'h74;        memory[48792] <=  8'h78;        memory[48793] <=  8'h61;        memory[48794] <=  8'h74;        memory[48795] <=  8'h6b;        memory[48796] <=  8'h73;        memory[48797] <=  8'h68;        memory[48798] <=  8'h63;        memory[48799] <=  8'h66;        memory[48800] <=  8'h69;        memory[48801] <=  8'h77;        memory[48802] <=  8'h68;        memory[48803] <=  8'h61;        memory[48804] <=  8'h74;        memory[48805] <=  8'h61;        memory[48806] <=  8'h6e;        memory[48807] <=  8'h61;        memory[48808] <=  8'h62;        memory[48809] <=  8'h61;        memory[48810] <=  8'h63;        memory[48811] <=  8'h61;        memory[48812] <=  8'h74;        memory[48813] <=  8'h61;        memory[48814] <=  8'h62;        memory[48815] <=  8'h61;        memory[48816] <=  8'h72;        memory[48817] <=  8'h63;        memory[48818] <=  8'h61;        memory[48819] <=  8'h68;        memory[48820] <=  8'h64;        memory[48821] <=  8'h75;        memory[48822] <=  8'h63;        memory[48823] <=  8'h74;        memory[48824] <=  8'h61;        memory[48825] <=  8'h64;        memory[48826] <=  8'h61;        memory[48827] <=  8'h61;        memory[48828] <=  8'h63;        memory[48829] <=  8'h61;        memory[48830] <=  8'h72;        memory[48831] <=  8'h62;        memory[48832] <=  8'h61;        memory[48833] <=  8'h72;        memory[48834] <=  8'h74;        memory[48835] <=  8'h78;        memory[48836] <=  8'h61;        memory[48837] <=  8'h74;        memory[48838] <=  8'h6b;        memory[48839] <=  8'h73;        memory[48840] <=  8'h68;        memory[48841] <=  8'h63;        memory[48842] <=  8'h66;        memory[48843] <=  8'h69;        memory[48844] <=  8'h77;        memory[48845] <=  8'h68;        memory[48846] <=  8'h61;        memory[48847] <=  8'h74;        memory[48848] <=  8'h61;        memory[48849] <=  8'h6e;        memory[48850] <=  8'h61;        memory[48851] <=  8'h62;        memory[48852] <=  8'h61;        memory[48853] <=  8'h63;        memory[48854] <=  8'h61;        memory[48855] <=  8'h74;        memory[48856] <=  8'h61;        memory[48857] <=  8'h62;        memory[48858] <=  8'h61;        memory[48859] <=  8'h72;        memory[48860] <=  8'h63;        memory[48861] <=  8'h61;        memory[48862] <=  8'h68;        memory[48863] <=  8'h64;        memory[48864] <=  8'h75;        memory[48865] <=  8'h63;        memory[48866] <=  8'h74;        memory[48867] <=  8'h61;        memory[48868] <=  8'h64;        memory[48869] <=  8'h61;        memory[48870] <=  8'h61;        memory[48871] <=  8'h63;        memory[48872] <=  8'h61;        memory[48873] <=  8'h72;        memory[48874] <=  8'h62;        memory[48875] <=  8'h61;        memory[48876] <=  8'h72;        memory[48877] <=  8'h74;        memory[48878] <=  8'h78;        memory[48879] <=  8'h61;        memory[48880] <=  8'h74;        memory[48881] <=  8'h6b;        memory[48882] <=  8'h73;        memory[48883] <=  8'h68;        memory[48884] <=  8'h63;        memory[48885] <=  8'h66;        memory[48886] <=  8'h69;        memory[48887] <=  8'h77;        memory[48888] <=  8'h68;        memory[48889] <=  8'h61;        memory[48890] <=  8'h74;        memory[48891] <=  8'h61;        memory[48892] <=  8'h6e;        memory[48893] <=  8'h61;        memory[48894] <=  8'h62;        memory[48895] <=  8'h61;        memory[48896] <=  8'h63;        memory[48897] <=  8'h61;        memory[48898] <=  8'h74;        memory[48899] <=  8'h61;        memory[48900] <=  8'h62;        memory[48901] <=  8'h61;        memory[48902] <=  8'h72;        memory[48903] <=  8'h63;        memory[48904] <=  8'h61;        memory[48905] <=  8'h68;        memory[48906] <=  8'h64;        memory[48907] <=  8'h75;        memory[48908] <=  8'h63;        memory[48909] <=  8'h74;        memory[48910] <=  8'h61;        memory[48911] <=  8'h64;        memory[48912] <=  8'h61;        memory[48913] <=  8'h61;        memory[48914] <=  8'h63;        memory[48915] <=  8'h61;        memory[48916] <=  8'h72;        memory[48917] <=  8'h62;        memory[48918] <=  8'h61;        memory[48919] <=  8'h72;        memory[48920] <=  8'h74;        memory[48921] <=  8'h74;        memory[48922] <=  8'h62;        memory[48923] <=  8'h61;        memory[48924] <=  8'h72;        memory[48925] <=  8'h74;        memory[48926] <=  8'h78;        memory[48927] <=  8'h61;        memory[48928] <=  8'h74;        memory[48929] <=  8'h6b;        memory[48930] <=  8'h73;        memory[48931] <=  8'h68;        memory[48932] <=  8'h63;        memory[48933] <=  8'h66;        memory[48934] <=  8'h69;        memory[48935] <=  8'h77;        memory[48936] <=  8'h68;        memory[48937] <=  8'h61;        memory[48938] <=  8'h74;        memory[48939] <=  8'h61;        memory[48940] <=  8'h6e;        memory[48941] <=  8'h61;        memory[48942] <=  8'h62;        memory[48943] <=  8'h61;        memory[48944] <=  8'h63;        memory[48945] <=  8'h61;        memory[48946] <=  8'h74;        memory[48947] <=  8'h61;        memory[48948] <=  8'h62;        memory[48949] <=  8'h61;        memory[48950] <=  8'h72;        memory[48951] <=  8'h63;        memory[48952] <=  8'h61;        memory[48953] <=  8'h68;        memory[48954] <=  8'h64;        memory[48955] <=  8'h75;        memory[48956] <=  8'h63;        memory[48957] <=  8'h74;        memory[48958] <=  8'h61;        memory[48959] <=  8'h64;        memory[48960] <=  8'h61;        memory[48961] <=  8'h61;        memory[48962] <=  8'h63;        memory[48963] <=  8'h61;        memory[48964] <=  8'h72;        memory[48965] <=  8'h63;        memory[48966] <=  8'h74;        memory[48967] <=  8'h72;        memory[48968] <=  8'h63;        memory[48969] <=  8'h61;        memory[48970] <=  8'h74;        memory[48971] <=  8'h72;        memory[48972] <=  8'h63;        memory[48973] <=  8'h61;        memory[48974] <=  8'h74;        memory[48975] <=  8'h63;        memory[48976] <=  8'h62;        memory[48977] <=  8'h61;        memory[48978] <=  8'h74;        memory[48979] <=  8'h62;        memory[48980] <=  8'h72;        memory[48981] <=  8'h63;        memory[48982] <=  8'h61;        memory[48983] <=  8'h72;        memory[48984] <=  8'h62;        memory[48985] <=  8'h78;        memory[48986] <=  8'h74;        memory[48987] <=  8'h61;        memory[48988] <=  8'h72;        memory[48989] <=  8'h64;        memory[48990] <=  8'h66;        memory[48991] <=  8'h73;        memory[48992] <=  8'h67;        memory[48993] <=  8'h76;        memory[48994] <=  8'h68;        memory[48995] <=  8'h62;        memory[48996] <=  8'h6b;        memory[48997] <=  8'h6a;        memory[48998] <=  8'h6e;        memory[48999] <=  8'h6d;        memory[49000] <=  8'h62;        memory[49001] <=  8'h76;        memory[49002] <=  8'h78;        memory[49003] <=  8'h63;        memory[49004] <=  8'h73;        memory[49005] <=  8'h66;        memory[49006] <=  8'h72;        memory[49007] <=  8'h74;        memory[49008] <=  8'h79;        memory[49009] <=  8'h75;        memory[49010] <=  8'h6a;        memory[49011] <=  8'h6e;        memory[49012] <=  8'h62;        memory[49013] <=  8'h76;        memory[49014] <=  8'h63;        memory[49015] <=  8'h64;        memory[49016] <=  8'h74;        memory[49017] <=  8'h79;        memory[49018] <=  8'h75;        memory[49019] <=  8'h69;        memory[49020] <=  8'h6b;        memory[49021] <=  8'h6d;        memory[49022] <=  8'h6e;        memory[49023] <=  8'h62;        memory[49024] <=  8'h76;        memory[49025] <=  8'h63;        memory[49026] <=  8'h78;        memory[49027] <=  8'h73;        memory[49028] <=  8'h64;        memory[49029] <=  8'h72;        memory[49030] <=  8'h74;        memory[49031] <=  8'h79;        memory[49032] <=  8'h75;        memory[49033] <=  8'h69;        memory[49034] <=  8'h6b;        memory[49035] <=  8'h6d;        memory[49036] <=  8'h6e;        memory[49037] <=  8'h62;        memory[49038] <=  8'h76;        memory[49039] <=  8'h63;        memory[49040] <=  8'h73;        memory[49041] <=  8'h77;        memory[49042] <=  8'h33;        memory[49043] <=  8'h34;        memory[49044] <=  8'h35;        memory[49045] <=  8'h36;        memory[49046] <=  8'h37;        memory[49047] <=  8'h38;        memory[49048] <=  8'h69;        memory[49049] <=  8'h6b;        memory[49050] <=  8'h6d;        memory[49051] <=  8'h6e;        memory[49052] <=  8'h62;        memory[49053] <=  8'h76;        memory[49054] <=  8'h63;        memory[49055] <=  8'h64;        memory[49056] <=  8'h65;        memory[49057] <=  8'h72;        memory[49058] <=  8'h36;        memory[49059] <=  8'h37;        memory[49060] <=  8'h38;        memory[49061] <=  8'h69;        memory[49062] <=  8'h6f;        memory[49063] <=  8'h6b;        memory[49064] <=  8'h6a;        memory[49065] <=  8'h6e;        memory[49066] <=  8'h62;        memory[49067] <=  8'h76;        memory[49068] <=  8'h63;        memory[49069] <=  8'h64;        memory[49070] <=  8'h72;        memory[49071] <=  8'h74;        memory[49072] <=  8'h79;        memory[49073] <=  8'h75;        memory[49074] <=  8'h73;        memory[49075] <=  8'h6a;        memory[49076] <=  8'h63;        memory[49077] <=  8'h6e;        memory[49078] <=  8'h62;        memory[49079] <=  8'h64;        memory[49080] <=  8'h66;        memory[49081] <=  8'h73;        memory[49082] <=  8'h74;        memory[49083] <=  8'h79;        memory[49084] <=  8'h75;        memory[49085] <=  8'h61;        memory[49086] <=  8'h69;        memory[49087] <=  8'h6b;        memory[49088] <=  8'h78;        memory[49089] <=  8'h6d;        memory[49090] <=  8'h6e;        memory[49091] <=  8'h73;        memory[49092] <=  8'h6a;        memory[49093] <=  8'h6f;        memory[49094] <=  8'h64;        memory[49095] <=  8'h6c;        memory[49096] <=  8'h63;        memory[49097] <=  8'h78;        memory[49098] <=  8'h2c;        memory[49099] <=  8'h6d;        memory[49100] <=  8'h73;        memory[49101] <=  8'h6b;        memory[49102] <=  8'h64;        memory[49103] <=  8'h6c;        memory[49104] <=  8'h70;        memory[49105] <=  8'h5b;        memory[49106] <=  8'h3b;        memory[49107] <=  8'h73;        memory[49108] <=  8'h6c;        memory[49109] <=  8'h64;        memory[49110] <=  8'h70;        memory[49111] <=  8'h76;        memory[49112] <=  8'h63;        memory[49113] <=  8'h5b;        memory[49114] <=  8'h78;        memory[49115] <=  8'h76;        memory[49116] <=  8'h63;        memory[49117] <=  8'h5b;        memory[49118] <=  8'h78;        memory[49119] <=  8'h70;        memory[49120] <=  8'h6f;        memory[49121] <=  8'h20;        memory[49122] <=  8'h62;        memory[49123] <=  8'h61;        memory[49124] <=  8'h72;        memory[49125] <=  8'h74;        memory[49126] <=  8'h74;        memory[49127] <=  8'h62;        memory[49128] <=  8'h61;        memory[49129] <=  8'h72;        memory[49130] <=  8'h74;        memory[49131] <=  8'h78;        memory[49132] <=  8'h61;        memory[49133] <=  8'h74;        memory[49134] <=  8'h6b;        memory[49135] <=  8'h73;        memory[49136] <=  8'h68;        memory[49137] <=  8'h63;        memory[49138] <=  8'h66;        memory[49139] <=  8'h69;        memory[49140] <=  8'h77;        memory[49141] <=  8'h68;        memory[49142] <=  8'h61;        memory[49143] <=  8'h69;        memory[49144] <=  8'h6a;        memory[49145] <=  8'h78;        memory[49146] <=  8'h5d;        memory[49147] <=  8'h65;        memory[49148] <=  8'h6b;        memory[49149] <=  8'h6f;        memory[49150] <=  8'h39;        memory[49151] <=  8'h64;        memory[49152] <=  8'h75;        memory[49153] <=  8'h38;        memory[49154] <=  8'h79;        memory[49155] <=  8'h20;        memory[49156] <=  8'h37;        memory[49157] <=  8'h63;        memory[49158] <=  8'h67;        memory[49159] <=  8'h78;        memory[49160] <=  8'h63;        memory[49161] <=  8'h75;        memory[49162] <=  8'h68;        memory[49163] <=  8'h69;        memory[49164] <=  8'h6a;        memory[49165] <=  8'h77;        memory[49166] <=  8'h69;        memory[49167] <=  8'h64;        memory[49168] <=  8'h66;        memory[49169] <=  8'h68;        memory[49170] <=  8'h75;        memory[49171] <=  8'h76;        memory[49172] <=  8'h64;        memory[49173] <=  8'h62;        memory[49174] <=  8'h66;        memory[49175] <=  8'h6a;        memory[49176] <=  8'h6e;        memory[49177] <=  8'h6b;        memory[49178] <=  8'h6a;        memory[49179] <=  8'h65;        memory[49180] <=  8'h38;        memory[49181] <=  8'h66;        memory[49182] <=  8'h37;        memory[49183] <=  8'h67;        memory[49184] <=  8'h79;        memory[49185] <=  8'h76;        memory[49186] <=  8'h63;        memory[49187] <=  8'h68;        memory[49188] <=  8'h69;        memory[49189] <=  8'h6a;        memory[49190] <=  8'h33;        memory[49191] <=  8'h65;        memory[49192] <=  8'h67;        memory[49193] <=  8'h79;        memory[49194] <=  8'h72;        memory[49195] <=  8'h64;        memory[49196] <=  8'h62;        memory[49197] <=  8'h6e;        memory[49198] <=  8'h63;        memory[49199] <=  8'h7a;        memory[49200] <=  8'h6a;        memory[49201] <=  8'h6f;        memory[49202] <=  8'h66;        memory[49203] <=  8'h78;        memory[49204] <=  8'h6a;        memory[49205] <=  8'h69;        memory[49206] <=  8'h63;        memory[49207] <=  8'h68;        memory[49208] <=  8'h62;        memory[49209] <=  8'h6e;        memory[49210] <=  8'h6d;        memory[49211] <=  8'h63;        memory[49212] <=  8'h73;        memory[49213] <=  8'h6c;        memory[49214] <=  8'h6b;        memory[49215] <=  8'h6a;        memory[49216] <=  8'h69;        memory[49217] <=  8'h68;        memory[49218] <=  8'h76;        memory[49219] <=  8'h75;        memory[49220] <=  8'h69;        memory[49221] <=  8'h64;        memory[49222] <=  8'h68;        memory[49223] <=  8'h75;        memory[49224] <=  8'h67;        memory[49225] <=  8'h79;        memory[49226] <=  8'h62;        memory[49227] <=  8'h68;        memory[49228] <=  8'h65;        memory[49229] <=  8'h6a;        memory[49230] <=  8'h72;        memory[49231] <=  8'h6b;        memory[49232] <=  8'h6a;        memory[49233] <=  8'h6f;        memory[49234] <=  8'h64;        memory[49235] <=  8'h67;        memory[49236] <=  8'h69;        memory[49237] <=  8'h75;        memory[49238] <=  8'h69;        memory[49239] <=  8'h67;        memory[49240] <=  8'h76;        memory[49241] <=  8'h79;        memory[49242] <=  8'h75;        memory[49243] <=  8'h67;        memory[49244] <=  8'h78;        memory[49245] <=  8'h68;        memory[49246] <=  8'h63;        memory[49247] <=  8'h20;        memory[49248] <=  8'h20;        memory[49249] <=  8'h20;        memory[49250] <=  8'h78;        memory[49251] <=  8'h76;        memory[49252] <=  8'h20;        memory[49253] <=  8'h63;        memory[49254] <=  8'h78;        memory[49255] <=  8'h67;        memory[49256] <=  8'h79;        memory[49257] <=  8'h63;        memory[49258] <=  8'h75;        memory[49259] <=  8'h68;        memory[49260] <=  8'h6a;        memory[49261] <=  8'h6b;        memory[49262] <=  8'h61;        memory[49263] <=  8'h6c;        memory[49264] <=  8'h78;        memory[49265] <=  8'h76;        memory[49266] <=  8'h70;        memory[49267] <=  8'h6f;        memory[49268] <=  8'h69;        memory[49269] <=  8'h6a;        memory[49270] <=  8'h69;        memory[49271] <=  8'h68;        memory[49272] <=  8'h6a;        memory[49273] <=  8'h62;        memory[49274] <=  8'h77;        memory[49275] <=  8'h65;        memory[49276] <=  8'h6e;        memory[49277] <=  8'h61;        memory[49278] <=  8'h66;        memory[49279] <=  8'h6d;        memory[49280] <=  8'h64;        memory[49281] <=  8'h6b;        memory[49282] <=  8'h6d;        memory[49283] <=  8'h76;        memory[49284] <=  8'h6c;        memory[49285] <=  8'h63;        memory[49286] <=  8'h6f;        memory[49287] <=  8'h64;        memory[49288] <=  8'h69;        memory[49289] <=  8'h75;        memory[49290] <=  8'h68;        memory[49291] <=  8'h73;        memory[49292] <=  8'h66;        memory[49293] <=  8'h65;        memory[49294] <=  8'h62;        memory[49295] <=  8'h6e;        memory[49296] <=  8'h64;        memory[49297] <=  8'h73;        memory[49298] <=  8'h63;        memory[49299] <=  8'h6b;        memory[49300] <=  8'h20;        memory[49301] <=  8'h78;        memory[49302] <=  8'h6a;        memory[49303] <=  8'h78;        memory[49304] <=  8'h63;        memory[49305] <=  8'h73;        memory[49306] <=  8'h64;        memory[49307] <=  8'h66;        memory[49308] <=  8'h6b;        memory[49309] <=  8'h64;        memory[49310] <=  8'h6e;        memory[49311] <=  8'h6d;        memory[49312] <=  8'h64;        memory[49313] <=  8'h73;        memory[49314] <=  8'h63;        memory[49315] <=  8'h6b;        memory[49316] <=  8'h78;        memory[49317] <=  8'h6c;        memory[49318] <=  8'h6f;        memory[49319] <=  8'h66;        memory[49320] <=  8'h6a;        memory[49321] <=  8'h69;        memory[49322] <=  8'h61;        memory[49323] <=  8'h62;        memory[49324] <=  8'h6e;        memory[49325] <=  8'h20;        memory[49326] <=  8'h78;        memory[49327] <=  8'h6b;        memory[49328] <=  8'h6d;        memory[49329] <=  8'h20;        memory[49330] <=  8'h6f;        memory[49331] <=  8'h63;        memory[49332] <=  8'h76;        memory[49333] <=  8'h73;        memory[49334] <=  8'h64;        memory[49335] <=  8'h69;        memory[49336] <=  8'h66;        memory[49337] <=  8'h68;        memory[49338] <=  8'h65;        memory[49339] <=  8'h71;        memory[49340] <=  8'h6a;        memory[49341] <=  8'h77;        memory[49342] <=  8'h62;        memory[49343] <=  8'h65;        memory[49344] <=  8'h6e;        memory[49345] <=  8'h20;        memory[49346] <=  8'h6d;        memory[49347] <=  8'h64;        memory[49348] <=  8'h73;        memory[49349] <=  8'h6c;        memory[49350] <=  8'h76;        memory[49351] <=  8'h6b;        memory[49352] <=  8'h63;        memory[49353] <=  8'h78;        memory[49354] <=  8'h20;        memory[49355] <=  8'h6f;        memory[49356] <=  8'h78;        memory[49357] <=  8'h69;        memory[49358] <=  8'h63;        memory[49359] <=  8'h6a;        memory[49360] <=  8'h76;        memory[49361] <=  8'h64;        memory[49362] <=  8'h66;        memory[49363] <=  8'h65;        memory[49364] <=  8'h71;        memory[49365] <=  8'h6e;        memory[49366] <=  8'h20;        memory[49367] <=  8'h64;        memory[49368] <=  8'h6d;        memory[49369] <=  8'h73;        memory[49370] <=  8'h6c;        memory[49371] <=  8'h63;        memory[49372] <=  8'h78;        memory[49373] <=  8'h6b;        memory[49374] <=  8'h20;        memory[49375] <=  8'h6f;        memory[49376] <=  8'h78;        memory[49377] <=  8'h63;        memory[49378] <=  8'h76;        memory[49379] <=  8'h6a;        memory[49380] <=  8'h64;        memory[49381] <=  8'h62;        memory[49382] <=  8'h71;        memory[49383] <=  8'h77;        memory[49384] <=  8'h65;        memory[49385] <=  8'h6e;        memory[49386] <=  8'h6d;        memory[49387] <=  8'h64;        memory[49388] <=  8'h6c;        memory[49389] <=  8'h73;        memory[49390] <=  8'h2c;        memory[49391] <=  8'h76;        memory[49392] <=  8'h63;        memory[49393] <=  8'h78;        memory[49394] <=  8'h20;        memory[49395] <=  8'h63;        memory[49396] <=  8'h6f;        memory[49397] <=  8'h69;        memory[49398] <=  8'h76;        memory[49399] <=  8'h68;        memory[49400] <=  8'h73;        memory[49401] <=  8'h64;        memory[49402] <=  8'h62;        memory[49403] <=  8'h71;        memory[49404] <=  8'h77;        memory[49405] <=  8'h65;        memory[49406] <=  8'h6e;        memory[49407] <=  8'h64;        memory[49408] <=  8'h6b;        memory[49409] <=  8'h73;        memory[49410] <=  8'h76;        memory[49411] <=  8'h6f;        memory[49412] <=  8'h63;        memory[49413] <=  8'h20;        memory[49414] <=  8'h76;        memory[49415] <=  8'h69;        memory[49416] <=  8'h75;        memory[49417] <=  8'h69;        memory[49418] <=  8'h68;        memory[49419] <=  8'h63;        memory[49420] <=  8'h78;        memory[49421] <=  8'h69;        memory[49422] <=  8'h6f;        memory[49423] <=  8'h76;        memory[49424] <=  8'h73;        memory[49425] <=  8'h64;        memory[49426] <=  8'h61;        memory[49427] <=  8'h64;        memory[49428] <=  8'h6e;        memory[49429] <=  8'h77;        memory[49430] <=  8'h71;        memory[49431] <=  8'h6b;        memory[49432] <=  8'h6c;        memory[49433] <=  8'h73;        memory[49434] <=  8'h76;        memory[49435] <=  8'h6e;        memory[49436] <=  8'h62;        memory[49437] <=  8'h20;        memory[49438] <=  8'h64;        memory[49439] <=  8'h66;        memory[49440] <=  8'h6a;        memory[49441] <=  8'h6b;        memory[49442] <=  8'h71;        memory[49443] <=  8'h64;        memory[49444] <=  8'h77;        memory[49445] <=  8'h65;        memory[49446] <=  8'h6e;        memory[49447] <=  8'h62;        memory[49448] <=  8'h20;        memory[49449] <=  8'h64;        memory[49450] <=  8'h73;        memory[49451] <=  8'h76;        memory[49452] <=  8'h68;        memory[49453] <=  8'h64;        memory[49454] <=  8'h61;        memory[49455] <=  8'h71;        memory[49456] <=  8'h77;        memory[49457] <=  8'h6a;        memory[49458] <=  8'h65;        memory[49459] <=  8'h6e;        memory[49460] <=  8'h64;        memory[49461] <=  8'h20;        memory[49462] <=  8'h61;        memory[49463] <=  8'h63;        memory[49464] <=  8'h62;        memory[49465] <=  8'h68;        memory[49466] <=  8'h64;        memory[49467] <=  8'h61;        memory[49468] <=  8'h77;        memory[49469] <=  8'h71;        memory[49470] <=  8'h6e;        memory[49471] <=  8'h20;        memory[49472] <=  8'h62;        memory[49473] <=  8'h73;        memory[49474] <=  8'h76;        memory[49475] <=  8'h61;        memory[49476] <=  8'h67;        memory[49477] <=  8'h76;        memory[49478] <=  8'h68;        memory[49479] <=  8'h67;        memory[49480] <=  8'h61;        memory[49481] <=  8'h73;        memory[49482] <=  8'h6a;        memory[49483] <=  8'h6b;        memory[49484] <=  8'h63;        memory[49485] <=  8'h78;        memory[49486] <=  8'h76;        memory[49487] <=  8'h6e;        memory[49488] <=  8'h73;        memory[49489] <=  8'h64;        memory[49490] <=  8'h20;        memory[49491] <=  8'h66;        memory[49492] <=  8'h62;        memory[49493] <=  8'h64;        memory[49494] <=  8'h61;        memory[49495] <=  8'h73;        memory[49496] <=  8'h76;        memory[49497] <=  8'h67;        memory[49498] <=  8'h63;        memory[49499] <=  8'h79;        memory[49500] <=  8'h7a;        memory[49501] <=  8'h78;        memory[49502] <=  8'h79;        memory[49503] <=  8'h75;        memory[49504] <=  8'h20;        memory[49505] <=  8'h69;        memory[49506] <=  8'h6a;        memory[49507] <=  8'h64;        memory[49508] <=  8'h66;        memory[49509] <=  8'h6b;        memory[49510] <=  8'h61;        memory[49511] <=  8'h64;        memory[49512] <=  8'h63;        memory[49513] <=  8'h78;        memory[49514] <=  8'h68;        memory[49515] <=  8'h20;        memory[49516] <=  8'h67;        memory[49517] <=  8'h61;        memory[49518] <=  8'h68;        memory[49519] <=  8'h75;        memory[49520] <=  8'h64;        memory[49521] <=  8'h73;        memory[49522] <=  8'h69;        memory[49523] <=  8'h6a;        memory[49524] <=  8'h61;        memory[49525] <=  8'h6b;        memory[49526] <=  8'h63;        memory[49527] <=  8'h62;        memory[49528] <=  8'h61;        memory[49529] <=  8'h72;        memory[49530] <=  8'h73;        memory[49531] <=  8'h68;        memory[49532] <=  8'h64;        memory[49533] <=  8'h66;        memory[49534] <=  8'h67;        memory[49535] <=  8'h73;        memory[49536] <=  8'h68;        memory[49537] <=  8'h64;        memory[49538] <=  8'h66;        memory[49539] <=  8'h68;        memory[49540] <=  8'h64;        memory[49541] <=  8'h6a;        memory[49542] <=  8'h68;        memory[49543] <=  8'h62;        memory[49544] <=  8'h67;        memory[49545] <=  8'h63;        memory[49546] <=  8'h61;        memory[49547] <=  8'h66;        memory[49548] <=  8'h73;        memory[49549] <=  8'h79;        memory[49550] <=  8'h67;        memory[49551] <=  8'h6b;        memory[49552] <=  8'h75;        memory[49553] <=  8'h64;        memory[49554] <=  8'h68;        memory[49555] <=  8'h62;        memory[49556] <=  8'h77;        memory[49557] <=  8'h76;        memory[49558] <=  8'h67;        memory[49559] <=  8'h61;        memory[49560] <=  8'h66;        memory[49561] <=  8'h64;        memory[49562] <=  8'h74;        memory[49563] <=  8'h75;        memory[49564] <=  8'h66;        memory[49565] <=  8'h79;        memory[49566] <=  8'h67;        memory[49567] <=  8'h69;        memory[49568] <=  8'h75;        memory[49569] <=  8'h68;        memory[49570] <=  8'h6c;        memory[49571] <=  8'h6a;        memory[49572] <=  8'h62;        memory[49573] <=  8'h6b;        memory[49574] <=  8'h68;        memory[49575] <=  8'h76;        memory[49576] <=  8'h67;        memory[49577] <=  8'h63;        memory[49578] <=  8'h66;        memory[49579] <=  8'h78;        memory[49580] <=  8'h64;        memory[49581] <=  8'h74;        memory[49582] <=  8'h75;        memory[49583] <=  8'h79;        memory[49584] <=  8'h69;        memory[49585] <=  8'h75;        memory[49586] <=  8'h68;        memory[49587] <=  8'h6c;        memory[49588] <=  8'h6a;        memory[49589] <=  8'h6b;        memory[49590] <=  8'h67;        memory[49591] <=  8'h6a;        memory[49592] <=  8'h63;        memory[49593] <=  8'h66;        memory[49594] <=  8'h68;        memory[49595] <=  8'h64;        memory[49596] <=  8'h67;        memory[49597] <=  8'h72;        memory[49598] <=  8'h79;        memory[49599] <=  8'h74;        memory[49600] <=  8'h66;        memory[49601] <=  8'h75;        memory[49602] <=  8'h79;        memory[49603] <=  8'h69;        memory[49604] <=  8'h68;        memory[49605] <=  8'h6c;        memory[49606] <=  8'h62;        memory[49607] <=  8'h6d;        memory[49608] <=  8'h76;        memory[49609] <=  8'h6e;        memory[49610] <=  8'h63;        memory[49611] <=  8'h66;        memory[49612] <=  8'h68;        memory[49613] <=  8'h64;        memory[49614] <=  8'h74;        memory[49615] <=  8'h75;        memory[49616] <=  8'h67;        memory[49617] <=  8'h79;        memory[49618] <=  8'h69;        memory[49619] <=  8'h68;        memory[49620] <=  8'h75;        memory[49621] <=  8'h6a;        memory[49622] <=  8'h6c;        memory[49623] <=  8'h62;        memory[49624] <=  8'h6d;        memory[49625] <=  8'h76;        memory[49626] <=  8'h6e;        memory[49627] <=  8'h63;        memory[49628] <=  8'h66;        memory[49629] <=  8'h68;        memory[49630] <=  8'h67;        memory[49631] <=  8'h79;        memory[49632] <=  8'h68;        memory[49633] <=  8'h75;        memory[49634] <=  8'h6a;        memory[49635] <=  8'h6e;        memory[49636] <=  8'h2c;        memory[49637] <=  8'h62;        memory[49638] <=  8'h6e;        memory[49639] <=  8'h6d;        memory[49640] <=  8'h76;        memory[49641] <=  8'h6e;        memory[49642] <=  8'h63;        memory[49643] <=  8'h66;        memory[49644] <=  8'h68;        memory[49645] <=  8'h74;        memory[49646] <=  8'h79;        memory[49647] <=  8'h69;        memory[49648] <=  8'h75;        memory[49649] <=  8'h6c;        memory[49650] <=  8'h6a;        memory[49651] <=  8'h62;        memory[49652] <=  8'h6d;        memory[49653] <=  8'h76;        memory[49654] <=  8'h6e;        memory[49655] <=  8'h63;        memory[49656] <=  8'h66;        memory[49657] <=  8'h74;        memory[49658] <=  8'h75;        memory[49659] <=  8'h79;        memory[49660] <=  8'h69;        memory[49661] <=  8'h68;        memory[49662] <=  8'h6b;        memory[49663] <=  8'h62;        memory[49664] <=  8'h76;        memory[49665] <=  8'h63;        memory[49666] <=  8'h66;        memory[49667] <=  8'h67;        memory[49668] <=  8'h74;        memory[49669] <=  8'h75;        memory[49670] <=  8'h79;        memory[49671] <=  8'h69;        memory[49672] <=  8'h75;        memory[49673] <=  8'h68;        memory[49674] <=  8'h6a;        memory[49675] <=  8'h6b;        memory[49676] <=  8'h62;        memory[49677] <=  8'h76;        memory[49678] <=  8'h63;        memory[49679] <=  8'h66;        memory[49680] <=  8'h74;        memory[49681] <=  8'h75;        memory[49682] <=  8'h79;        memory[49683] <=  8'h69;        memory[49684] <=  8'h75;        memory[49685] <=  8'h6a;        memory[49686] <=  8'h6b;        memory[49687] <=  8'h6e;        memory[49688] <=  8'h62;        memory[49689] <=  8'h76;        memory[49690] <=  8'h67;        memory[49691] <=  8'h66;        memory[49692] <=  8'h74;        memory[49693] <=  8'h79;        memory[49694] <=  8'h75;        memory[49695] <=  8'h75;        memory[49696] <=  8'h69;        memory[49697] <=  8'h6a;        memory[49698] <=  8'h6b;        memory[49699] <=  8'h68;        memory[49700] <=  8'h62;        memory[49701] <=  8'h6a;        memory[49702] <=  8'h67;        memory[49703] <=  8'h68;        memory[49704] <=  8'h66;        memory[49705] <=  8'h79;        memory[49706] <=  8'h74;        memory[49707] <=  8'h79;        memory[49708] <=  8'h69;        memory[49709] <=  8'h75;        memory[49710] <=  8'h64;        memory[49711] <=  8'h6a;        memory[49712] <=  8'h6b;        memory[49713] <=  8'h68;        memory[49714] <=  8'h63;        memory[49715] <=  8'h7a;        memory[49716] <=  8'h67;        memory[49717] <=  8'h68;        memory[49718] <=  8'h74;        memory[49719] <=  8'h75;        memory[49720] <=  8'h79;        memory[49721] <=  8'h69;        memory[49722] <=  8'h61;        memory[49723] <=  8'h73;        memory[49724] <=  8'h75;        memory[49725] <=  8'h6a;        memory[49726] <=  8'h6b;        memory[49727] <=  8'h62;        memory[49728] <=  8'h6e;        memory[49729] <=  8'h61;        memory[49730] <=  8'h76;        memory[49731] <=  8'h63;        memory[49732] <=  8'h66;        memory[49733] <=  8'h68;        memory[49734] <=  8'h75;        memory[49735] <=  8'h61;        memory[49736] <=  8'h73;        memory[49737] <=  8'h79;        memory[49738] <=  8'h64;        memory[49739] <=  8'h75;        memory[49740] <=  8'h69;        memory[49741] <=  8'h6a;        memory[49742] <=  8'h61;        memory[49743] <=  8'h6b;        memory[49744] <=  8'h62;        memory[49745] <=  8'h63;        memory[49746] <=  8'h78;        memory[49747] <=  8'h68;        memory[49748] <=  8'h67;        memory[49749] <=  8'h79;        memory[49750] <=  8'h75;        memory[49751] <=  8'h7a;        memory[49752] <=  8'h63;        memory[49753] <=  8'h61;        memory[49754] <=  8'h73;        memory[49755] <=  8'h69;        memory[49756] <=  8'h75;        memory[49757] <=  8'h6f;        memory[49758] <=  8'h69;        memory[49759] <=  8'h6a;        memory[49760] <=  8'h61;        memory[49761] <=  8'h6c;        memory[49762] <=  8'h63;        memory[49763] <=  8'h78;        memory[49764] <=  8'h62;        memory[49765] <=  8'h63;        memory[49766] <=  8'h20;        memory[49767] <=  8'h6e;        memory[49768] <=  8'h76;        memory[49769] <=  8'h63;        memory[49770] <=  8'h61;        memory[49771] <=  8'h64;        memory[49772] <=  8'h73;        memory[49773] <=  8'h67;        memory[49774] <=  8'h79;        memory[49775] <=  8'h68;        memory[49776] <=  8'h75;        memory[49777] <=  8'h61;        memory[49778] <=  8'h6a;        memory[49779] <=  8'h6b;        memory[49780] <=  8'h78;        memory[49781] <=  8'h62;        memory[49782] <=  8'h20;        memory[49783] <=  8'h6e;        memory[49784] <=  8'h76;        memory[49785] <=  8'h63;        memory[49786] <=  8'h61;        memory[49787] <=  8'h73;        memory[49788] <=  8'h67;        memory[49789] <=  8'h68;        memory[49790] <=  8'h75;        memory[49791] <=  8'h6a;        memory[49792] <=  8'h6c;        memory[49793] <=  8'h6b;        memory[49794] <=  8'h63;        memory[49795] <=  8'h78;        memory[49796] <=  8'h20;        memory[49797] <=  8'h6a;        memory[49798] <=  8'h6b;        memory[49799] <=  8'h68;        memory[49800] <=  8'h61;        memory[49801] <=  8'h73;        memory[49802] <=  8'h76;        memory[49803] <=  8'h64;        memory[49804] <=  8'h6e;        memory[49805] <=  8'h20;        memory[49806] <=  8'h62;        memory[49807] <=  8'h6e;        memory[49808] <=  8'h6d;        memory[49809] <=  8'h6b;        memory[49810] <=  8'h77;        memory[49811] <=  8'h64;        memory[49812] <=  8'h6f;        memory[49813] <=  8'h77;        memory[49814] <=  8'h69;        memory[49815] <=  8'h6f;        memory[49816] <=  8'h75;        memory[49817] <=  8'h69;        memory[49818] <=  8'h68;        memory[49819] <=  8'h62;        memory[49820] <=  8'h6e;        memory[49821] <=  8'h6b;        memory[49822] <=  8'h77;        memory[49823] <=  8'h69;        memory[49824] <=  8'h6f;        memory[49825] <=  8'h75;        memory[49826] <=  8'h71;        memory[49827] <=  8'h69;        memory[49828] <=  8'h79;        memory[49829] <=  8'h67;        memory[49830] <=  8'h6a;        memory[49831] <=  8'h64;        memory[49832] <=  8'h61;        memory[49833] <=  8'h76;        memory[49834] <=  8'h62;        memory[49835] <=  8'h6e;        memory[49836] <=  8'h6b;        memory[49837] <=  8'h6f;        memory[49838] <=  8'h70;        memory[49839] <=  8'h64;        memory[49840] <=  8'h76;        memory[49841] <=  8'h69;        memory[49842] <=  8'h6f;        memory[49843] <=  8'h75;        memory[49844] <=  8'h69;        memory[49845] <=  8'h48;        memory[49846] <=  8'h42;        memory[49847] <=  8'h6b;        memory[49848] <=  8'h64;        memory[49849] <=  8'h6e;        memory[49850] <=  8'h6c;        memory[49851] <=  8'h71;        memory[49852] <=  8'h6b;        memory[49853] <=  8'h6d;        memory[49854] <=  8'h6a;        memory[49855] <=  8'h70;        memory[49856] <=  8'h69;        memory[49857] <=  8'h6f;        memory[49858] <=  8'h68;        memory[49859] <=  8'h65;        memory[49860] <=  8'h66;        memory[49861] <=  8'h75;        memory[49862] <=  8'h67;        memory[49863] <=  8'h69;        memory[49864] <=  8'h73;        memory[49865] <=  8'h61;        memory[49866] <=  8'h62;        memory[49867] <=  8'h64;        memory[49868] <=  8'h6b;        memory[49869] <=  8'h6a;        memory[49870] <=  8'h6b;        memory[49871] <=  8'h6c;        memory[49872] <=  8'h6a;        memory[49873] <=  8'h69;        memory[49874] <=  8'h73;        memory[49875] <=  8'h6f;        memory[49876] <=  8'h71;        memory[49877] <=  8'h68;        memory[49878] <=  8'h77;        memory[49879] <=  8'h67;        memory[49880] <=  8'h69;        memory[49881] <=  8'h79;        memory[49882] <=  8'h6a;        memory[49883] <=  8'h64;        memory[49884] <=  8'h76;        memory[49885] <=  8'h62;        memory[49886] <=  8'h6e;        memory[49887] <=  8'h61;        memory[49888] <=  8'h73;        memory[49889] <=  8'h66;        memory[49890] <=  8'h6c;        memory[49891] <=  8'h6b;        memory[49892] <=  8'h64;        memory[49893] <=  8'h6a;        memory[49894] <=  8'h68;        memory[49895] <=  8'h63;        memory[49896] <=  8'h67;        memory[49897] <=  8'h6a;        memory[49898] <=  8'h76;        memory[49899] <=  8'h73;        memory[49900] <=  8'h64;        memory[49901] <=  8'h62;        memory[49902] <=  8'h62;        memory[49903] <=  8'h61;        memory[49904] <=  8'h72;        memory[49905] <=  8'h62;        memory[49906] <=  8'h62;        memory[49907] <=  8'h73;        memory[49908] <=  8'h62;        memory[49909] <=  8'h67;        memory[49910] <=  8'h73;        memory[49911] <=  8'h66;        memory[49912] <=  8'h67;        memory[49913] <=  8'h61;        memory[49914] <=  8'h68;        memory[49915] <=  8'h66;        memory[49916] <=  8'h73;        memory[49917] <=  8'h68;        memory[49918] <=  8'h61;        memory[49919] <=  8'h66;        memory[49920] <=  8'h73;        memory[49921] <=  8'h66;        memory[49922] <=  8'h68;        memory[49923] <=  8'h61;        memory[49924] <=  8'h69;        memory[49925] <=  8'h64;        memory[49926] <=  8'h75;        memory[49927] <=  8'h67;        memory[49928] <=  8'h64;        memory[49929] <=  8'h77;        memory[49930] <=  8'h62;        memory[49931] <=  8'h61;        memory[49932] <=  8'h62;        memory[49933] <=  8'h72;        memory[49934] <=  8'h62;        memory[49935] <=  8'h61;        memory[49936] <=  8'h62;        memory[49937] <=  8'h62;        memory[49938] <=  8'h74;        memory[49939] <=  8'h62;        memory[49940] <=  8'h62;        memory[49941] <=  8'h62;        memory[49942] <=  8'h62;        memory[49943] <=  8'h62;        memory[49944] <=  8'h62;        memory[49945] <=  8'h62;        memory[49946] <=  8'h62;        memory[49947] <=  8'h61;        memory[49948] <=  8'h62;        memory[49949] <=  8'h62;        memory[49950] <=  8'h72;        memory[49951] <=  8'h74;        memory[49952] <=  8'h62;        memory[49953] <=  8'h62;        memory[49954] <=  8'h61;        memory[49955] <=  8'h62;        memory[49956] <=  8'h72;        memory[49957] <=  8'h62;        memory[49958] <=  8'h74;        memory[49959] <=  8'h62;        memory[49960] <=  8'h62;        memory[49961] <=  8'h62;        memory[49962] <=  8'h63;        memory[49963] <=  8'h61;        memory[49964] <=  8'h72;        memory[49965] <=  8'h74;        memory[49966] <=  8'h73;        memory[49967] <=  8'h62;        memory[49968] <=  8'h61;        memory[49969] <=  8'h72;        memory[49970] <=  8'h74;        memory[49971] <=  8'h74;        memory[49972] <=  8'h62;        memory[49973] <=  8'h61;        memory[49974] <=  8'h72;        memory[49975] <=  8'h74;        memory[49976] <=  8'h78;        memory[49977] <=  8'h61;        memory[49978] <=  8'h74;        memory[49979] <=  8'h6b;        memory[49980] <=  8'h73;        memory[49981] <=  8'h68;        memory[49982] <=  8'h63;        memory[49983] <=  8'h66;        memory[49984] <=  8'h69;        memory[49985] <=  8'h77;        memory[49986] <=  8'h68;        memory[49987] <=  8'h61;        memory[49988] <=  8'h74;        memory[49989] <=  8'h61;        memory[49990] <=  8'h6e;        memory[49991] <=  8'h61;        memory[49992] <=  8'h62;        memory[49993] <=  8'h61;        memory[49994] <=  8'h63;        memory[49995] <=  8'h61;        memory[49996] <=  8'h74;        memory[49997] <=  8'h61;        memory[49998] <=  8'h62;        memory[49999] <=  8'h61;        memory[50000] <=  8'h72;        memory[50001] <=  8'h63;        memory[50002] <=  8'h61;        memory[50003] <=  8'h68;        memory[50004] <=  8'h64;        memory[50005] <=  8'h75;        memory[50006] <=  8'h63;        memory[50007] <=  8'h74;        memory[50008] <=  8'h61;        memory[50009] <=  8'h64;        memory[50010] <=  8'h61;        memory[50011] <=  8'h61;        memory[50012] <=  8'h63;        memory[50013] <=  8'h61;        memory[50014] <=  8'h72;        memory[50015] <=  8'h63;        memory[50016] <=  8'h74;        memory[50017] <=  8'h72;        memory[50018] <=  8'h63;        memory[50019] <=  8'h61;        memory[50020] <=  8'h74;        memory[50021] <=  8'h72;        memory[50022] <=  8'h63;        memory[50023] <=  8'h61;        memory[50024] <=  8'h74;        memory[50025] <=  8'h63;        memory[50026] <=  8'h62;        memory[50027] <=  8'h61;        memory[50028] <=  8'h74;        memory[50029] <=  8'h62;        memory[50030] <=  8'h72;        memory[50031] <=  8'h63;        memory[50032] <=  8'h61;        memory[50033] <=  8'h74;        memory[50034] <=  8'h72;        memory[50035] <=  8'h6e;        memory[50036] <=  8'h62;        memory[50037] <=  8'h61;        memory[50038] <=  8'h63;        memory[50039] <=  8'h61;        memory[50040] <=  8'h74;        memory[50041] <=  8'h79;        memory[50042] <=  8'h73;        memory[50043] <=  8'h6e;        memory[50044] <=  8'h63;        memory[50045] <=  8'h74;        memory[50046] <=  8'h61;        memory[50047] <=  8'h6e;        memory[50048] <=  8'h62;        memory[50049] <=  8'h61;        memory[50050] <=  8'h63;        memory[50051] <=  8'h72;        memory[50052] <=  8'h6e;        memory[50053] <=  8'h74;        memory[50054] <=  8'h61;        memory[50055] <=  8'h62;        memory[50056] <=  8'h74;        memory[50057] <=  8'h6e;        memory[50058] <=  8'h61;        memory[50059] <=  8'h72;        memory[50060] <=  8'h62;        memory[50061] <=  8'h78;        memory[50062] <=  8'h74;        memory[50063] <=  8'h61;        memory[50064] <=  8'h72;        memory[50065] <=  8'h62;        memory[50066] <=  8'h61;        memory[50067] <=  8'h72;        memory[50068] <=  8'h74;        memory[50069] <=  8'h74;        memory[50070] <=  8'h62;        memory[50071] <=  8'h61;        memory[50072] <=  8'h72;        memory[50073] <=  8'h74;        memory[50074] <=  8'h78;        memory[50075] <=  8'h61;        memory[50076] <=  8'h74;        memory[50077] <=  8'h6b;        memory[50078] <=  8'h73;        memory[50079] <=  8'h68;        memory[50080] <=  8'h63;        memory[50081] <=  8'h66;        memory[50082] <=  8'h69;        memory[50083] <=  8'h77;        memory[50084] <=  8'h68;        memory[50085] <=  8'h61;        memory[50086] <=  8'h74;        memory[50087] <=  8'h61;        memory[50088] <=  8'h6e;        memory[50089] <=  8'h61;        memory[50090] <=  8'h62;        memory[50091] <=  8'h61;        memory[50092] <=  8'h63;        memory[50093] <=  8'h61;        memory[50094] <=  8'h74;        memory[50095] <=  8'h61;        memory[50096] <=  8'h62;        memory[50097] <=  8'h61;        memory[50098] <=  8'h72;        memory[50099] <=  8'h63;        memory[50100] <=  8'h61;        memory[50101] <=  8'h68;        memory[50102] <=  8'h64;        memory[50103] <=  8'h75;        memory[50104] <=  8'h63;        memory[50105] <=  8'h74;        memory[50106] <=  8'h61;        memory[50107] <=  8'h64;        memory[50108] <=  8'h61;        memory[50109] <=  8'h61;        memory[50110] <=  8'h63;        memory[50111] <=  8'h61;        memory[50112] <=  8'h72;        memory[50113] <=  8'h63;        memory[50114] <=  8'h74;        memory[50115] <=  8'h72;        memory[50116] <=  8'h63;        memory[50117] <=  8'h61;        memory[50118] <=  8'h74;        memory[50119] <=  8'h72;        memory[50120] <=  8'h63;        memory[50121] <=  8'h61;        memory[50122] <=  8'h74;        memory[50123] <=  8'h63;        memory[50124] <=  8'h62;        memory[50125] <=  8'h61;        memory[50126] <=  8'h74;        memory[50127] <=  8'h62;        memory[50128] <=  8'h72;        memory[50129] <=  8'h63;        memory[50130] <=  8'h61;        memory[50131] <=  8'h74;        memory[50132] <=  8'h72;        memory[50133] <=  8'h6e;        memory[50134] <=  8'h62;        memory[50135] <=  8'h61;        memory[50136] <=  8'h63;        memory[50137] <=  8'h61;        memory[50138] <=  8'h74;        memory[50139] <=  8'h79;        memory[50140] <=  8'h73;        memory[50141] <=  8'h6e;        memory[50142] <=  8'h63;        memory[50143] <=  8'h74;        memory[50144] <=  8'h61;        memory[50145] <=  8'h6e;        memory[50146] <=  8'h62;        memory[50147] <=  8'h61;        memory[50148] <=  8'h63;        memory[50149] <=  8'h72;        memory[50150] <=  8'h6e;        memory[50151] <=  8'h74;        memory[50152] <=  8'h61;        memory[50153] <=  8'h62;        memory[50154] <=  8'h74;        memory[50155] <=  8'h6e;        memory[50156] <=  8'h61;        memory[50157] <=  8'h72;        memory[50158] <=  8'h62;        memory[50159] <=  8'h78;        memory[50160] <=  8'h74;        memory[50161] <=  8'h61;        memory[50162] <=  8'h72;        memory[50163] <=  8'h62;        memory[50164] <=  8'h61;        memory[50165] <=  8'h72;        memory[50166] <=  8'h74;        memory[50167] <=  8'h74;        memory[50168] <=  8'h62;        memory[50169] <=  8'h61;        memory[50170] <=  8'h72;        memory[50171] <=  8'h74;        memory[50172] <=  8'h78;        memory[50173] <=  8'h61;        memory[50174] <=  8'h74;        memory[50175] <=  8'h6b;        memory[50176] <=  8'h73;        memory[50177] <=  8'h68;        memory[50178] <=  8'h63;        memory[50179] <=  8'h66;        memory[50180] <=  8'h69;        memory[50181] <=  8'h77;        memory[50182] <=  8'h68;        memory[50183] <=  8'h61;        memory[50184] <=  8'h74;        memory[50185] <=  8'h61;        memory[50186] <=  8'h6e;        memory[50187] <=  8'h61;        memory[50188] <=  8'h62;        memory[50189] <=  8'h61;        memory[50190] <=  8'h63;        memory[50191] <=  8'h61;        memory[50192] <=  8'h74;        memory[50193] <=  8'h61;        memory[50194] <=  8'h62;        memory[50195] <=  8'h61;        memory[50196] <=  8'h72;        memory[50197] <=  8'h63;        memory[50198] <=  8'h61;        memory[50199] <=  8'h68;        memory[50200] <=  8'h64;        memory[50201] <=  8'h75;        memory[50202] <=  8'h63;        memory[50203] <=  8'h74;        memory[50204] <=  8'h61;        memory[50205] <=  8'h64;        memory[50206] <=  8'h61;        memory[50207] <=  8'h61;        memory[50208] <=  8'h63;        memory[50209] <=  8'h61;        memory[50210] <=  8'h72;        memory[50211] <=  8'h63;        memory[50212] <=  8'h74;        memory[50213] <=  8'h72;        memory[50214] <=  8'h63;        memory[50215] <=  8'h61;        memory[50216] <=  8'h74;        memory[50217] <=  8'h72;        memory[50218] <=  8'h63;        memory[50219] <=  8'h61;        memory[50220] <=  8'h74;        memory[50221] <=  8'h63;        memory[50222] <=  8'h62;        memory[50223] <=  8'h61;        memory[50224] <=  8'h74;        memory[50225] <=  8'h62;        memory[50226] <=  8'h72;        memory[50227] <=  8'h63;        memory[50228] <=  8'h61;        memory[50229] <=  8'h74;        memory[50230] <=  8'h72;        memory[50231] <=  8'h6e;        memory[50232] <=  8'h62;        memory[50233] <=  8'h61;        memory[50234] <=  8'h63;        memory[50235] <=  8'h61;        memory[50236] <=  8'h74;        memory[50237] <=  8'h79;        memory[50238] <=  8'h73;        memory[50239] <=  8'h6e;        memory[50240] <=  8'h63;        memory[50241] <=  8'h74;        memory[50242] <=  8'h61;        memory[50243] <=  8'h6e;        memory[50244] <=  8'h62;        memory[50245] <=  8'h61;        memory[50246] <=  8'h63;        memory[50247] <=  8'h72;        memory[50248] <=  8'h6e;        memory[50249] <=  8'h74;        memory[50250] <=  8'h61;        memory[50251] <=  8'h62;        memory[50252] <=  8'h74;        memory[50253] <=  8'h6e;        memory[50254] <=  8'h61;        memory[50255] <=  8'h72;        memory[50256] <=  8'h62;        memory[50257] <=  8'h78;        memory[50258] <=  8'h74;        memory[50259] <=  8'h61;        memory[50260] <=  8'h72;        memory[50261] <=  8'h5d;        memory[50262] <=  8'h5d;        memory[50263] <=  8'h65;        memory[50264] <=  8'h66;        memory[50265] <=  8'h77;        memory[50266] <=  8'h65;        memory[50267] <=  8'h5d;        memory[50268] <=  8'h65;        memory[50269] <=  8'h67;        memory[50270] <=  8'h73;        memory[50271] <=  8'h67;        memory[50272] <=  8'h66;        memory[50273] <=  8'h62;        memory[50274] <=  8'h61;        memory[50275] <=  8'h72;        memory[50276] <=  8'h74;        memory[50277] <=  8'h74;        memory[50278] <=  8'h62;        memory[50279] <=  8'h61;        memory[50280] <=  8'h72;        memory[50281] <=  8'h74;        memory[50282] <=  8'h78;        memory[50283] <=  8'h61;        memory[50284] <=  8'h74;        memory[50285] <=  8'h6b;        memory[50286] <=  8'h73;        memory[50287] <=  8'h68;        memory[50288] <=  8'h63;        memory[50289] <=  8'h66;        memory[50290] <=  8'h69;        memory[50291] <=  8'h77;        memory[50292] <=  8'h68;        memory[50293] <=  8'h61;        memory[50294] <=  8'h74;        memory[50295] <=  8'h61;        memory[50296] <=  8'h6e;        memory[50297] <=  8'h61;        memory[50298] <=  8'h62;        memory[50299] <=  8'h61;        memory[50300] <=  8'h63;        memory[50301] <=  8'h61;        memory[50302] <=  8'h74;        memory[50303] <=  8'h61;        memory[50304] <=  8'h62;        memory[50305] <=  8'h61;        memory[50306] <=  8'h72;        memory[50307] <=  8'h63;        memory[50308] <=  8'h61;        memory[50309] <=  8'h68;        memory[50310] <=  8'h64;        memory[50311] <=  8'h75;        memory[50312] <=  8'h63;        memory[50313] <=  8'h74;        memory[50314] <=  8'h61;        memory[50315] <=  8'h64;        memory[50316] <=  8'h61;        memory[50317] <=  8'h61;        memory[50318] <=  8'h63;        memory[50319] <=  8'h61;        memory[50320] <=  8'h72;        memory[50321] <=  8'h63;        memory[50322] <=  8'h74;        memory[50323] <=  8'h72;        memory[50324] <=  8'h63;        memory[50325] <=  8'h61;        memory[50326] <=  8'h74;        memory[50327] <=  8'h72;        memory[50328] <=  8'h63;        memory[50329] <=  8'h61;        memory[50330] <=  8'h74;        memory[50331] <=  8'h63;        memory[50332] <=  8'h62;        memory[50333] <=  8'h61;        memory[50334] <=  8'h74;        memory[50335] <=  8'h62;        memory[50336] <=  8'h72;        memory[50337] <=  8'h63;        memory[50338] <=  8'h61;        memory[50339] <=  8'h74;        memory[50340] <=  8'h72;        memory[50341] <=  8'h6e;        memory[50342] <=  8'h62;        memory[50343] <=  8'h61;        memory[50344] <=  8'h63;        memory[50345] <=  8'h61;        memory[50346] <=  8'h74;        memory[50347] <=  8'h79;        memory[50348] <=  8'h73;        memory[50349] <=  8'h6e;        memory[50350] <=  8'h63;        memory[50351] <=  8'h74;        memory[50352] <=  8'h61;        memory[50353] <=  8'h6e;        memory[50354] <=  8'h62;        memory[50355] <=  8'h61;        memory[50356] <=  8'h63;        memory[50357] <=  8'h72;        memory[50358] <=  8'h6e;        memory[50359] <=  8'h74;        memory[50360] <=  8'h61;        memory[50361] <=  8'h62;        memory[50362] <=  8'h74;        memory[50363] <=  8'h6e;        memory[50364] <=  8'h61;        memory[50365] <=  8'h72;        memory[50366] <=  8'h62;        memory[50367] <=  8'h78;        memory[50368] <=  8'h74;        memory[50369] <=  8'h61;        memory[50370] <=  8'h72;        memory[50371] <=  8'h62;        memory[50372] <=  8'h61;        memory[50373] <=  8'h72;        memory[50374] <=  8'h74;        memory[50375] <=  8'h74;        memory[50376] <=  8'h62;        memory[50377] <=  8'h61;        memory[50378] <=  8'h72;        memory[50379] <=  8'h74;        memory[50380] <=  8'h78;        memory[50381] <=  8'h61;        memory[50382] <=  8'h74;        memory[50383] <=  8'h6b;        memory[50384] <=  8'h73;        memory[50385] <=  8'h68;        memory[50386] <=  8'h63;        memory[50387] <=  8'h66;        memory[50388] <=  8'h69;        memory[50389] <=  8'h77;        memory[50390] <=  8'h68;        memory[50391] <=  8'h61;        memory[50392] <=  8'h74;        memory[50393] <=  8'h61;        memory[50394] <=  8'h6e;        memory[50395] <=  8'h61;        memory[50396] <=  8'h62;        memory[50397] <=  8'h61;        memory[50398] <=  8'h63;        memory[50399] <=  8'h61;        memory[50400] <=  8'h74;        memory[50401] <=  8'h61;        memory[50402] <=  8'h62;        memory[50403] <=  8'h61;        memory[50404] <=  8'h72;        memory[50405] <=  8'h63;        memory[50406] <=  8'h61;        memory[50407] <=  8'h68;        memory[50408] <=  8'h64;        memory[50409] <=  8'h75;        memory[50410] <=  8'h63;        memory[50411] <=  8'h74;        memory[50412] <=  8'h61;        memory[50413] <=  8'h64;        memory[50414] <=  8'h61;        memory[50415] <=  8'h61;        memory[50416] <=  8'h63;        memory[50417] <=  8'h61;        memory[50418] <=  8'h72;        memory[50419] <=  8'h63;        memory[50420] <=  8'h74;        memory[50421] <=  8'h72;        memory[50422] <=  8'h63;        memory[50423] <=  8'h61;        memory[50424] <=  8'h74;        memory[50425] <=  8'h72;        memory[50426] <=  8'h63;        memory[50427] <=  8'h61;        memory[50428] <=  8'h74;        memory[50429] <=  8'h63;        memory[50430] <=  8'h62;        memory[50431] <=  8'h61;        memory[50432] <=  8'h74;        memory[50433] <=  8'h62;        memory[50434] <=  8'h72;        memory[50435] <=  8'h63;        memory[50436] <=  8'h61;        memory[50437] <=  8'h74;        memory[50438] <=  8'h72;        memory[50439] <=  8'h6e;        memory[50440] <=  8'h62;        memory[50441] <=  8'h61;        memory[50442] <=  8'h63;        memory[50443] <=  8'h61;        memory[50444] <=  8'h74;        memory[50445] <=  8'h79;        memory[50446] <=  8'h73;        memory[50447] <=  8'h6e;        memory[50448] <=  8'h63;        memory[50449] <=  8'h74;        memory[50450] <=  8'h61;        memory[50451] <=  8'h6e;        memory[50452] <=  8'h62;        memory[50453] <=  8'h61;        memory[50454] <=  8'h63;        memory[50455] <=  8'h72;        memory[50456] <=  8'h6e;        memory[50457] <=  8'h74;        memory[50458] <=  8'h61;        memory[50459] <=  8'h62;        memory[50460] <=  8'h74;        memory[50461] <=  8'h6e;        memory[50462] <=  8'h61;        memory[50463] <=  8'h72;        memory[50464] <=  8'h62;        memory[50465] <=  8'h78;        memory[50466] <=  8'h74;        memory[50467] <=  8'h61;        memory[50468] <=  8'h72;        memory[50469] <=  8'h64;        memory[50470] <=  8'h66;        memory[50471] <=  8'h73;        memory[50472] <=  8'h67;        memory[50473] <=  8'h76;        memory[50474] <=  8'h68;        memory[50475] <=  8'h62;        memory[50476] <=  8'h6b;        memory[50477] <=  8'h6a;        memory[50478] <=  8'h6e;        memory[50479] <=  8'h6d;        memory[50480] <=  8'h62;        memory[50481] <=  8'h76;        memory[50482] <=  8'h78;        memory[50483] <=  8'h63;        memory[50484] <=  8'h73;        memory[50485] <=  8'h66;        memory[50486] <=  8'h72;        memory[50487] <=  8'h74;        memory[50488] <=  8'h79;        memory[50489] <=  8'h75;        memory[50490] <=  8'h6a;        memory[50491] <=  8'h6e;        memory[50492] <=  8'h62;        memory[50493] <=  8'h76;        memory[50494] <=  8'h63;        memory[50495] <=  8'h64;        memory[50496] <=  8'h74;        memory[50497] <=  8'h79;        memory[50498] <=  8'h75;        memory[50499] <=  8'h69;        memory[50500] <=  8'h6b;        memory[50501] <=  8'h6d;        memory[50502] <=  8'h6e;        memory[50503] <=  8'h62;        memory[50504] <=  8'h76;        memory[50505] <=  8'h63;        memory[50506] <=  8'h78;        memory[50507] <=  8'h73;        memory[50508] <=  8'h64;        memory[50509] <=  8'h72;        memory[50510] <=  8'h74;        memory[50511] <=  8'h79;        memory[50512] <=  8'h75;        memory[50513] <=  8'h69;        memory[50514] <=  8'h6b;        memory[50515] <=  8'h6d;        memory[50516] <=  8'h6e;        memory[50517] <=  8'h62;        memory[50518] <=  8'h76;        memory[50519] <=  8'h63;        memory[50520] <=  8'h73;        memory[50521] <=  8'h77;        memory[50522] <=  8'h33;        memory[50523] <=  8'h34;        memory[50524] <=  8'h35;        memory[50525] <=  8'h36;        memory[50526] <=  8'h37;        memory[50527] <=  8'h38;        memory[50528] <=  8'h69;        memory[50529] <=  8'h6b;        memory[50530] <=  8'h6d;        memory[50531] <=  8'h6e;        memory[50532] <=  8'h62;        memory[50533] <=  8'h76;        memory[50534] <=  8'h63;        memory[50535] <=  8'h64;        memory[50536] <=  8'h65;        memory[50537] <=  8'h72;        memory[50538] <=  8'h36;        memory[50539] <=  8'h37;        memory[50540] <=  8'h38;        memory[50541] <=  8'h69;        memory[50542] <=  8'h6f;        memory[50543] <=  8'h6b;        memory[50544] <=  8'h6a;        memory[50545] <=  8'h6e;        memory[50546] <=  8'h62;        memory[50547] <=  8'h76;        memory[50548] <=  8'h63;        memory[50549] <=  8'h64;        memory[50550] <=  8'h72;        memory[50551] <=  8'h74;        memory[50552] <=  8'h79;        memory[50553] <=  8'h75;        memory[50554] <=  8'h73;        memory[50555] <=  8'h6a;        memory[50556] <=  8'h63;        memory[50557] <=  8'h6e;        memory[50558] <=  8'h62;        memory[50559] <=  8'h64;        memory[50560] <=  8'h66;        memory[50561] <=  8'h73;        memory[50562] <=  8'h74;        memory[50563] <=  8'h79;        memory[50564] <=  8'h75;        memory[50565] <=  8'h61;        memory[50566] <=  8'h69;        memory[50567] <=  8'h6b;        memory[50568] <=  8'h78;        memory[50569] <=  8'h6d;        memory[50570] <=  8'h6e;        memory[50571] <=  8'h73;        memory[50572] <=  8'h6a;        memory[50573] <=  8'h6f;        memory[50574] <=  8'h64;        memory[50575] <=  8'h6c;        memory[50576] <=  8'h63;        memory[50577] <=  8'h78;        memory[50578] <=  8'h62;        memory[50579] <=  8'h61;        memory[50580] <=  8'h72;        memory[50581] <=  8'h74;        memory[50582] <=  8'h78;        memory[50583] <=  8'h61;        memory[50584] <=  8'h74;        memory[50585] <=  8'h6b;        memory[50586] <=  8'h73;        memory[50587] <=  8'h68;        memory[50588] <=  8'h63;        memory[50589] <=  8'h66;        memory[50590] <=  8'h69;        memory[50591] <=  8'h77;        memory[50592] <=  8'h68;        memory[50593] <=  8'h61;        memory[50594] <=  8'h74;        memory[50595] <=  8'h61;        memory[50596] <=  8'h6e;        memory[50597] <=  8'h61;        memory[50598] <=  8'h62;        memory[50599] <=  8'h61;        memory[50600] <=  8'h63;        memory[50601] <=  8'h61;        memory[50602] <=  8'h74;        memory[50603] <=  8'h61;        memory[50604] <=  8'h62;        memory[50605] <=  8'h61;        memory[50606] <=  8'h72;        memory[50607] <=  8'h63;        memory[50608] <=  8'h61;        memory[50609] <=  8'h68;        memory[50610] <=  8'h64;        memory[50611] <=  8'h75;        memory[50612] <=  8'h63;        memory[50613] <=  8'h74;        memory[50614] <=  8'h61;        memory[50615] <=  8'h64;        memory[50616] <=  8'h61;        memory[50617] <=  8'h61;        memory[50618] <=  8'h63;        memory[50619] <=  8'h61;        memory[50620] <=  8'h72;        memory[50621] <=  8'h62;        memory[50622] <=  8'h61;        memory[50623] <=  8'h72;        memory[50624] <=  8'h74;        memory[50625] <=  8'h78;        memory[50626] <=  8'h61;        memory[50627] <=  8'h74;        memory[50628] <=  8'h6b;        memory[50629] <=  8'h73;        memory[50630] <=  8'h68;        memory[50631] <=  8'h63;        memory[50632] <=  8'h66;        memory[50633] <=  8'h69;        memory[50634] <=  8'h77;        memory[50635] <=  8'h68;        memory[50636] <=  8'h61;        memory[50637] <=  8'h74;        memory[50638] <=  8'h61;        memory[50639] <=  8'h6e;        memory[50640] <=  8'h61;        memory[50641] <=  8'h62;        memory[50642] <=  8'h61;        memory[50643] <=  8'h63;        memory[50644] <=  8'h61;        memory[50645] <=  8'h74;        memory[50646] <=  8'h61;        memory[50647] <=  8'h62;        memory[50648] <=  8'h61;        memory[50649] <=  8'h72;        memory[50650] <=  8'h63;        memory[50651] <=  8'h61;        memory[50652] <=  8'h68;        memory[50653] <=  8'h64;        memory[50654] <=  8'h75;        memory[50655] <=  8'h63;        memory[50656] <=  8'h74;        memory[50657] <=  8'h61;        memory[50658] <=  8'h64;        memory[50659] <=  8'h61;        memory[50660] <=  8'h61;        memory[50661] <=  8'h63;        memory[50662] <=  8'h61;        memory[50663] <=  8'h72;        memory[50664] <=  8'h62;        memory[50665] <=  8'h61;        memory[50666] <=  8'h72;        memory[50667] <=  8'h74;        memory[50668] <=  8'h78;        memory[50669] <=  8'h61;        memory[50670] <=  8'h74;        memory[50671] <=  8'h6b;        memory[50672] <=  8'h73;        memory[50673] <=  8'h68;        memory[50674] <=  8'h63;        memory[50675] <=  8'h66;        memory[50676] <=  8'h69;        memory[50677] <=  8'h77;        memory[50678] <=  8'h68;        memory[50679] <=  8'h61;        memory[50680] <=  8'h74;        memory[50681] <=  8'h61;        memory[50682] <=  8'h6e;        memory[50683] <=  8'h61;        memory[50684] <=  8'h62;        memory[50685] <=  8'h61;        memory[50686] <=  8'h63;        memory[50687] <=  8'h61;        memory[50688] <=  8'h74;        memory[50689] <=  8'h61;        memory[50690] <=  8'h62;        memory[50691] <=  8'h61;        memory[50692] <=  8'h72;        memory[50693] <=  8'h63;        memory[50694] <=  8'h61;        memory[50695] <=  8'h68;        memory[50696] <=  8'h64;        memory[50697] <=  8'h75;        memory[50698] <=  8'h63;        memory[50699] <=  8'h74;        memory[50700] <=  8'h61;        memory[50701] <=  8'h64;        memory[50702] <=  8'h61;        memory[50703] <=  8'h61;        memory[50704] <=  8'h63;        memory[50705] <=  8'h61;        memory[50706] <=  8'h72;        memory[50707] <=  8'h62;        memory[50708] <=  8'h61;        memory[50709] <=  8'h72;        memory[50710] <=  8'h74;        memory[50711] <=  8'h78;        memory[50712] <=  8'h61;        memory[50713] <=  8'h74;        memory[50714] <=  8'h6b;        memory[50715] <=  8'h73;        memory[50716] <=  8'h68;        memory[50717] <=  8'h63;        memory[50718] <=  8'h66;        memory[50719] <=  8'h69;        memory[50720] <=  8'h77;        memory[50721] <=  8'h68;        memory[50722] <=  8'h61;        memory[50723] <=  8'h74;        memory[50724] <=  8'h61;        memory[50725] <=  8'h6e;        memory[50726] <=  8'h61;        memory[50727] <=  8'h62;        memory[50728] <=  8'h61;        memory[50729] <=  8'h63;        memory[50730] <=  8'h61;        memory[50731] <=  8'h74;        memory[50732] <=  8'h61;        memory[50733] <=  8'h62;        memory[50734] <=  8'h61;        memory[50735] <=  8'h72;        memory[50736] <=  8'h63;        memory[50737] <=  8'h61;        memory[50738] <=  8'h68;        memory[50739] <=  8'h64;        memory[50740] <=  8'h75;        memory[50741] <=  8'h63;        memory[50742] <=  8'h74;        memory[50743] <=  8'h61;        memory[50744] <=  8'h64;        memory[50745] <=  8'h61;        memory[50746] <=  8'h61;        memory[50747] <=  8'h63;        memory[50748] <=  8'h61;        memory[50749] <=  8'h72;        memory[50750] <=  8'h62;        memory[50751] <=  8'h61;        memory[50752] <=  8'h72;        memory[50753] <=  8'h74;        memory[50754] <=  8'h78;        memory[50755] <=  8'h61;        memory[50756] <=  8'h74;        memory[50757] <=  8'h6b;        memory[50758] <=  8'h73;        memory[50759] <=  8'h68;        memory[50760] <=  8'h63;        memory[50761] <=  8'h66;        memory[50762] <=  8'h69;        memory[50763] <=  8'h77;        memory[50764] <=  8'h68;        memory[50765] <=  8'h61;        memory[50766] <=  8'h74;        memory[50767] <=  8'h61;        memory[50768] <=  8'h6e;        memory[50769] <=  8'h61;        memory[50770] <=  8'h62;        memory[50771] <=  8'h61;        memory[50772] <=  8'h63;        memory[50773] <=  8'h61;        memory[50774] <=  8'h74;        memory[50775] <=  8'h61;        memory[50776] <=  8'h62;        memory[50777] <=  8'h61;        memory[50778] <=  8'h72;        memory[50779] <=  8'h63;        memory[50780] <=  8'h61;        memory[50781] <=  8'h68;        memory[50782] <=  8'h64;        memory[50783] <=  8'h75;        memory[50784] <=  8'h63;        memory[50785] <=  8'h74;        memory[50786] <=  8'h61;        memory[50787] <=  8'h64;        memory[50788] <=  8'h61;        memory[50789] <=  8'h61;        memory[50790] <=  8'h63;        memory[50791] <=  8'h61;        memory[50792] <=  8'h72;        memory[50793] <=  8'h62;        memory[50794] <=  8'h61;        memory[50795] <=  8'h72;        memory[50796] <=  8'h74;        memory[50797] <=  8'h78;        memory[50798] <=  8'h61;        memory[50799] <=  8'h74;        memory[50800] <=  8'h6b;        memory[50801] <=  8'h73;        memory[50802] <=  8'h68;        memory[50803] <=  8'h63;        memory[50804] <=  8'h66;        memory[50805] <=  8'h69;        memory[50806] <=  8'h77;        memory[50807] <=  8'h68;        memory[50808] <=  8'h61;        memory[50809] <=  8'h74;        memory[50810] <=  8'h61;        memory[50811] <=  8'h6e;        memory[50812] <=  8'h61;        memory[50813] <=  8'h62;        memory[50814] <=  8'h61;        memory[50815] <=  8'h63;        memory[50816] <=  8'h61;        memory[50817] <=  8'h74;        memory[50818] <=  8'h61;        memory[50819] <=  8'h62;        memory[50820] <=  8'h61;        memory[50821] <=  8'h72;        memory[50822] <=  8'h63;        memory[50823] <=  8'h61;        memory[50824] <=  8'h68;        memory[50825] <=  8'h64;        memory[50826] <=  8'h75;        memory[50827] <=  8'h63;        memory[50828] <=  8'h74;        memory[50829] <=  8'h61;        memory[50830] <=  8'h64;        memory[50831] <=  8'h61;        memory[50832] <=  8'h61;        memory[50833] <=  8'h63;        memory[50834] <=  8'h61;        memory[50835] <=  8'h72;        memory[50836] <=  8'h62;        memory[50837] <=  8'h61;        memory[50838] <=  8'h72;        memory[50839] <=  8'h74;        memory[50840] <=  8'h78;        memory[50841] <=  8'h61;        memory[50842] <=  8'h74;        memory[50843] <=  8'h6b;        memory[50844] <=  8'h73;        memory[50845] <=  8'h68;        memory[50846] <=  8'h63;        memory[50847] <=  8'h66;        memory[50848] <=  8'h69;        memory[50849] <=  8'h77;        memory[50850] <=  8'h68;        memory[50851] <=  8'h61;        memory[50852] <=  8'h74;        memory[50853] <=  8'h61;        memory[50854] <=  8'h6e;        memory[50855] <=  8'h61;        memory[50856] <=  8'h62;        memory[50857] <=  8'h61;        memory[50858] <=  8'h63;        memory[50859] <=  8'h61;        memory[50860] <=  8'h74;        memory[50861] <=  8'h61;        memory[50862] <=  8'h62;        memory[50863] <=  8'h61;        memory[50864] <=  8'h72;        memory[50865] <=  8'h63;        memory[50866] <=  8'h61;        memory[50867] <=  8'h68;        memory[50868] <=  8'h64;        memory[50869] <=  8'h75;        memory[50870] <=  8'h63;        memory[50871] <=  8'h74;        memory[50872] <=  8'h61;        memory[50873] <=  8'h64;        memory[50874] <=  8'h61;        memory[50875] <=  8'h61;        memory[50876] <=  8'h63;        memory[50877] <=  8'h61;        memory[50878] <=  8'h72;        memory[50879] <=  8'h62;        memory[50880] <=  8'h61;        memory[50881] <=  8'h72;        memory[50882] <=  8'h74;        memory[50883] <=  8'h78;        memory[50884] <=  8'h61;        memory[50885] <=  8'h74;        memory[50886] <=  8'h6b;        memory[50887] <=  8'h73;        memory[50888] <=  8'h68;        memory[50889] <=  8'h63;        memory[50890] <=  8'h66;        memory[50891] <=  8'h69;        memory[50892] <=  8'h77;        memory[50893] <=  8'h68;        memory[50894] <=  8'h61;        memory[50895] <=  8'h74;        memory[50896] <=  8'h61;        memory[50897] <=  8'h6e;        memory[50898] <=  8'h61;        memory[50899] <=  8'h62;        memory[50900] <=  8'h61;        memory[50901] <=  8'h63;        memory[50902] <=  8'h61;        memory[50903] <=  8'h74;        memory[50904] <=  8'h61;        memory[50905] <=  8'h62;        memory[50906] <=  8'h61;        memory[50907] <=  8'h72;        memory[50908] <=  8'h63;        memory[50909] <=  8'h61;        memory[50910] <=  8'h68;        memory[50911] <=  8'h64;        memory[50912] <=  8'h75;        memory[50913] <=  8'h63;        memory[50914] <=  8'h74;        memory[50915] <=  8'h61;        memory[50916] <=  8'h64;        memory[50917] <=  8'h61;        memory[50918] <=  8'h61;        memory[50919] <=  8'h63;        memory[50920] <=  8'h61;        memory[50921] <=  8'h72;        memory[50922] <=  8'h62;        memory[50923] <=  8'h61;        memory[50924] <=  8'h72;        memory[50925] <=  8'h74;        memory[50926] <=  8'h78;        memory[50927] <=  8'h61;        memory[50928] <=  8'h74;        memory[50929] <=  8'h6b;        memory[50930] <=  8'h73;        memory[50931] <=  8'h68;        memory[50932] <=  8'h63;        memory[50933] <=  8'h66;        memory[50934] <=  8'h69;        memory[50935] <=  8'h77;        memory[50936] <=  8'h68;        memory[50937] <=  8'h61;        memory[50938] <=  8'h74;        memory[50939] <=  8'h61;        memory[50940] <=  8'h6e;        memory[50941] <=  8'h61;        memory[50942] <=  8'h62;        memory[50943] <=  8'h61;        memory[50944] <=  8'h63;        memory[50945] <=  8'h61;        memory[50946] <=  8'h74;        memory[50947] <=  8'h61;        memory[50948] <=  8'h62;        memory[50949] <=  8'h61;        memory[50950] <=  8'h72;        memory[50951] <=  8'h63;        memory[50952] <=  8'h61;        memory[50953] <=  8'h68;        memory[50954] <=  8'h64;        memory[50955] <=  8'h75;        memory[50956] <=  8'h63;        memory[50957] <=  8'h74;        memory[50958] <=  8'h61;        memory[50959] <=  8'h64;        memory[50960] <=  8'h61;        memory[50961] <=  8'h61;        memory[50962] <=  8'h63;        memory[50963] <=  8'h61;        memory[50964] <=  8'h72;        memory[50965] <=  8'h62;        memory[50966] <=  8'h61;        memory[50967] <=  8'h72;        memory[50968] <=  8'h74;        memory[50969] <=  8'h74;        memory[50970] <=  8'h62;        memory[50971] <=  8'h61;        memory[50972] <=  8'h72;        memory[50973] <=  8'h74;        memory[50974] <=  8'h78;        memory[50975] <=  8'h61;        memory[50976] <=  8'h74;        memory[50977] <=  8'h6b;        memory[50978] <=  8'h73;        memory[50979] <=  8'h68;        memory[50980] <=  8'h63;        memory[50981] <=  8'h66;        memory[50982] <=  8'h69;        memory[50983] <=  8'h77;        memory[50984] <=  8'h68;        memory[50985] <=  8'h61;        memory[50986] <=  8'h74;        memory[50987] <=  8'h61;        memory[50988] <=  8'h6e;        memory[50989] <=  8'h61;        memory[50990] <=  8'h62;        memory[50991] <=  8'h61;        memory[50992] <=  8'h63;        memory[50993] <=  8'h61;        memory[50994] <=  8'h74;        memory[50995] <=  8'h61;        memory[50996] <=  8'h62;        memory[50997] <=  8'h61;        memory[50998] <=  8'h72;        memory[50999] <=  8'h63;        memory[51000] <=  8'h61;        memory[51001] <=  8'h68;        memory[51002] <=  8'h64;        memory[51003] <=  8'h75;        memory[51004] <=  8'h63;        memory[51005] <=  8'h74;        memory[51006] <=  8'h61;        memory[51007] <=  8'h64;        memory[51008] <=  8'h61;        memory[51009] <=  8'h61;        memory[51010] <=  8'h63;        memory[51011] <=  8'h61;        memory[51012] <=  8'h72;        memory[51013] <=  8'h63;        memory[51014] <=  8'h74;        memory[51015] <=  8'h72;        memory[51016] <=  8'h63;        memory[51017] <=  8'h61;        memory[51018] <=  8'h74;        memory[51019] <=  8'h72;        memory[51020] <=  8'h63;        memory[51021] <=  8'h61;        memory[51022] <=  8'h74;        memory[51023] <=  8'h63;        memory[51024] <=  8'h62;        memory[51025] <=  8'h61;        memory[51026] <=  8'h74;        memory[51027] <=  8'h62;        memory[51028] <=  8'h72;        memory[51029] <=  8'h63;        memory[51030] <=  8'h61;        memory[51031] <=  8'h72;        memory[51032] <=  8'h62;        memory[51033] <=  8'h78;        memory[51034] <=  8'h74;        memory[51035] <=  8'h61;        memory[51036] <=  8'h72;        memory[51037] <=  8'h64;        memory[51038] <=  8'h66;        memory[51039] <=  8'h73;        memory[51040] <=  8'h67;        memory[51041] <=  8'h76;        memory[51042] <=  8'h68;        memory[51043] <=  8'h62;        memory[51044] <=  8'h6b;        memory[51045] <=  8'h6a;        memory[51046] <=  8'h6e;        memory[51047] <=  8'h6d;        memory[51048] <=  8'h62;        memory[51049] <=  8'h76;        memory[51050] <=  8'h78;        memory[51051] <=  8'h63;        memory[51052] <=  8'h73;        memory[51053] <=  8'h66;        memory[51054] <=  8'h72;        memory[51055] <=  8'h74;        memory[51056] <=  8'h79;        memory[51057] <=  8'h75;        memory[51058] <=  8'h6a;        memory[51059] <=  8'h6e;        memory[51060] <=  8'h62;        memory[51061] <=  8'h76;        memory[51062] <=  8'h63;        memory[51063] <=  8'h64;        memory[51064] <=  8'h74;        memory[51065] <=  8'h79;        memory[51066] <=  8'h75;        memory[51067] <=  8'h69;        memory[51068] <=  8'h6b;        memory[51069] <=  8'h6d;        memory[51070] <=  8'h6e;        memory[51071] <=  8'h62;        memory[51072] <=  8'h76;        memory[51073] <=  8'h63;        memory[51074] <=  8'h78;        memory[51075] <=  8'h73;        memory[51076] <=  8'h64;        memory[51077] <=  8'h72;        memory[51078] <=  8'h74;        memory[51079] <=  8'h79;        memory[51080] <=  8'h75;        memory[51081] <=  8'h69;        memory[51082] <=  8'h6b;        memory[51083] <=  8'h6d;        memory[51084] <=  8'h6e;        memory[51085] <=  8'h62;        memory[51086] <=  8'h76;        memory[51087] <=  8'h63;        memory[51088] <=  8'h73;        memory[51089] <=  8'h77;        memory[51090] <=  8'h33;        memory[51091] <=  8'h34;        memory[51092] <=  8'h35;        memory[51093] <=  8'h36;        memory[51094] <=  8'h37;        memory[51095] <=  8'h38;        memory[51096] <=  8'h69;        memory[51097] <=  8'h6b;        memory[51098] <=  8'h6d;        memory[51099] <=  8'h6e;        memory[51100] <=  8'h62;        memory[51101] <=  8'h76;        memory[51102] <=  8'h63;        memory[51103] <=  8'h64;        memory[51104] <=  8'h65;        memory[51105] <=  8'h72;        memory[51106] <=  8'h36;        memory[51107] <=  8'h37;        memory[51108] <=  8'h38;        memory[51109] <=  8'h69;        memory[51110] <=  8'h6f;        memory[51111] <=  8'h6b;        memory[51112] <=  8'h6a;        memory[51113] <=  8'h6e;        memory[51114] <=  8'h62;        memory[51115] <=  8'h76;        memory[51116] <=  8'h63;        memory[51117] <=  8'h64;        memory[51118] <=  8'h72;        memory[51119] <=  8'h74;        memory[51120] <=  8'h79;        memory[51121] <=  8'h75;        memory[51122] <=  8'h73;        memory[51123] <=  8'h6a;        memory[51124] <=  8'h63;        memory[51125] <=  8'h6e;        memory[51126] <=  8'h62;        memory[51127] <=  8'h64;        memory[51128] <=  8'h66;        memory[51129] <=  8'h73;        memory[51130] <=  8'h74;        memory[51131] <=  8'h79;        memory[51132] <=  8'h75;        memory[51133] <=  8'h61;        memory[51134] <=  8'h69;        memory[51135] <=  8'h6b;        memory[51136] <=  8'h78;        memory[51137] <=  8'h6d;        memory[51138] <=  8'h6e;        memory[51139] <=  8'h73;        memory[51140] <=  8'h6a;        memory[51141] <=  8'h6f;        memory[51142] <=  8'h64;        memory[51143] <=  8'h6c;        memory[51144] <=  8'h63;        memory[51145] <=  8'h78;        memory[51146] <=  8'h2c;        memory[51147] <=  8'h6d;        memory[51148] <=  8'h73;        memory[51149] <=  8'h6b;        memory[51150] <=  8'h64;        memory[51151] <=  8'h6c;        memory[51152] <=  8'h70;        memory[51153] <=  8'h5b;        memory[51154] <=  8'h3b;        memory[51155] <=  8'h73;        memory[51156] <=  8'h6c;        memory[51157] <=  8'h64;        memory[51158] <=  8'h70;        memory[51159] <=  8'h76;        memory[51160] <=  8'h63;        memory[51161] <=  8'h5b;        memory[51162] <=  8'h78;        memory[51163] <=  8'h76;        memory[51164] <=  8'h63;        memory[51165] <=  8'h5b;        memory[51166] <=  8'h78;        memory[51167] <=  8'h70;        memory[51168] <=  8'h6f;        memory[51169] <=  8'h20;        memory[51170] <=  8'h62;        memory[51171] <=  8'h61;        memory[51172] <=  8'h72;        memory[51173] <=  8'h74;        memory[51174] <=  8'h74;        memory[51175] <=  8'h62;        memory[51176] <=  8'h61;        memory[51177] <=  8'h72;        memory[51178] <=  8'h74;        memory[51179] <=  8'h78;        memory[51180] <=  8'h61;        memory[51181] <=  8'h74;        memory[51182] <=  8'h6b;        memory[51183] <=  8'h73;        memory[51184] <=  8'h68;        memory[51185] <=  8'h63;        memory[51186] <=  8'h66;        memory[51187] <=  8'h69;        memory[51188] <=  8'h77;        memory[51189] <=  8'h68;        memory[51190] <=  8'h61;        memory[51191] <=  8'h69;        memory[51192] <=  8'h6a;        memory[51193] <=  8'h78;        memory[51194] <=  8'h5d;        memory[51195] <=  8'h65;        memory[51196] <=  8'h6b;        memory[51197] <=  8'h6f;        memory[51198] <=  8'h39;        memory[51199] <=  8'h64;        memory[51200] <=  8'h75;        memory[51201] <=  8'h38;        memory[51202] <=  8'h79;        memory[51203] <=  8'h20;        memory[51204] <=  8'h37;        memory[51205] <=  8'h63;        memory[51206] <=  8'h67;        memory[51207] <=  8'h78;        memory[51208] <=  8'h63;        memory[51209] <=  8'h75;        memory[51210] <=  8'h68;        memory[51211] <=  8'h69;        memory[51212] <=  8'h6a;        memory[51213] <=  8'h77;        memory[51214] <=  8'h69;        memory[51215] <=  8'h64;        memory[51216] <=  8'h66;        memory[51217] <=  8'h68;        memory[51218] <=  8'h75;        memory[51219] <=  8'h76;        memory[51220] <=  8'h64;        memory[51221] <=  8'h62;        memory[51222] <=  8'h66;        memory[51223] <=  8'h6a;        memory[51224] <=  8'h6e;        memory[51225] <=  8'h6b;        memory[51226] <=  8'h6a;        memory[51227] <=  8'h65;        memory[51228] <=  8'h38;        memory[51229] <=  8'h66;        memory[51230] <=  8'h37;        memory[51231] <=  8'h67;        memory[51232] <=  8'h79;        memory[51233] <=  8'h76;        memory[51234] <=  8'h63;        memory[51235] <=  8'h68;        memory[51236] <=  8'h69;        memory[51237] <=  8'h6a;        memory[51238] <=  8'h33;        memory[51239] <=  8'h65;        memory[51240] <=  8'h67;        memory[51241] <=  8'h79;        memory[51242] <=  8'h72;        memory[51243] <=  8'h64;        memory[51244] <=  8'h62;        memory[51245] <=  8'h6e;        memory[51246] <=  8'h63;        memory[51247] <=  8'h7a;        memory[51248] <=  8'h6a;        memory[51249] <=  8'h6f;        memory[51250] <=  8'h66;        memory[51251] <=  8'h78;        memory[51252] <=  8'h6a;        memory[51253] <=  8'h69;        memory[51254] <=  8'h63;        memory[51255] <=  8'h68;        memory[51256] <=  8'h62;        memory[51257] <=  8'h6e;        memory[51258] <=  8'h6d;        memory[51259] <=  8'h63;        memory[51260] <=  8'h73;        memory[51261] <=  8'h6c;        memory[51262] <=  8'h6b;        memory[51263] <=  8'h6a;        memory[51264] <=  8'h69;        memory[51265] <=  8'h68;        memory[51266] <=  8'h76;        memory[51267] <=  8'h75;        memory[51268] <=  8'h69;        memory[51269] <=  8'h64;        memory[51270] <=  8'h68;        memory[51271] <=  8'h75;        memory[51272] <=  8'h67;        memory[51273] <=  8'h79;        memory[51274] <=  8'h62;        memory[51275] <=  8'h68;        memory[51276] <=  8'h65;        memory[51277] <=  8'h6a;        memory[51278] <=  8'h72;        memory[51279] <=  8'h6b;        memory[51280] <=  8'h6a;        memory[51281] <=  8'h6f;        memory[51282] <=  8'h64;        memory[51283] <=  8'h67;        memory[51284] <=  8'h69;        memory[51285] <=  8'h75;        memory[51286] <=  8'h69;        memory[51287] <=  8'h67;        memory[51288] <=  8'h76;        memory[51289] <=  8'h79;        memory[51290] <=  8'h75;        memory[51291] <=  8'h67;        memory[51292] <=  8'h78;        memory[51293] <=  8'h68;        memory[51294] <=  8'h63;        memory[51295] <=  8'h20;        memory[51296] <=  8'h20;        memory[51297] <=  8'h20;        memory[51298] <=  8'h78;        memory[51299] <=  8'h76;        memory[51300] <=  8'h20;        memory[51301] <=  8'h63;        memory[51302] <=  8'h78;        memory[51303] <=  8'h67;        memory[51304] <=  8'h79;        memory[51305] <=  8'h63;        memory[51306] <=  8'h75;        memory[51307] <=  8'h68;        memory[51308] <=  8'h6a;        memory[51309] <=  8'h6b;        memory[51310] <=  8'h61;        memory[51311] <=  8'h6c;        memory[51312] <=  8'h78;        memory[51313] <=  8'h76;        memory[51314] <=  8'h70;        memory[51315] <=  8'h6f;        memory[51316] <=  8'h69;        memory[51317] <=  8'h6a;        memory[51318] <=  8'h69;        memory[51319] <=  8'h68;        memory[51320] <=  8'h6a;        memory[51321] <=  8'h62;        memory[51322] <=  8'h77;        memory[51323] <=  8'h65;        memory[51324] <=  8'h6e;        memory[51325] <=  8'h61;        memory[51326] <=  8'h66;        memory[51327] <=  8'h6d;        memory[51328] <=  8'h64;        memory[51329] <=  8'h6b;        memory[51330] <=  8'h6d;        memory[51331] <=  8'h76;        memory[51332] <=  8'h6c;        memory[51333] <=  8'h63;        memory[51334] <=  8'h6f;        memory[51335] <=  8'h64;        memory[51336] <=  8'h69;        memory[51337] <=  8'h75;        memory[51338] <=  8'h68;        memory[51339] <=  8'h73;        memory[51340] <=  8'h66;        memory[51341] <=  8'h65;        memory[51342] <=  8'h62;        memory[51343] <=  8'h6e;        memory[51344] <=  8'h64;        memory[51345] <=  8'h73;        memory[51346] <=  8'h63;        memory[51347] <=  8'h6b;        memory[51348] <=  8'h20;        memory[51349] <=  8'h78;        memory[51350] <=  8'h6a;        memory[51351] <=  8'h78;        memory[51352] <=  8'h63;        memory[51353] <=  8'h73;        memory[51354] <=  8'h64;        memory[51355] <=  8'h66;        memory[51356] <=  8'h6b;        memory[51357] <=  8'h64;        memory[51358] <=  8'h6e;        memory[51359] <=  8'h6d;        memory[51360] <=  8'h64;        memory[51361] <=  8'h73;        memory[51362] <=  8'h63;        memory[51363] <=  8'h6b;        memory[51364] <=  8'h78;        memory[51365] <=  8'h6c;        memory[51366] <=  8'h6f;        memory[51367] <=  8'h66;        memory[51368] <=  8'h6a;        memory[51369] <=  8'h69;        memory[51370] <=  8'h61;        memory[51371] <=  8'h62;        memory[51372] <=  8'h6e;        memory[51373] <=  8'h20;        memory[51374] <=  8'h78;        memory[51375] <=  8'h6b;        memory[51376] <=  8'h6d;        memory[51377] <=  8'h20;        memory[51378] <=  8'h6f;        memory[51379] <=  8'h63;        memory[51380] <=  8'h76;        memory[51381] <=  8'h73;        memory[51382] <=  8'h64;        memory[51383] <=  8'h69;        memory[51384] <=  8'h66;        memory[51385] <=  8'h68;        memory[51386] <=  8'h65;        memory[51387] <=  8'h71;        memory[51388] <=  8'h6a;        memory[51389] <=  8'h77;        memory[51390] <=  8'h62;        memory[51391] <=  8'h65;        memory[51392] <=  8'h6e;        memory[51393] <=  8'h20;        memory[51394] <=  8'h6d;        memory[51395] <=  8'h64;        memory[51396] <=  8'h73;        memory[51397] <=  8'h6c;        memory[51398] <=  8'h76;        memory[51399] <=  8'h6b;        memory[51400] <=  8'h63;        memory[51401] <=  8'h78;        memory[51402] <=  8'h20;        memory[51403] <=  8'h6f;        memory[51404] <=  8'h78;        memory[51405] <=  8'h69;        memory[51406] <=  8'h63;        memory[51407] <=  8'h6a;        memory[51408] <=  8'h76;        memory[51409] <=  8'h64;        memory[51410] <=  8'h66;        memory[51411] <=  8'h65;        memory[51412] <=  8'h71;        memory[51413] <=  8'h6e;        memory[51414] <=  8'h20;        memory[51415] <=  8'h64;        memory[51416] <=  8'h6d;        memory[51417] <=  8'h73;        memory[51418] <=  8'h6c;        memory[51419] <=  8'h63;        memory[51420] <=  8'h78;        memory[51421] <=  8'h6b;        memory[51422] <=  8'h20;        memory[51423] <=  8'h6f;        memory[51424] <=  8'h78;        memory[51425] <=  8'h63;        memory[51426] <=  8'h76;        memory[51427] <=  8'h6a;        memory[51428] <=  8'h64;        memory[51429] <=  8'h62;        memory[51430] <=  8'h71;        memory[51431] <=  8'h77;        memory[51432] <=  8'h65;        memory[51433] <=  8'h6e;        memory[51434] <=  8'h6d;        memory[51435] <=  8'h64;        memory[51436] <=  8'h6c;        memory[51437] <=  8'h73;        memory[51438] <=  8'h2c;        memory[51439] <=  8'h76;        memory[51440] <=  8'h63;        memory[51441] <=  8'h78;        memory[51442] <=  8'h20;        memory[51443] <=  8'h63;        memory[51444] <=  8'h6f;        memory[51445] <=  8'h69;        memory[51446] <=  8'h76;        memory[51447] <=  8'h68;        memory[51448] <=  8'h73;        memory[51449] <=  8'h64;        memory[51450] <=  8'h62;        memory[51451] <=  8'h71;        memory[51452] <=  8'h77;        memory[51453] <=  8'h65;        memory[51454] <=  8'h6e;        memory[51455] <=  8'h64;        memory[51456] <=  8'h6b;        memory[51457] <=  8'h73;        memory[51458] <=  8'h76;        memory[51459] <=  8'h6f;        memory[51460] <=  8'h63;        memory[51461] <=  8'h20;        memory[51462] <=  8'h76;        memory[51463] <=  8'h69;        memory[51464] <=  8'h75;        memory[51465] <=  8'h69;        memory[51466] <=  8'h68;        memory[51467] <=  8'h63;        memory[51468] <=  8'h78;        memory[51469] <=  8'h69;        memory[51470] <=  8'h6f;        memory[51471] <=  8'h76;        memory[51472] <=  8'h73;        memory[51473] <=  8'h64;        memory[51474] <=  8'h61;        memory[51475] <=  8'h64;        memory[51476] <=  8'h6e;        memory[51477] <=  8'h77;        memory[51478] <=  8'h71;        memory[51479] <=  8'h6b;        memory[51480] <=  8'h6c;        memory[51481] <=  8'h73;        memory[51482] <=  8'h76;        memory[51483] <=  8'h6e;        memory[51484] <=  8'h62;        memory[51485] <=  8'h20;        memory[51486] <=  8'h64;        memory[51487] <=  8'h66;        memory[51488] <=  8'h6a;        memory[51489] <=  8'h6b;        memory[51490] <=  8'h71;        memory[51491] <=  8'h64;        memory[51492] <=  8'h77;        memory[51493] <=  8'h65;        memory[51494] <=  8'h6e;        memory[51495] <=  8'h62;        memory[51496] <=  8'h20;        memory[51497] <=  8'h64;        memory[51498] <=  8'h73;        memory[51499] <=  8'h76;        memory[51500] <=  8'h68;        memory[51501] <=  8'h64;        memory[51502] <=  8'h61;        memory[51503] <=  8'h71;        memory[51504] <=  8'h77;        memory[51505] <=  8'h6a;        memory[51506] <=  8'h65;        memory[51507] <=  8'h6e;        memory[51508] <=  8'h64;        memory[51509] <=  8'h20;        memory[51510] <=  8'h61;        memory[51511] <=  8'h63;        memory[51512] <=  8'h62;        memory[51513] <=  8'h68;        memory[51514] <=  8'h64;        memory[51515] <=  8'h61;        memory[51516] <=  8'h77;        memory[51517] <=  8'h71;        memory[51518] <=  8'h6e;        memory[51519] <=  8'h20;        memory[51520] <=  8'h62;        memory[51521] <=  8'h73;        memory[51522] <=  8'h76;        memory[51523] <=  8'h61;        memory[51524] <=  8'h67;        memory[51525] <=  8'h76;        memory[51526] <=  8'h68;        memory[51527] <=  8'h67;        memory[51528] <=  8'h61;        memory[51529] <=  8'h73;        memory[51530] <=  8'h6a;        memory[51531] <=  8'h6b;        memory[51532] <=  8'h63;        memory[51533] <=  8'h78;        memory[51534] <=  8'h76;        memory[51535] <=  8'h6e;        memory[51536] <=  8'h73;        memory[51537] <=  8'h64;        memory[51538] <=  8'h20;        memory[51539] <=  8'h66;        memory[51540] <=  8'h62;        memory[51541] <=  8'h64;        memory[51542] <=  8'h61;        memory[51543] <=  8'h73;        memory[51544] <=  8'h76;        memory[51545] <=  8'h67;        memory[51546] <=  8'h63;        memory[51547] <=  8'h79;        memory[51548] <=  8'h7a;        memory[51549] <=  8'h78;        memory[51550] <=  8'h79;        memory[51551] <=  8'h75;        memory[51552] <=  8'h20;        memory[51553] <=  8'h69;        memory[51554] <=  8'h6a;        memory[51555] <=  8'h64;        memory[51556] <=  8'h66;        memory[51557] <=  8'h6b;        memory[51558] <=  8'h61;        memory[51559] <=  8'h64;        memory[51560] <=  8'h63;        memory[51561] <=  8'h78;        memory[51562] <=  8'h68;        memory[51563] <=  8'h20;        memory[51564] <=  8'h67;        memory[51565] <=  8'h61;        memory[51566] <=  8'h68;        memory[51567] <=  8'h75;        memory[51568] <=  8'h64;        memory[51569] <=  8'h73;        memory[51570] <=  8'h69;        memory[51571] <=  8'h6a;        memory[51572] <=  8'h61;        memory[51573] <=  8'h6b;        memory[51574] <=  8'h63;        memory[51575] <=  8'h62;        memory[51576] <=  8'h61;        memory[51577] <=  8'h72;        memory[51578] <=  8'h73;        memory[51579] <=  8'h68;        memory[51580] <=  8'h64;        memory[51581] <=  8'h66;        memory[51582] <=  8'h67;        memory[51583] <=  8'h73;        memory[51584] <=  8'h68;        memory[51585] <=  8'h64;        memory[51586] <=  8'h66;        memory[51587] <=  8'h68;        memory[51588] <=  8'h64;        memory[51589] <=  8'h6a;        memory[51590] <=  8'h68;        memory[51591] <=  8'h62;        memory[51592] <=  8'h67;        memory[51593] <=  8'h63;        memory[51594] <=  8'h61;        memory[51595] <=  8'h66;        memory[51596] <=  8'h73;        memory[51597] <=  8'h79;        memory[51598] <=  8'h67;        memory[51599] <=  8'h6b;        memory[51600] <=  8'h75;        memory[51601] <=  8'h64;        memory[51602] <=  8'h68;        memory[51603] <=  8'h62;        memory[51604] <=  8'h77;        memory[51605] <=  8'h76;        memory[51606] <=  8'h67;        memory[51607] <=  8'h61;        memory[51608] <=  8'h66;        memory[51609] <=  8'h64;        memory[51610] <=  8'h74;        memory[51611] <=  8'h75;        memory[51612] <=  8'h66;        memory[51613] <=  8'h79;        memory[51614] <=  8'h67;        memory[51615] <=  8'h69;        memory[51616] <=  8'h75;        memory[51617] <=  8'h68;        memory[51618] <=  8'h6c;        memory[51619] <=  8'h6a;        memory[51620] <=  8'h62;        memory[51621] <=  8'h6b;        memory[51622] <=  8'h68;        memory[51623] <=  8'h76;        memory[51624] <=  8'h67;        memory[51625] <=  8'h63;        memory[51626] <=  8'h66;        memory[51627] <=  8'h78;        memory[51628] <=  8'h64;        memory[51629] <=  8'h74;        memory[51630] <=  8'h75;        memory[51631] <=  8'h79;        memory[51632] <=  8'h69;        memory[51633] <=  8'h75;        memory[51634] <=  8'h68;        memory[51635] <=  8'h6c;        memory[51636] <=  8'h6a;        memory[51637] <=  8'h6b;        memory[51638] <=  8'h67;        memory[51639] <=  8'h6a;        memory[51640] <=  8'h63;        memory[51641] <=  8'h66;        memory[51642] <=  8'h68;        memory[51643] <=  8'h64;        memory[51644] <=  8'h67;        memory[51645] <=  8'h72;        memory[51646] <=  8'h79;        memory[51647] <=  8'h74;        memory[51648] <=  8'h66;        memory[51649] <=  8'h75;        memory[51650] <=  8'h79;        memory[51651] <=  8'h69;        memory[51652] <=  8'h68;        memory[51653] <=  8'h6c;        memory[51654] <=  8'h62;        memory[51655] <=  8'h6d;        memory[51656] <=  8'h76;        memory[51657] <=  8'h6e;        memory[51658] <=  8'h63;        memory[51659] <=  8'h66;        memory[51660] <=  8'h68;        memory[51661] <=  8'h64;        memory[51662] <=  8'h74;        memory[51663] <=  8'h75;        memory[51664] <=  8'h67;        memory[51665] <=  8'h79;        memory[51666] <=  8'h69;        memory[51667] <=  8'h68;        memory[51668] <=  8'h75;        memory[51669] <=  8'h6a;        memory[51670] <=  8'h6c;        memory[51671] <=  8'h62;        memory[51672] <=  8'h6d;        memory[51673] <=  8'h76;        memory[51674] <=  8'h6e;        memory[51675] <=  8'h63;        memory[51676] <=  8'h66;        memory[51677] <=  8'h68;        memory[51678] <=  8'h67;        memory[51679] <=  8'h79;        memory[51680] <=  8'h68;        memory[51681] <=  8'h75;        memory[51682] <=  8'h6a;        memory[51683] <=  8'h6e;        memory[51684] <=  8'h2c;        memory[51685] <=  8'h62;        memory[51686] <=  8'h6e;        memory[51687] <=  8'h6d;        memory[51688] <=  8'h76;        memory[51689] <=  8'h6e;        memory[51690] <=  8'h63;        memory[51691] <=  8'h66;        memory[51692] <=  8'h68;        memory[51693] <=  8'h74;        memory[51694] <=  8'h79;        memory[51695] <=  8'h69;        memory[51696] <=  8'h75;        memory[51697] <=  8'h6c;        memory[51698] <=  8'h6a;        memory[51699] <=  8'h62;        memory[51700] <=  8'h6d;        memory[51701] <=  8'h76;        memory[51702] <=  8'h6e;        memory[51703] <=  8'h63;        memory[51704] <=  8'h66;        memory[51705] <=  8'h74;        memory[51706] <=  8'h75;        memory[51707] <=  8'h79;        memory[51708] <=  8'h69;        memory[51709] <=  8'h68;        memory[51710] <=  8'h6b;        memory[51711] <=  8'h62;        memory[51712] <=  8'h76;        memory[51713] <=  8'h63;        memory[51714] <=  8'h66;        memory[51715] <=  8'h67;        memory[51716] <=  8'h74;        memory[51717] <=  8'h75;        memory[51718] <=  8'h79;        memory[51719] <=  8'h69;        memory[51720] <=  8'h75;        memory[51721] <=  8'h68;        memory[51722] <=  8'h6a;        memory[51723] <=  8'h6b;        memory[51724] <=  8'h62;        memory[51725] <=  8'h76;        memory[51726] <=  8'h63;        memory[51727] <=  8'h66;        memory[51728] <=  8'h74;        memory[51729] <=  8'h75;        memory[51730] <=  8'h79;        memory[51731] <=  8'h69;        memory[51732] <=  8'h75;        memory[51733] <=  8'h6a;        memory[51734] <=  8'h6b;        memory[51735] <=  8'h6e;        memory[51736] <=  8'h62;        memory[51737] <=  8'h76;        memory[51738] <=  8'h67;        memory[51739] <=  8'h66;        memory[51740] <=  8'h74;        memory[51741] <=  8'h79;        memory[51742] <=  8'h75;        memory[51743] <=  8'h75;        memory[51744] <=  8'h69;        memory[51745] <=  8'h6a;        memory[51746] <=  8'h6b;        memory[51747] <=  8'h68;        memory[51748] <=  8'h62;        memory[51749] <=  8'h6a;        memory[51750] <=  8'h67;        memory[51751] <=  8'h68;        memory[51752] <=  8'h66;        memory[51753] <=  8'h79;        memory[51754] <=  8'h74;        memory[51755] <=  8'h79;        memory[51756] <=  8'h69;        memory[51757] <=  8'h75;        memory[51758] <=  8'h64;        memory[51759] <=  8'h6a;        memory[51760] <=  8'h6b;        memory[51761] <=  8'h68;        memory[51762] <=  8'h63;        memory[51763] <=  8'h7a;        memory[51764] <=  8'h67;        memory[51765] <=  8'h68;        memory[51766] <=  8'h74;        memory[51767] <=  8'h75;        memory[51768] <=  8'h79;        memory[51769] <=  8'h69;        memory[51770] <=  8'h61;        memory[51771] <=  8'h73;        memory[51772] <=  8'h75;        memory[51773] <=  8'h6a;        memory[51774] <=  8'h6b;        memory[51775] <=  8'h62;        memory[51776] <=  8'h6e;        memory[51777] <=  8'h61;        memory[51778] <=  8'h76;        memory[51779] <=  8'h63;        memory[51780] <=  8'h66;        memory[51781] <=  8'h68;        memory[51782] <=  8'h75;        memory[51783] <=  8'h61;        memory[51784] <=  8'h73;        memory[51785] <=  8'h79;        memory[51786] <=  8'h64;        memory[51787] <=  8'h75;        memory[51788] <=  8'h69;        memory[51789] <=  8'h6a;        memory[51790] <=  8'h61;        memory[51791] <=  8'h6b;        memory[51792] <=  8'h62;        memory[51793] <=  8'h63;        memory[51794] <=  8'h78;        memory[51795] <=  8'h68;        memory[51796] <=  8'h67;        memory[51797] <=  8'h79;        memory[51798] <=  8'h75;        memory[51799] <=  8'h7a;        memory[51800] <=  8'h63;        memory[51801] <=  8'h61;        memory[51802] <=  8'h73;        memory[51803] <=  8'h69;        memory[51804] <=  8'h75;        memory[51805] <=  8'h6f;        memory[51806] <=  8'h69;        memory[51807] <=  8'h6a;        memory[51808] <=  8'h61;        memory[51809] <=  8'h6c;        memory[51810] <=  8'h63;        memory[51811] <=  8'h78;        memory[51812] <=  8'h62;        memory[51813] <=  8'h63;        memory[51814] <=  8'h20;        memory[51815] <=  8'h6e;        memory[51816] <=  8'h76;        memory[51817] <=  8'h63;        memory[51818] <=  8'h61;        memory[51819] <=  8'h64;        memory[51820] <=  8'h73;        memory[51821] <=  8'h67;        memory[51822] <=  8'h79;        memory[51823] <=  8'h68;        memory[51824] <=  8'h75;        memory[51825] <=  8'h61;        memory[51826] <=  8'h6a;        memory[51827] <=  8'h6b;        memory[51828] <=  8'h78;        memory[51829] <=  8'h62;        memory[51830] <=  8'h20;        memory[51831] <=  8'h6e;        memory[51832] <=  8'h76;        memory[51833] <=  8'h63;        memory[51834] <=  8'h61;        memory[51835] <=  8'h73;        memory[51836] <=  8'h67;        memory[51837] <=  8'h68;        memory[51838] <=  8'h75;        memory[51839] <=  8'h6a;        memory[51840] <=  8'h6c;        memory[51841] <=  8'h6b;        memory[51842] <=  8'h63;        memory[51843] <=  8'h78;        memory[51844] <=  8'h20;        memory[51845] <=  8'h6a;        memory[51846] <=  8'h6b;        memory[51847] <=  8'h68;        memory[51848] <=  8'h61;        memory[51849] <=  8'h73;        memory[51850] <=  8'h76;        memory[51851] <=  8'h64;        memory[51852] <=  8'h6e;        memory[51853] <=  8'h20;        memory[51854] <=  8'h62;        memory[51855] <=  8'h6e;        memory[51856] <=  8'h6d;        memory[51857] <=  8'h6b;        memory[51858] <=  8'h77;        memory[51859] <=  8'h64;        memory[51860] <=  8'h6f;        memory[51861] <=  8'h77;        memory[51862] <=  8'h69;        memory[51863] <=  8'h6f;        memory[51864] <=  8'h75;        memory[51865] <=  8'h69;        memory[51866] <=  8'h68;        memory[51867] <=  8'h62;        memory[51868] <=  8'h6e;        memory[51869] <=  8'h6b;        memory[51870] <=  8'h77;        memory[51871] <=  8'h69;        memory[51872] <=  8'h6f;        memory[51873] <=  8'h75;        memory[51874] <=  8'h71;        memory[51875] <=  8'h69;        memory[51876] <=  8'h79;        memory[51877] <=  8'h67;        memory[51878] <=  8'h6a;        memory[51879] <=  8'h64;        memory[51880] <=  8'h61;        memory[51881] <=  8'h76;        memory[51882] <=  8'h62;        memory[51883] <=  8'h6e;        memory[51884] <=  8'h6b;        memory[51885] <=  8'h6f;        memory[51886] <=  8'h70;        memory[51887] <=  8'h64;        memory[51888] <=  8'h76;        memory[51889] <=  8'h69;        memory[51890] <=  8'h6f;        memory[51891] <=  8'h75;        memory[51892] <=  8'h69;        memory[51893] <=  8'h48;        memory[51894] <=  8'h42;        memory[51895] <=  8'h6b;        memory[51896] <=  8'h64;        memory[51897] <=  8'h6e;        memory[51898] <=  8'h6c;        memory[51899] <=  8'h71;        memory[51900] <=  8'h6b;        memory[51901] <=  8'h6d;        memory[51902] <=  8'h6a;        memory[51903] <=  8'h70;        memory[51904] <=  8'h69;        memory[51905] <=  8'h6f;        memory[51906] <=  8'h68;        memory[51907] <=  8'h65;        memory[51908] <=  8'h66;        memory[51909] <=  8'h75;        memory[51910] <=  8'h67;        memory[51911] <=  8'h69;        memory[51912] <=  8'h73;        memory[51913] <=  8'h61;        memory[51914] <=  8'h62;        memory[51915] <=  8'h64;        memory[51916] <=  8'h6b;        memory[51917] <=  8'h6a;        memory[51918] <=  8'h6b;        memory[51919] <=  8'h6c;        memory[51920] <=  8'h6a;        memory[51921] <=  8'h69;        memory[51922] <=  8'h73;        memory[51923] <=  8'h6f;        memory[51924] <=  8'h71;        memory[51925] <=  8'h68;        memory[51926] <=  8'h77;        memory[51927] <=  8'h67;        memory[51928] <=  8'h69;        memory[51929] <=  8'h79;        memory[51930] <=  8'h6a;        memory[51931] <=  8'h64;        memory[51932] <=  8'h76;        memory[51933] <=  8'h62;        memory[51934] <=  8'h6e;        memory[51935] <=  8'h61;        memory[51936] <=  8'h73;        memory[51937] <=  8'h66;        memory[51938] <=  8'h6c;        memory[51939] <=  8'h6b;        memory[51940] <=  8'h64;        memory[51941] <=  8'h6a;        memory[51942] <=  8'h68;        memory[51943] <=  8'h63;        memory[51944] <=  8'h67;        memory[51945] <=  8'h6a;        memory[51946] <=  8'h76;        memory[51947] <=  8'h73;        memory[51948] <=  8'h64;        memory[51949] <=  8'h62;        memory[51950] <=  8'h62;        memory[51951] <=  8'h61;        memory[51952] <=  8'h72;        memory[51953] <=  8'h62;        memory[51954] <=  8'h62;        memory[51955] <=  8'h73;        memory[51956] <=  8'h62;        memory[51957] <=  8'h67;        memory[51958] <=  8'h73;        memory[51959] <=  8'h66;        memory[51960] <=  8'h67;        memory[51961] <=  8'h61;        memory[51962] <=  8'h68;        memory[51963] <=  8'h66;        memory[51964] <=  8'h73;        memory[51965] <=  8'h68;        memory[51966] <=  8'h61;        memory[51967] <=  8'h66;        memory[51968] <=  8'h73;        memory[51969] <=  8'h66;        memory[51970] <=  8'h68;        memory[51971] <=  8'h61;        memory[51972] <=  8'h69;        memory[51973] <=  8'h64;        memory[51974] <=  8'h75;        memory[51975] <=  8'h67;        memory[51976] <=  8'h64;        memory[51977] <=  8'h77;        memory[51978] <=  8'h62;        memory[51979] <=  8'h61;        memory[51980] <=  8'h62;        memory[51981] <=  8'h72;        memory[51982] <=  8'h62;        memory[51983] <=  8'h61;        memory[51984] <=  8'h62;        memory[51985] <=  8'h62;        memory[51986] <=  8'h74;        memory[51987] <=  8'h62;        memory[51988] <=  8'h62;        memory[51989] <=  8'h62;        memory[51990] <=  8'h62;        memory[51991] <=  8'h62;        memory[51992] <=  8'h62;        memory[51993] <=  8'h62;        memory[51994] <=  8'h62;        memory[51995] <=  8'h61;        memory[51996] <=  8'h62;        memory[51997] <=  8'h62;        memory[51998] <=  8'h72;        memory[51999] <=  8'h74;        memory[52000] <=  8'h62;        memory[52001] <=  8'h62;        memory[52002] <=  8'h61;        memory[52003] <=  8'h62;        memory[52004] <=  8'h72;        memory[52005] <=  8'h62;        memory[52006] <=  8'h74;        memory[52007] <=  8'h62;        memory[52008] <=  8'h62;        memory[52009] <=  8'h62;        memory[52010] <=  8'h63;        memory[52011] <=  8'h61;        memory[52012] <=  8'h72;        memory[52013] <=  8'h74;        memory[52014] <=  8'h73;        memory[52015] <=  8'h62;        memory[52016] <=  8'h61;        memory[52017] <=  8'h72;        memory[52018] <=  8'h74;        memory[52019] <=  8'h74;        memory[52020] <=  8'h62;        memory[52021] <=  8'h61;        memory[52022] <=  8'h72;        memory[52023] <=  8'h74;        memory[52024] <=  8'h78;        memory[52025] <=  8'h61;        memory[52026] <=  8'h74;        memory[52027] <=  8'h6b;        memory[52028] <=  8'h73;        memory[52029] <=  8'h68;        memory[52030] <=  8'h63;        memory[52031] <=  8'h66;        memory[52032] <=  8'h69;        memory[52033] <=  8'h77;        memory[52034] <=  8'h68;        memory[52035] <=  8'h61;        memory[52036] <=  8'h74;        memory[52037] <=  8'h61;        memory[52038] <=  8'h6e;        memory[52039] <=  8'h61;        memory[52040] <=  8'h62;        memory[52041] <=  8'h61;        memory[52042] <=  8'h63;        memory[52043] <=  8'h61;        memory[52044] <=  8'h74;        memory[52045] <=  8'h61;        memory[52046] <=  8'h62;        memory[52047] <=  8'h61;        memory[52048] <=  8'h72;        memory[52049] <=  8'h63;        memory[52050] <=  8'h61;        memory[52051] <=  8'h68;        memory[52052] <=  8'h64;        memory[52053] <=  8'h75;        memory[52054] <=  8'h63;        memory[52055] <=  8'h74;        memory[52056] <=  8'h61;        memory[52057] <=  8'h64;        memory[52058] <=  8'h61;        memory[52059] <=  8'h61;        memory[52060] <=  8'h63;        memory[52061] <=  8'h61;        memory[52062] <=  8'h72;        memory[52063] <=  8'h63;        memory[52064] <=  8'h74;        memory[52065] <=  8'h72;        memory[52066] <=  8'h63;        memory[52067] <=  8'h61;        memory[52068] <=  8'h74;        memory[52069] <=  8'h72;        memory[52070] <=  8'h63;        memory[52071] <=  8'h61;        memory[52072] <=  8'h74;        memory[52073] <=  8'h63;        memory[52074] <=  8'h62;        memory[52075] <=  8'h61;        memory[52076] <=  8'h74;        memory[52077] <=  8'h62;        memory[52078] <=  8'h72;        memory[52079] <=  8'h63;        memory[52080] <=  8'h61;        memory[52081] <=  8'h74;        memory[52082] <=  8'h72;        memory[52083] <=  8'h6e;        memory[52084] <=  8'h62;        memory[52085] <=  8'h61;        memory[52086] <=  8'h63;        memory[52087] <=  8'h61;        memory[52088] <=  8'h74;        memory[52089] <=  8'h79;        memory[52090] <=  8'h73;        memory[52091] <=  8'h6e;        memory[52092] <=  8'h63;        memory[52093] <=  8'h74;        memory[52094] <=  8'h61;        memory[52095] <=  8'h6e;        memory[52096] <=  8'h62;        memory[52097] <=  8'h61;        memory[52098] <=  8'h63;        memory[52099] <=  8'h72;        memory[52100] <=  8'h6e;        memory[52101] <=  8'h74;        memory[52102] <=  8'h61;        memory[52103] <=  8'h62;        memory[52104] <=  8'h74;        memory[52105] <=  8'h6e;        memory[52106] <=  8'h61;        memory[52107] <=  8'h72;        memory[52108] <=  8'h62;        memory[52109] <=  8'h78;        memory[52110] <=  8'h74;        memory[52111] <=  8'h61;        memory[52112] <=  8'h72;        memory[52113] <=  8'h62;        memory[52114] <=  8'h61;        memory[52115] <=  8'h72;        memory[52116] <=  8'h74;        memory[52117] <=  8'h74;        memory[52118] <=  8'h62;        memory[52119] <=  8'h61;        memory[52120] <=  8'h72;        memory[52121] <=  8'h74;        memory[52122] <=  8'h78;        memory[52123] <=  8'h61;        memory[52124] <=  8'h74;        memory[52125] <=  8'h6b;        memory[52126] <=  8'h73;        memory[52127] <=  8'h68;        memory[52128] <=  8'h63;        memory[52129] <=  8'h66;        memory[52130] <=  8'h69;        memory[52131] <=  8'h77;        memory[52132] <=  8'h68;        memory[52133] <=  8'h61;        memory[52134] <=  8'h74;        memory[52135] <=  8'h61;        memory[52136] <=  8'h6e;        memory[52137] <=  8'h61;        memory[52138] <=  8'h62;        memory[52139] <=  8'h61;        memory[52140] <=  8'h63;        memory[52141] <=  8'h61;        memory[52142] <=  8'h74;        memory[52143] <=  8'h61;        memory[52144] <=  8'h62;        memory[52145] <=  8'h61;        memory[52146] <=  8'h72;        memory[52147] <=  8'h63;        memory[52148] <=  8'h61;        memory[52149] <=  8'h68;        memory[52150] <=  8'h64;        memory[52151] <=  8'h75;        memory[52152] <=  8'h63;        memory[52153] <=  8'h74;        memory[52154] <=  8'h61;        memory[52155] <=  8'h64;        memory[52156] <=  8'h61;        memory[52157] <=  8'h61;        memory[52158] <=  8'h63;        memory[52159] <=  8'h61;        memory[52160] <=  8'h72;        memory[52161] <=  8'h63;        memory[52162] <=  8'h74;        memory[52163] <=  8'h72;        memory[52164] <=  8'h63;        memory[52165] <=  8'h61;        memory[52166] <=  8'h74;        memory[52167] <=  8'h72;        memory[52168] <=  8'h63;        memory[52169] <=  8'h61;        memory[52170] <=  8'h74;        memory[52171] <=  8'h63;        memory[52172] <=  8'h62;        memory[52173] <=  8'h61;        memory[52174] <=  8'h74;        memory[52175] <=  8'h62;        memory[52176] <=  8'h72;        memory[52177] <=  8'h63;        memory[52178] <=  8'h61;        memory[52179] <=  8'h74;        memory[52180] <=  8'h72;        memory[52181] <=  8'h6e;        memory[52182] <=  8'h62;        memory[52183] <=  8'h61;        memory[52184] <=  8'h63;        memory[52185] <=  8'h61;        memory[52186] <=  8'h74;        memory[52187] <=  8'h79;        memory[52188] <=  8'h73;        memory[52189] <=  8'h6e;        memory[52190] <=  8'h63;        memory[52191] <=  8'h74;        memory[52192] <=  8'h61;        memory[52193] <=  8'h6e;        memory[52194] <=  8'h62;        memory[52195] <=  8'h61;        memory[52196] <=  8'h63;        memory[52197] <=  8'h72;        memory[52198] <=  8'h6e;        memory[52199] <=  8'h74;        memory[52200] <=  8'h61;        memory[52201] <=  8'h62;        memory[52202] <=  8'h74;        memory[52203] <=  8'h6e;        memory[52204] <=  8'h61;        memory[52205] <=  8'h72;        memory[52206] <=  8'h62;        memory[52207] <=  8'h78;        memory[52208] <=  8'h74;        memory[52209] <=  8'h61;        memory[52210] <=  8'h72;        memory[52211] <=  8'h62;        memory[52212] <=  8'h61;        memory[52213] <=  8'h72;        memory[52214] <=  8'h74;        memory[52215] <=  8'h74;        memory[52216] <=  8'h62;        memory[52217] <=  8'h61;        memory[52218] <=  8'h72;        memory[52219] <=  8'h74;        memory[52220] <=  8'h78;        memory[52221] <=  8'h61;        memory[52222] <=  8'h74;        memory[52223] <=  8'h6b;        memory[52224] <=  8'h73;        memory[52225] <=  8'h68;        memory[52226] <=  8'h63;        memory[52227] <=  8'h66;        memory[52228] <=  8'h69;        memory[52229] <=  8'h77;        memory[52230] <=  8'h68;        memory[52231] <=  8'h61;        memory[52232] <=  8'h74;        memory[52233] <=  8'h61;        memory[52234] <=  8'h6e;        memory[52235] <=  8'h61;        memory[52236] <=  8'h62;        memory[52237] <=  8'h61;        memory[52238] <=  8'h63;        memory[52239] <=  8'h61;        memory[52240] <=  8'h74;        memory[52241] <=  8'h61;        memory[52242] <=  8'h62;        memory[52243] <=  8'h61;        memory[52244] <=  8'h72;        memory[52245] <=  8'h63;        memory[52246] <=  8'h61;        memory[52247] <=  8'h68;        memory[52248] <=  8'h64;        memory[52249] <=  8'h75;        memory[52250] <=  8'h63;        memory[52251] <=  8'h74;        memory[52252] <=  8'h61;        memory[52253] <=  8'h64;        memory[52254] <=  8'h61;        memory[52255] <=  8'h61;        memory[52256] <=  8'h63;        memory[52257] <=  8'h61;        memory[52258] <=  8'h72;        memory[52259] <=  8'h63;        memory[52260] <=  8'h74;        memory[52261] <=  8'h72;        memory[52262] <=  8'h63;        memory[52263] <=  8'h61;        memory[52264] <=  8'h74;        memory[52265] <=  8'h72;        memory[52266] <=  8'h63;        memory[52267] <=  8'h61;        memory[52268] <=  8'h74;        memory[52269] <=  8'h63;        memory[52270] <=  8'h62;        memory[52271] <=  8'h61;        memory[52272] <=  8'h74;        memory[52273] <=  8'h62;        memory[52274] <=  8'h72;        memory[52275] <=  8'h63;        memory[52276] <=  8'h61;        memory[52277] <=  8'h74;        memory[52278] <=  8'h72;        memory[52279] <=  8'h6e;        memory[52280] <=  8'h62;        memory[52281] <=  8'h61;        memory[52282] <=  8'h63;        memory[52283] <=  8'h61;        memory[52284] <=  8'h74;        memory[52285] <=  8'h79;        memory[52286] <=  8'h73;        memory[52287] <=  8'h6e;        memory[52288] <=  8'h63;        memory[52289] <=  8'h74;        memory[52290] <=  8'h61;        memory[52291] <=  8'h6e;        memory[52292] <=  8'h62;        memory[52293] <=  8'h61;        memory[52294] <=  8'h63;        memory[52295] <=  8'h72;        memory[52296] <=  8'h6e;        memory[52297] <=  8'h74;        memory[52298] <=  8'h61;        memory[52299] <=  8'h62;        memory[52300] <=  8'h74;        memory[52301] <=  8'h6e;        memory[52302] <=  8'h61;        memory[52303] <=  8'h72;        memory[52304] <=  8'h62;        memory[52305] <=  8'h78;        memory[52306] <=  8'h74;        memory[52307] <=  8'h61;        memory[52308] <=  8'h72;        memory[52309] <=  8'h5d;        memory[52310] <=  8'h5d;        memory[52311] <=  8'h65;        memory[52312] <=  8'h66;        memory[52313] <=  8'h77;        memory[52314] <=  8'h65;        memory[52315] <=  8'h5d;        memory[52316] <=  8'h65;        memory[52317] <=  8'h67;        memory[52318] <=  8'h73;        memory[52319] <=  8'h67;        memory[52320] <=  8'h66;        memory[52321] <=  8'h62;        memory[52322] <=  8'h61;        memory[52323] <=  8'h72;        memory[52324] <=  8'h74;        memory[52325] <=  8'h74;        memory[52326] <=  8'h62;        memory[52327] <=  8'h61;        memory[52328] <=  8'h72;        memory[52329] <=  8'h74;        memory[52330] <=  8'h78;        memory[52331] <=  8'h61;        memory[52332] <=  8'h74;        memory[52333] <=  8'h6b;        memory[52334] <=  8'h73;        memory[52335] <=  8'h68;        memory[52336] <=  8'h63;        memory[52337] <=  8'h66;        memory[52338] <=  8'h69;        memory[52339] <=  8'h77;        memory[52340] <=  8'h68;        memory[52341] <=  8'h61;        memory[52342] <=  8'h74;        memory[52343] <=  8'h61;        memory[52344] <=  8'h6e;        memory[52345] <=  8'h61;        memory[52346] <=  8'h62;        memory[52347] <=  8'h61;        memory[52348] <=  8'h63;        memory[52349] <=  8'h61;        memory[52350] <=  8'h74;        memory[52351] <=  8'h61;        memory[52352] <=  8'h62;        memory[52353] <=  8'h61;        memory[52354] <=  8'h72;        memory[52355] <=  8'h63;        memory[52356] <=  8'h61;        memory[52357] <=  8'h68;        memory[52358] <=  8'h64;        memory[52359] <=  8'h75;        memory[52360] <=  8'h63;        memory[52361] <=  8'h74;        memory[52362] <=  8'h61;        memory[52363] <=  8'h64;        memory[52364] <=  8'h61;        memory[52365] <=  8'h61;        memory[52366] <=  8'h63;        memory[52367] <=  8'h61;        memory[52368] <=  8'h72;        memory[52369] <=  8'h63;        memory[52370] <=  8'h74;        memory[52371] <=  8'h72;        memory[52372] <=  8'h63;        memory[52373] <=  8'h61;        memory[52374] <=  8'h74;        memory[52375] <=  8'h72;        memory[52376] <=  8'h63;        memory[52377] <=  8'h61;        memory[52378] <=  8'h74;        memory[52379] <=  8'h63;        memory[52380] <=  8'h62;        memory[52381] <=  8'h61;        memory[52382] <=  8'h74;        memory[52383] <=  8'h62;        memory[52384] <=  8'h72;        memory[52385] <=  8'h63;        memory[52386] <=  8'h61;        memory[52387] <=  8'h74;        memory[52388] <=  8'h72;        memory[52389] <=  8'h6e;        memory[52390] <=  8'h62;        memory[52391] <=  8'h61;        memory[52392] <=  8'h63;        memory[52393] <=  8'h61;        memory[52394] <=  8'h74;        memory[52395] <=  8'h79;        memory[52396] <=  8'h73;        memory[52397] <=  8'h6e;        memory[52398] <=  8'h63;        memory[52399] <=  8'h74;        memory[52400] <=  8'h61;        memory[52401] <=  8'h6e;        memory[52402] <=  8'h62;        memory[52403] <=  8'h61;        memory[52404] <=  8'h63;        memory[52405] <=  8'h72;        memory[52406] <=  8'h6e;        memory[52407] <=  8'h74;        memory[52408] <=  8'h61;        memory[52409] <=  8'h62;        memory[52410] <=  8'h74;        memory[52411] <=  8'h6e;        memory[52412] <=  8'h61;        memory[52413] <=  8'h72;        memory[52414] <=  8'h62;        memory[52415] <=  8'h78;        memory[52416] <=  8'h74;        memory[52417] <=  8'h61;        memory[52418] <=  8'h72;        memory[52419] <=  8'h62;        memory[52420] <=  8'h61;        memory[52421] <=  8'h72;        memory[52422] <=  8'h74;        memory[52423] <=  8'h74;        memory[52424] <=  8'h62;        memory[52425] <=  8'h61;        memory[52426] <=  8'h72;        memory[52427] <=  8'h74;        memory[52428] <=  8'h78;        memory[52429] <=  8'h61;        memory[52430] <=  8'h74;        memory[52431] <=  8'h6b;        memory[52432] <=  8'h73;        memory[52433] <=  8'h68;        memory[52434] <=  8'h63;        memory[52435] <=  8'h66;        memory[52436] <=  8'h69;        memory[52437] <=  8'h77;        memory[52438] <=  8'h68;        memory[52439] <=  8'h61;        memory[52440] <=  8'h74;        memory[52441] <=  8'h61;        memory[52442] <=  8'h6e;        memory[52443] <=  8'h61;        memory[52444] <=  8'h62;        memory[52445] <=  8'h61;        memory[52446] <=  8'h63;        memory[52447] <=  8'h61;        memory[52448] <=  8'h74;        memory[52449] <=  8'h61;        memory[52450] <=  8'h62;        memory[52451] <=  8'h61;        memory[52452] <=  8'h72;        memory[52453] <=  8'h63;        memory[52454] <=  8'h61;        memory[52455] <=  8'h68;        memory[52456] <=  8'h64;        memory[52457] <=  8'h75;        memory[52458] <=  8'h63;        memory[52459] <=  8'h74;        memory[52460] <=  8'h61;        memory[52461] <=  8'h64;        memory[52462] <=  8'h61;        memory[52463] <=  8'h61;        memory[52464] <=  8'h63;        memory[52465] <=  8'h61;        memory[52466] <=  8'h72;        memory[52467] <=  8'h63;        memory[52468] <=  8'h74;        memory[52469] <=  8'h72;        memory[52470] <=  8'h63;        memory[52471] <=  8'h61;        memory[52472] <=  8'h74;        memory[52473] <=  8'h72;        memory[52474] <=  8'h63;        memory[52475] <=  8'h61;        memory[52476] <=  8'h74;        memory[52477] <=  8'h63;        memory[52478] <=  8'h62;        memory[52479] <=  8'h61;        memory[52480] <=  8'h74;        memory[52481] <=  8'h62;        memory[52482] <=  8'h72;        memory[52483] <=  8'h63;        memory[52484] <=  8'h61;        memory[52485] <=  8'h74;        memory[52486] <=  8'h72;        memory[52487] <=  8'h6e;        memory[52488] <=  8'h62;        memory[52489] <=  8'h61;        memory[52490] <=  8'h63;        memory[52491] <=  8'h61;        memory[52492] <=  8'h74;        memory[52493] <=  8'h79;        memory[52494] <=  8'h73;        memory[52495] <=  8'h6e;        memory[52496] <=  8'h63;        memory[52497] <=  8'h74;        memory[52498] <=  8'h61;        memory[52499] <=  8'h6e;        memory[52500] <=  8'h62;        memory[52501] <=  8'h61;        memory[52502] <=  8'h63;        memory[52503] <=  8'h72;        memory[52504] <=  8'h6e;        memory[52505] <=  8'h74;        memory[52506] <=  8'h61;        memory[52507] <=  8'h62;        memory[52508] <=  8'h74;        memory[52509] <=  8'h6e;        memory[52510] <=  8'h61;        memory[52511] <=  8'h72;        memory[52512] <=  8'h62;        memory[52513] <=  8'h78;        memory[52514] <=  8'h74;        memory[52515] <=  8'h61;        memory[52516] <=  8'h72;        memory[52517] <=  8'h64;        memory[52518] <=  8'h66;        memory[52519] <=  8'h73;        memory[52520] <=  8'h67;        memory[52521] <=  8'h76;        memory[52522] <=  8'h68;        memory[52523] <=  8'h62;        memory[52524] <=  8'h6b;        memory[52525] <=  8'h6a;        memory[52526] <=  8'h6e;        memory[52527] <=  8'h6d;        memory[52528] <=  8'h62;        memory[52529] <=  8'h76;        memory[52530] <=  8'h78;        memory[52531] <=  8'h63;        memory[52532] <=  8'h73;        memory[52533] <=  8'h66;        memory[52534] <=  8'h72;        memory[52535] <=  8'h74;        memory[52536] <=  8'h79;        memory[52537] <=  8'h75;        memory[52538] <=  8'h6a;        memory[52539] <=  8'h6e;        memory[52540] <=  8'h62;        memory[52541] <=  8'h76;        memory[52542] <=  8'h63;        memory[52543] <=  8'h64;        memory[52544] <=  8'h74;        memory[52545] <=  8'h79;        memory[52546] <=  8'h75;        memory[52547] <=  8'h69;        memory[52548] <=  8'h6b;        memory[52549] <=  8'h6d;        memory[52550] <=  8'h6e;        memory[52551] <=  8'h62;        memory[52552] <=  8'h76;        memory[52553] <=  8'h63;        memory[52554] <=  8'h78;        memory[52555] <=  8'h73;        memory[52556] <=  8'h64;        memory[52557] <=  8'h72;        memory[52558] <=  8'h74;        memory[52559] <=  8'h79;        memory[52560] <=  8'h75;        memory[52561] <=  8'h69;        memory[52562] <=  8'h6b;        memory[52563] <=  8'h6d;        memory[52564] <=  8'h6e;        memory[52565] <=  8'h62;        memory[52566] <=  8'h76;        memory[52567] <=  8'h63;        memory[52568] <=  8'h73;        memory[52569] <=  8'h77;        memory[52570] <=  8'h33;        memory[52571] <=  8'h34;        memory[52572] <=  8'h35;        memory[52573] <=  8'h36;        memory[52574] <=  8'h37;        memory[52575] <=  8'h38;        memory[52576] <=  8'h69;        memory[52577] <=  8'h6b;        memory[52578] <=  8'h6d;        memory[52579] <=  8'h6e;        memory[52580] <=  8'h62;        memory[52581] <=  8'h76;        memory[52582] <=  8'h63;        memory[52583] <=  8'h64;        memory[52584] <=  8'h65;        memory[52585] <=  8'h72;        memory[52586] <=  8'h36;        memory[52587] <=  8'h37;        memory[52588] <=  8'h38;        memory[52589] <=  8'h69;        memory[52590] <=  8'h6f;        memory[52591] <=  8'h6b;        memory[52592] <=  8'h6a;        memory[52593] <=  8'h6e;        memory[52594] <=  8'h62;        memory[52595] <=  8'h76;        memory[52596] <=  8'h63;        memory[52597] <=  8'h64;        memory[52598] <=  8'h72;        memory[52599] <=  8'h74;        memory[52600] <=  8'h79;        memory[52601] <=  8'h75;        memory[52602] <=  8'h73;        memory[52603] <=  8'h6a;        memory[52604] <=  8'h63;        memory[52605] <=  8'h6e;        memory[52606] <=  8'h62;        memory[52607] <=  8'h64;        memory[52608] <=  8'h66;        memory[52609] <=  8'h73;        memory[52610] <=  8'h74;        memory[52611] <=  8'h79;        memory[52612] <=  8'h75;        memory[52613] <=  8'h61;        memory[52614] <=  8'h69;        memory[52615] <=  8'h6b;        memory[52616] <=  8'h78;        memory[52617] <=  8'h6d;        memory[52618] <=  8'h6e;        memory[52619] <=  8'h73;        memory[52620] <=  8'h6a;        memory[52621] <=  8'h6f;        memory[52622] <=  8'h64;        memory[52623] <=  8'h6c;        memory[52624] <=  8'h63;        memory[52625] <=  8'h78;        memory[52626] <=  8'h62;        memory[52627] <=  8'h61;        memory[52628] <=  8'h72;        memory[52629] <=  8'h74;        memory[52630] <=  8'h78;        memory[52631] <=  8'h61;        memory[52632] <=  8'h74;        memory[52633] <=  8'h6b;        memory[52634] <=  8'h73;        memory[52635] <=  8'h68;        memory[52636] <=  8'h63;        memory[52637] <=  8'h66;        memory[52638] <=  8'h69;        memory[52639] <=  8'h77;        memory[52640] <=  8'h68;        memory[52641] <=  8'h61;        memory[52642] <=  8'h74;        memory[52643] <=  8'h61;        memory[52644] <=  8'h6e;        memory[52645] <=  8'h61;        memory[52646] <=  8'h62;        memory[52647] <=  8'h61;        memory[52648] <=  8'h63;        memory[52649] <=  8'h61;        memory[52650] <=  8'h74;        memory[52651] <=  8'h61;        memory[52652] <=  8'h62;        memory[52653] <=  8'h61;        memory[52654] <=  8'h72;        memory[52655] <=  8'h63;        memory[52656] <=  8'h61;        memory[52657] <=  8'h68;        memory[52658] <=  8'h64;        memory[52659] <=  8'h75;        memory[52660] <=  8'h63;        memory[52661] <=  8'h74;        memory[52662] <=  8'h61;        memory[52663] <=  8'h64;        memory[52664] <=  8'h61;        memory[52665] <=  8'h61;        memory[52666] <=  8'h63;        memory[52667] <=  8'h61;        memory[52668] <=  8'h72;        memory[52669] <=  8'h62;        memory[52670] <=  8'h61;        memory[52671] <=  8'h72;        memory[52672] <=  8'h74;        memory[52673] <=  8'h78;        memory[52674] <=  8'h61;        memory[52675] <=  8'h74;        memory[52676] <=  8'h6b;        memory[52677] <=  8'h73;        memory[52678] <=  8'h68;        memory[52679] <=  8'h63;        memory[52680] <=  8'h66;        memory[52681] <=  8'h69;        memory[52682] <=  8'h77;        memory[52683] <=  8'h68;        memory[52684] <=  8'h61;        memory[52685] <=  8'h74;        memory[52686] <=  8'h61;        memory[52687] <=  8'h6e;        memory[52688] <=  8'h61;        memory[52689] <=  8'h62;        memory[52690] <=  8'h61;        memory[52691] <=  8'h63;        memory[52692] <=  8'h61;        memory[52693] <=  8'h74;        memory[52694] <=  8'h61;        memory[52695] <=  8'h62;        memory[52696] <=  8'h61;        memory[52697] <=  8'h72;        memory[52698] <=  8'h63;        memory[52699] <=  8'h61;        memory[52700] <=  8'h68;        memory[52701] <=  8'h64;        memory[52702] <=  8'h75;        memory[52703] <=  8'h63;        memory[52704] <=  8'h74;        memory[52705] <=  8'h61;        memory[52706] <=  8'h64;        memory[52707] <=  8'h61;        memory[52708] <=  8'h61;        memory[52709] <=  8'h63;        memory[52710] <=  8'h61;        memory[52711] <=  8'h72;        memory[52712] <=  8'h62;        memory[52713] <=  8'h61;        memory[52714] <=  8'h72;        memory[52715] <=  8'h74;        memory[52716] <=  8'h78;        memory[52717] <=  8'h61;        memory[52718] <=  8'h74;        memory[52719] <=  8'h6b;        memory[52720] <=  8'h73;        memory[52721] <=  8'h68;        memory[52722] <=  8'h63;        memory[52723] <=  8'h66;        memory[52724] <=  8'h69;        memory[52725] <=  8'h77;        memory[52726] <=  8'h68;        memory[52727] <=  8'h61;        memory[52728] <=  8'h74;        memory[52729] <=  8'h61;        memory[52730] <=  8'h6e;        memory[52731] <=  8'h61;        memory[52732] <=  8'h62;        memory[52733] <=  8'h61;        memory[52734] <=  8'h63;        memory[52735] <=  8'h61;        memory[52736] <=  8'h74;        memory[52737] <=  8'h61;        memory[52738] <=  8'h62;        memory[52739] <=  8'h61;        memory[52740] <=  8'h72;        memory[52741] <=  8'h63;        memory[52742] <=  8'h61;        memory[52743] <=  8'h68;        memory[52744] <=  8'h64;        memory[52745] <=  8'h75;        memory[52746] <=  8'h63;        memory[52747] <=  8'h74;        memory[52748] <=  8'h61;        memory[52749] <=  8'h64;        memory[52750] <=  8'h61;        memory[52751] <=  8'h61;        memory[52752] <=  8'h63;        memory[52753] <=  8'h61;        memory[52754] <=  8'h72;        memory[52755] <=  8'h62;        memory[52756] <=  8'h61;        memory[52757] <=  8'h72;        memory[52758] <=  8'h74;        memory[52759] <=  8'h78;        memory[52760] <=  8'h61;        memory[52761] <=  8'h74;        memory[52762] <=  8'h6b;        memory[52763] <=  8'h73;        memory[52764] <=  8'h68;        memory[52765] <=  8'h63;        memory[52766] <=  8'h66;        memory[52767] <=  8'h69;        memory[52768] <=  8'h77;        memory[52769] <=  8'h68;        memory[52770] <=  8'h61;        memory[52771] <=  8'h74;        memory[52772] <=  8'h61;        memory[52773] <=  8'h6e;        memory[52774] <=  8'h61;        memory[52775] <=  8'h62;        memory[52776] <=  8'h61;        memory[52777] <=  8'h63;        memory[52778] <=  8'h61;        memory[52779] <=  8'h74;        memory[52780] <=  8'h61;        memory[52781] <=  8'h62;        memory[52782] <=  8'h61;        memory[52783] <=  8'h72;        memory[52784] <=  8'h63;        memory[52785] <=  8'h61;        memory[52786] <=  8'h68;        memory[52787] <=  8'h64;        memory[52788] <=  8'h75;        memory[52789] <=  8'h63;        memory[52790] <=  8'h74;        memory[52791] <=  8'h61;        memory[52792] <=  8'h64;        memory[52793] <=  8'h61;        memory[52794] <=  8'h61;        memory[52795] <=  8'h63;        memory[52796] <=  8'h61;        memory[52797] <=  8'h72;        memory[52798] <=  8'h62;        memory[52799] <=  8'h61;        memory[52800] <=  8'h72;        memory[52801] <=  8'h74;        memory[52802] <=  8'h78;        memory[52803] <=  8'h61;        memory[52804] <=  8'h74;        memory[52805] <=  8'h6b;        memory[52806] <=  8'h73;        memory[52807] <=  8'h68;        memory[52808] <=  8'h63;        memory[52809] <=  8'h66;        memory[52810] <=  8'h69;        memory[52811] <=  8'h77;        memory[52812] <=  8'h68;        memory[52813] <=  8'h61;        memory[52814] <=  8'h74;        memory[52815] <=  8'h61;        memory[52816] <=  8'h6e;        memory[52817] <=  8'h61;        memory[52818] <=  8'h62;        memory[52819] <=  8'h61;        memory[52820] <=  8'h63;        memory[52821] <=  8'h61;        memory[52822] <=  8'h74;        memory[52823] <=  8'h61;        memory[52824] <=  8'h62;        memory[52825] <=  8'h61;        memory[52826] <=  8'h72;        memory[52827] <=  8'h63;        memory[52828] <=  8'h61;        memory[52829] <=  8'h68;        memory[52830] <=  8'h64;        memory[52831] <=  8'h75;        memory[52832] <=  8'h63;        memory[52833] <=  8'h74;        memory[52834] <=  8'h61;        memory[52835] <=  8'h64;        memory[52836] <=  8'h61;        memory[52837] <=  8'h61;        memory[52838] <=  8'h63;        memory[52839] <=  8'h61;        memory[52840] <=  8'h72;        memory[52841] <=  8'h62;        memory[52842] <=  8'h61;        memory[52843] <=  8'h72;        memory[52844] <=  8'h74;        memory[52845] <=  8'h78;        memory[52846] <=  8'h61;        memory[52847] <=  8'h74;        memory[52848] <=  8'h6b;        memory[52849] <=  8'h73;        memory[52850] <=  8'h68;        memory[52851] <=  8'h63;        memory[52852] <=  8'h66;        memory[52853] <=  8'h69;        memory[52854] <=  8'h77;        memory[52855] <=  8'h68;        memory[52856] <=  8'h61;        memory[52857] <=  8'h74;        memory[52858] <=  8'h61;        memory[52859] <=  8'h6e;        memory[52860] <=  8'h61;        memory[52861] <=  8'h62;        memory[52862] <=  8'h61;        memory[52863] <=  8'h63;        memory[52864] <=  8'h61;        memory[52865] <=  8'h74;        memory[52866] <=  8'h61;        memory[52867] <=  8'h62;        memory[52868] <=  8'h61;        memory[52869] <=  8'h72;        memory[52870] <=  8'h63;        memory[52871] <=  8'h61;        memory[52872] <=  8'h68;        memory[52873] <=  8'h64;        memory[52874] <=  8'h75;        memory[52875] <=  8'h63;        memory[52876] <=  8'h74;        memory[52877] <=  8'h61;        memory[52878] <=  8'h64;        memory[52879] <=  8'h61;        memory[52880] <=  8'h61;        memory[52881] <=  8'h63;        memory[52882] <=  8'h61;        memory[52883] <=  8'h72;        memory[52884] <=  8'h62;        memory[52885] <=  8'h61;        memory[52886] <=  8'h72;        memory[52887] <=  8'h74;        memory[52888] <=  8'h78;        memory[52889] <=  8'h61;        memory[52890] <=  8'h74;        memory[52891] <=  8'h6b;        memory[52892] <=  8'h73;        memory[52893] <=  8'h68;        memory[52894] <=  8'h63;        memory[52895] <=  8'h66;        memory[52896] <=  8'h69;        memory[52897] <=  8'h77;        memory[52898] <=  8'h68;        memory[52899] <=  8'h61;        memory[52900] <=  8'h74;        memory[52901] <=  8'h61;        memory[52902] <=  8'h6e;        memory[52903] <=  8'h61;        memory[52904] <=  8'h62;        memory[52905] <=  8'h61;        memory[52906] <=  8'h63;        memory[52907] <=  8'h61;        memory[52908] <=  8'h74;        memory[52909] <=  8'h61;        memory[52910] <=  8'h62;        memory[52911] <=  8'h61;        memory[52912] <=  8'h72;        memory[52913] <=  8'h63;        memory[52914] <=  8'h61;        memory[52915] <=  8'h68;        memory[52916] <=  8'h64;        memory[52917] <=  8'h75;        memory[52918] <=  8'h63;        memory[52919] <=  8'h74;        memory[52920] <=  8'h61;        memory[52921] <=  8'h64;        memory[52922] <=  8'h61;        memory[52923] <=  8'h61;        memory[52924] <=  8'h63;        memory[52925] <=  8'h61;        memory[52926] <=  8'h72;        memory[52927] <=  8'h62;        memory[52928] <=  8'h61;        memory[52929] <=  8'h72;        memory[52930] <=  8'h74;        memory[52931] <=  8'h78;        memory[52932] <=  8'h61;        memory[52933] <=  8'h74;        memory[52934] <=  8'h6b;        memory[52935] <=  8'h73;        memory[52936] <=  8'h68;        memory[52937] <=  8'h63;        memory[52938] <=  8'h66;        memory[52939] <=  8'h69;        memory[52940] <=  8'h77;        memory[52941] <=  8'h68;        memory[52942] <=  8'h61;        memory[52943] <=  8'h74;        memory[52944] <=  8'h61;        memory[52945] <=  8'h6e;        memory[52946] <=  8'h61;        memory[52947] <=  8'h62;        memory[52948] <=  8'h61;        memory[52949] <=  8'h63;        memory[52950] <=  8'h61;        memory[52951] <=  8'h74;        memory[52952] <=  8'h61;        memory[52953] <=  8'h62;        memory[52954] <=  8'h61;        memory[52955] <=  8'h72;        memory[52956] <=  8'h63;        memory[52957] <=  8'h61;        memory[52958] <=  8'h68;        memory[52959] <=  8'h64;        memory[52960] <=  8'h75;        memory[52961] <=  8'h63;        memory[52962] <=  8'h74;        memory[52963] <=  8'h61;        memory[52964] <=  8'h64;        memory[52965] <=  8'h61;        memory[52966] <=  8'h61;        memory[52967] <=  8'h63;        memory[52968] <=  8'h61;        memory[52969] <=  8'h72;        memory[52970] <=  8'h62;        memory[52971] <=  8'h61;        memory[52972] <=  8'h72;        memory[52973] <=  8'h74;        memory[52974] <=  8'h78;        memory[52975] <=  8'h61;        memory[52976] <=  8'h74;        memory[52977] <=  8'h6b;        memory[52978] <=  8'h73;        memory[52979] <=  8'h68;        memory[52980] <=  8'h63;        memory[52981] <=  8'h66;        memory[52982] <=  8'h69;        memory[52983] <=  8'h77;        memory[52984] <=  8'h68;        memory[52985] <=  8'h61;        memory[52986] <=  8'h74;        memory[52987] <=  8'h61;        memory[52988] <=  8'h6e;        memory[52989] <=  8'h61;        memory[52990] <=  8'h62;        memory[52991] <=  8'h61;        memory[52992] <=  8'h63;        memory[52993] <=  8'h61;        memory[52994] <=  8'h74;        memory[52995] <=  8'h61;        memory[52996] <=  8'h62;        memory[52997] <=  8'h61;        memory[52998] <=  8'h72;        memory[52999] <=  8'h63;        memory[53000] <=  8'h61;        memory[53001] <=  8'h68;        memory[53002] <=  8'h64;        memory[53003] <=  8'h75;        memory[53004] <=  8'h63;        memory[53005] <=  8'h74;        memory[53006] <=  8'h61;        memory[53007] <=  8'h64;        memory[53008] <=  8'h61;        memory[53009] <=  8'h61;        memory[53010] <=  8'h63;        memory[53011] <=  8'h61;        memory[53012] <=  8'h72;        memory[53013] <=  8'h62;        memory[53014] <=  8'h61;        memory[53015] <=  8'h72;        memory[53016] <=  8'h74;        memory[53017] <=  8'h74;        memory[53018] <=  8'h62;        memory[53019] <=  8'h61;        memory[53020] <=  8'h72;        memory[53021] <=  8'h74;        memory[53022] <=  8'h78;        memory[53023] <=  8'h61;        memory[53024] <=  8'h74;        memory[53025] <=  8'h6b;        memory[53026] <=  8'h73;        memory[53027] <=  8'h68;        memory[53028] <=  8'h63;        memory[53029] <=  8'h66;        memory[53030] <=  8'h69;        memory[53031] <=  8'h77;        memory[53032] <=  8'h68;        memory[53033] <=  8'h61;        memory[53034] <=  8'h74;        memory[53035] <=  8'h61;        memory[53036] <=  8'h6e;        memory[53037] <=  8'h61;        memory[53038] <=  8'h62;        memory[53039] <=  8'h61;        memory[53040] <=  8'h63;        memory[53041] <=  8'h61;        memory[53042] <=  8'h74;        memory[53043] <=  8'h61;        memory[53044] <=  8'h62;        memory[53045] <=  8'h61;        memory[53046] <=  8'h72;        memory[53047] <=  8'h63;        memory[53048] <=  8'h61;        memory[53049] <=  8'h68;        memory[53050] <=  8'h64;        memory[53051] <=  8'h75;        memory[53052] <=  8'h63;        memory[53053] <=  8'h74;        memory[53054] <=  8'h61;        memory[53055] <=  8'h64;        memory[53056] <=  8'h61;        memory[53057] <=  8'h61;        memory[53058] <=  8'h63;        memory[53059] <=  8'h61;        memory[53060] <=  8'h72;        memory[53061] <=  8'h63;        memory[53062] <=  8'h74;        memory[53063] <=  8'h72;        memory[53064] <=  8'h63;        memory[53065] <=  8'h61;        memory[53066] <=  8'h74;        memory[53067] <=  8'h72;        memory[53068] <=  8'h63;        memory[53069] <=  8'h61;        memory[53070] <=  8'h74;        memory[53071] <=  8'h63;        memory[53072] <=  8'h62;        memory[53073] <=  8'h61;        memory[53074] <=  8'h74;        memory[53075] <=  8'h62;        memory[53076] <=  8'h72;        memory[53077] <=  8'h63;        memory[53078] <=  8'h61;        memory[53079] <=  8'h72;        memory[53080] <=  8'h62;        memory[53081] <=  8'h78;        memory[53082] <=  8'h74;        memory[53083] <=  8'h61;        memory[53084] <=  8'h72;        memory[53085] <=  8'h64;        memory[53086] <=  8'h66;        memory[53087] <=  8'h73;        memory[53088] <=  8'h67;        memory[53089] <=  8'h76;        memory[53090] <=  8'h68;        memory[53091] <=  8'h62;        memory[53092] <=  8'h6b;        memory[53093] <=  8'h6a;        memory[53094] <=  8'h6e;        memory[53095] <=  8'h6d;        memory[53096] <=  8'h62;        memory[53097] <=  8'h76;        memory[53098] <=  8'h78;        memory[53099] <=  8'h63;        memory[53100] <=  8'h73;        memory[53101] <=  8'h66;        memory[53102] <=  8'h72;        memory[53103] <=  8'h74;        memory[53104] <=  8'h79;        memory[53105] <=  8'h75;        memory[53106] <=  8'h6a;        memory[53107] <=  8'h6e;        memory[53108] <=  8'h62;        memory[53109] <=  8'h76;        memory[53110] <=  8'h63;        memory[53111] <=  8'h64;        memory[53112] <=  8'h74;        memory[53113] <=  8'h79;        memory[53114] <=  8'h75;        memory[53115] <=  8'h69;        memory[53116] <=  8'h6b;        memory[53117] <=  8'h6d;        memory[53118] <=  8'h6e;        memory[53119] <=  8'h62;        memory[53120] <=  8'h76;        memory[53121] <=  8'h63;        memory[53122] <=  8'h78;        memory[53123] <=  8'h73;        memory[53124] <=  8'h64;        memory[53125] <=  8'h72;        memory[53126] <=  8'h74;        memory[53127] <=  8'h79;        memory[53128] <=  8'h75;        memory[53129] <=  8'h69;        memory[53130] <=  8'h6b;        memory[53131] <=  8'h6d;        memory[53132] <=  8'h6e;        memory[53133] <=  8'h62;        memory[53134] <=  8'h76;        memory[53135] <=  8'h63;        memory[53136] <=  8'h73;        memory[53137] <=  8'h77;        memory[53138] <=  8'h33;        memory[53139] <=  8'h34;        memory[53140] <=  8'h35;        memory[53141] <=  8'h36;        memory[53142] <=  8'h37;        memory[53143] <=  8'h38;        memory[53144] <=  8'h69;        memory[53145] <=  8'h6b;        memory[53146] <=  8'h6d;        memory[53147] <=  8'h6e;        memory[53148] <=  8'h62;        memory[53149] <=  8'h76;        memory[53150] <=  8'h63;        memory[53151] <=  8'h64;        memory[53152] <=  8'h65;        memory[53153] <=  8'h72;        memory[53154] <=  8'h36;        memory[53155] <=  8'h37;        memory[53156] <=  8'h38;        memory[53157] <=  8'h69;        memory[53158] <=  8'h6f;        memory[53159] <=  8'h6b;        memory[53160] <=  8'h6a;        memory[53161] <=  8'h6e;        memory[53162] <=  8'h62;        memory[53163] <=  8'h76;        memory[53164] <=  8'h63;        memory[53165] <=  8'h64;        memory[53166] <=  8'h72;        memory[53167] <=  8'h74;        memory[53168] <=  8'h79;        memory[53169] <=  8'h75;        memory[53170] <=  8'h73;        memory[53171] <=  8'h6a;        memory[53172] <=  8'h63;        memory[53173] <=  8'h6e;        memory[53174] <=  8'h62;        memory[53175] <=  8'h64;        memory[53176] <=  8'h66;        memory[53177] <=  8'h73;        memory[53178] <=  8'h74;        memory[53179] <=  8'h79;        memory[53180] <=  8'h75;        memory[53181] <=  8'h61;        memory[53182] <=  8'h69;        memory[53183] <=  8'h6b;        memory[53184] <=  8'h78;        memory[53185] <=  8'h6d;        memory[53186] <=  8'h6e;        memory[53187] <=  8'h73;        memory[53188] <=  8'h6a;        memory[53189] <=  8'h6f;        memory[53190] <=  8'h64;        memory[53191] <=  8'h6c;        memory[53192] <=  8'h63;        memory[53193] <=  8'h78;        memory[53194] <=  8'h2c;        memory[53195] <=  8'h6d;        memory[53196] <=  8'h73;        memory[53197] <=  8'h6b;        memory[53198] <=  8'h64;        memory[53199] <=  8'h6c;        memory[53200] <=  8'h70;        memory[53201] <=  8'h5b;        memory[53202] <=  8'h3b;        memory[53203] <=  8'h73;        memory[53204] <=  8'h6c;        memory[53205] <=  8'h64;        memory[53206] <=  8'h70;        memory[53207] <=  8'h76;        memory[53208] <=  8'h63;        memory[53209] <=  8'h5b;        memory[53210] <=  8'h78;        memory[53211] <=  8'h76;        memory[53212] <=  8'h63;        memory[53213] <=  8'h5b;        memory[53214] <=  8'h78;        memory[53215] <=  8'h70;        memory[53216] <=  8'h6f;        memory[53217] <=  8'h20;        memory[53218] <=  8'h62;        memory[53219] <=  8'h61;        memory[53220] <=  8'h72;        memory[53221] <=  8'h74;        memory[53222] <=  8'h74;        memory[53223] <=  8'h62;        memory[53224] <=  8'h61;        memory[53225] <=  8'h72;        memory[53226] <=  8'h74;        memory[53227] <=  8'h78;        memory[53228] <=  8'h61;        memory[53229] <=  8'h74;        memory[53230] <=  8'h6b;        memory[53231] <=  8'h73;        memory[53232] <=  8'h68;        memory[53233] <=  8'h63;        memory[53234] <=  8'h66;        memory[53235] <=  8'h69;        memory[53236] <=  8'h77;        memory[53237] <=  8'h68;        memory[53238] <=  8'h61;        memory[53239] <=  8'h69;        memory[53240] <=  8'h6a;        memory[53241] <=  8'h78;        memory[53242] <=  8'h5d;        memory[53243] <=  8'h65;        memory[53244] <=  8'h6b;        memory[53245] <=  8'h6f;        memory[53246] <=  8'h39;        memory[53247] <=  8'h64;        memory[53248] <=  8'h75;        memory[53249] <=  8'h38;        memory[53250] <=  8'h79;        memory[53251] <=  8'h20;        memory[53252] <=  8'h37;        memory[53253] <=  8'h63;        memory[53254] <=  8'h67;        memory[53255] <=  8'h78;        memory[53256] <=  8'h63;        memory[53257] <=  8'h75;        memory[53258] <=  8'h68;        memory[53259] <=  8'h69;        memory[53260] <=  8'h6a;        memory[53261] <=  8'h77;        memory[53262] <=  8'h69;        memory[53263] <=  8'h64;        memory[53264] <=  8'h66;        memory[53265] <=  8'h68;        memory[53266] <=  8'h75;        memory[53267] <=  8'h76;        memory[53268] <=  8'h64;        memory[53269] <=  8'h62;        memory[53270] <=  8'h66;        memory[53271] <=  8'h6a;        memory[53272] <=  8'h6e;        memory[53273] <=  8'h6b;        memory[53274] <=  8'h6a;        memory[53275] <=  8'h65;        memory[53276] <=  8'h38;        memory[53277] <=  8'h66;        memory[53278] <=  8'h37;        memory[53279] <=  8'h67;        memory[53280] <=  8'h79;        memory[53281] <=  8'h76;        memory[53282] <=  8'h63;        memory[53283] <=  8'h68;        memory[53284] <=  8'h69;        memory[53285] <=  8'h6a;        memory[53286] <=  8'h33;        memory[53287] <=  8'h65;        memory[53288] <=  8'h67;        memory[53289] <=  8'h79;        memory[53290] <=  8'h72;        memory[53291] <=  8'h64;        memory[53292] <=  8'h62;        memory[53293] <=  8'h6e;        memory[53294] <=  8'h63;        memory[53295] <=  8'h7a;        memory[53296] <=  8'h6a;        memory[53297] <=  8'h6f;        memory[53298] <=  8'h66;        memory[53299] <=  8'h78;        memory[53300] <=  8'h6a;        memory[53301] <=  8'h69;        memory[53302] <=  8'h63;        memory[53303] <=  8'h68;        memory[53304] <=  8'h62;        memory[53305] <=  8'h6e;        memory[53306] <=  8'h6d;        memory[53307] <=  8'h63;        memory[53308] <=  8'h73;        memory[53309] <=  8'h6c;        memory[53310] <=  8'h6b;        memory[53311] <=  8'h6a;        memory[53312] <=  8'h69;        memory[53313] <=  8'h68;        memory[53314] <=  8'h76;        memory[53315] <=  8'h75;        memory[53316] <=  8'h69;        memory[53317] <=  8'h64;        memory[53318] <=  8'h68;        memory[53319] <=  8'h75;        memory[53320] <=  8'h67;        memory[53321] <=  8'h79;        memory[53322] <=  8'h62;        memory[53323] <=  8'h68;        memory[53324] <=  8'h65;        memory[53325] <=  8'h6a;        memory[53326] <=  8'h72;        memory[53327] <=  8'h6b;        memory[53328] <=  8'h6a;        memory[53329] <=  8'h6f;        memory[53330] <=  8'h64;        memory[53331] <=  8'h67;        memory[53332] <=  8'h69;        memory[53333] <=  8'h75;        memory[53334] <=  8'h69;        memory[53335] <=  8'h67;        memory[53336] <=  8'h76;        memory[53337] <=  8'h79;        memory[53338] <=  8'h75;        memory[53339] <=  8'h67;        memory[53340] <=  8'h78;        memory[53341] <=  8'h68;        memory[53342] <=  8'h63;        memory[53343] <=  8'h20;        memory[53344] <=  8'h20;        memory[53345] <=  8'h20;        memory[53346] <=  8'h78;        memory[53347] <=  8'h76;        memory[53348] <=  8'h20;        memory[53349] <=  8'h63;        memory[53350] <=  8'h78;        memory[53351] <=  8'h67;        memory[53352] <=  8'h79;        memory[53353] <=  8'h63;        memory[53354] <=  8'h75;        memory[53355] <=  8'h68;        memory[53356] <=  8'h6a;        memory[53357] <=  8'h6b;        memory[53358] <=  8'h61;        memory[53359] <=  8'h6c;        memory[53360] <=  8'h78;        memory[53361] <=  8'h76;        memory[53362] <=  8'h70;        memory[53363] <=  8'h6f;        memory[53364] <=  8'h69;        memory[53365] <=  8'h6a;        memory[53366] <=  8'h69;        memory[53367] <=  8'h68;        memory[53368] <=  8'h6a;        memory[53369] <=  8'h62;        memory[53370] <=  8'h77;        memory[53371] <=  8'h65;        memory[53372] <=  8'h6e;        memory[53373] <=  8'h61;        memory[53374] <=  8'h66;        memory[53375] <=  8'h6d;        memory[53376] <=  8'h64;        memory[53377] <=  8'h6b;        memory[53378] <=  8'h6d;        memory[53379] <=  8'h76;        memory[53380] <=  8'h6c;        memory[53381] <=  8'h63;        memory[53382] <=  8'h6f;        memory[53383] <=  8'h64;        memory[53384] <=  8'h69;        memory[53385] <=  8'h75;        memory[53386] <=  8'h68;        memory[53387] <=  8'h73;        memory[53388] <=  8'h66;        memory[53389] <=  8'h65;        memory[53390] <=  8'h62;        memory[53391] <=  8'h6e;        memory[53392] <=  8'h64;        memory[53393] <=  8'h73;        memory[53394] <=  8'h63;        memory[53395] <=  8'h6b;        memory[53396] <=  8'h20;        memory[53397] <=  8'h78;        memory[53398] <=  8'h6a;        memory[53399] <=  8'h78;        memory[53400] <=  8'h63;        memory[53401] <=  8'h73;        memory[53402] <=  8'h64;        memory[53403] <=  8'h66;        memory[53404] <=  8'h6b;        memory[53405] <=  8'h64;        memory[53406] <=  8'h6e;        memory[53407] <=  8'h6d;        memory[53408] <=  8'h64;        memory[53409] <=  8'h73;        memory[53410] <=  8'h63;        memory[53411] <=  8'h6b;        memory[53412] <=  8'h78;        memory[53413] <=  8'h6c;        memory[53414] <=  8'h6f;        memory[53415] <=  8'h66;        memory[53416] <=  8'h6a;        memory[53417] <=  8'h69;        memory[53418] <=  8'h61;        memory[53419] <=  8'h62;        memory[53420] <=  8'h6e;        memory[53421] <=  8'h20;        memory[53422] <=  8'h78;        memory[53423] <=  8'h6b;        memory[53424] <=  8'h6d;        memory[53425] <=  8'h20;        memory[53426] <=  8'h6f;        memory[53427] <=  8'h63;        memory[53428] <=  8'h76;        memory[53429] <=  8'h73;        memory[53430] <=  8'h64;        memory[53431] <=  8'h69;        memory[53432] <=  8'h66;        memory[53433] <=  8'h68;        memory[53434] <=  8'h65;        memory[53435] <=  8'h71;        memory[53436] <=  8'h6a;        memory[53437] <=  8'h77;        memory[53438] <=  8'h62;        memory[53439] <=  8'h65;        memory[53440] <=  8'h6e;        memory[53441] <=  8'h20;        memory[53442] <=  8'h6d;        memory[53443] <=  8'h64;        memory[53444] <=  8'h73;        memory[53445] <=  8'h6c;        memory[53446] <=  8'h76;        memory[53447] <=  8'h6b;        memory[53448] <=  8'h63;        memory[53449] <=  8'h78;        memory[53450] <=  8'h20;        memory[53451] <=  8'h6f;        memory[53452] <=  8'h78;        memory[53453] <=  8'h69;        memory[53454] <=  8'h63;        memory[53455] <=  8'h6a;        memory[53456] <=  8'h76;        memory[53457] <=  8'h64;        memory[53458] <=  8'h66;        memory[53459] <=  8'h65;        memory[53460] <=  8'h71;        memory[53461] <=  8'h6e;        memory[53462] <=  8'h20;        memory[53463] <=  8'h64;        memory[53464] <=  8'h6d;        memory[53465] <=  8'h73;        memory[53466] <=  8'h6c;        memory[53467] <=  8'h63;        memory[53468] <=  8'h78;        memory[53469] <=  8'h6b;        memory[53470] <=  8'h20;        memory[53471] <=  8'h6f;        memory[53472] <=  8'h78;        memory[53473] <=  8'h63;        memory[53474] <=  8'h76;        memory[53475] <=  8'h6a;        memory[53476] <=  8'h64;        memory[53477] <=  8'h62;        memory[53478] <=  8'h71;        memory[53479] <=  8'h77;        memory[53480] <=  8'h65;        memory[53481] <=  8'h6e;        memory[53482] <=  8'h6d;        memory[53483] <=  8'h64;        memory[53484] <=  8'h6c;        memory[53485] <=  8'h73;        memory[53486] <=  8'h2c;        memory[53487] <=  8'h76;        memory[53488] <=  8'h63;        memory[53489] <=  8'h78;        memory[53490] <=  8'h20;        memory[53491] <=  8'h63;        memory[53492] <=  8'h6f;        memory[53493] <=  8'h69;        memory[53494] <=  8'h76;        memory[53495] <=  8'h68;        memory[53496] <=  8'h73;        memory[53497] <=  8'h64;        memory[53498] <=  8'h62;        memory[53499] <=  8'h71;        memory[53500] <=  8'h77;        memory[53501] <=  8'h65;        memory[53502] <=  8'h6e;        memory[53503] <=  8'h64;        memory[53504] <=  8'h6b;        memory[53505] <=  8'h73;        memory[53506] <=  8'h76;        memory[53507] <=  8'h6f;        memory[53508] <=  8'h63;        memory[53509] <=  8'h20;        memory[53510] <=  8'h76;        memory[53511] <=  8'h69;        memory[53512] <=  8'h75;        memory[53513] <=  8'h69;        memory[53514] <=  8'h68;        memory[53515] <=  8'h63;        memory[53516] <=  8'h78;        memory[53517] <=  8'h69;        memory[53518] <=  8'h6f;        memory[53519] <=  8'h76;        memory[53520] <=  8'h73;        memory[53521] <=  8'h64;        memory[53522] <=  8'h61;        memory[53523] <=  8'h64;        memory[53524] <=  8'h6e;        memory[53525] <=  8'h77;        memory[53526] <=  8'h71;        memory[53527] <=  8'h6b;        memory[53528] <=  8'h6c;        memory[53529] <=  8'h73;        memory[53530] <=  8'h76;        memory[53531] <=  8'h6e;        memory[53532] <=  8'h62;        memory[53533] <=  8'h20;        memory[53534] <=  8'h64;        memory[53535] <=  8'h66;        memory[53536] <=  8'h6a;        memory[53537] <=  8'h6b;        memory[53538] <=  8'h71;        memory[53539] <=  8'h64;        memory[53540] <=  8'h77;        memory[53541] <=  8'h65;        memory[53542] <=  8'h6e;        memory[53543] <=  8'h62;        memory[53544] <=  8'h20;        memory[53545] <=  8'h64;        memory[53546] <=  8'h73;        memory[53547] <=  8'h76;        memory[53548] <=  8'h68;        memory[53549] <=  8'h64;        memory[53550] <=  8'h61;        memory[53551] <=  8'h71;        memory[53552] <=  8'h77;        memory[53553] <=  8'h6a;        memory[53554] <=  8'h65;        memory[53555] <=  8'h6e;        memory[53556] <=  8'h64;        memory[53557] <=  8'h20;        memory[53558] <=  8'h61;        memory[53559] <=  8'h63;        memory[53560] <=  8'h62;        memory[53561] <=  8'h68;        memory[53562] <=  8'h64;        memory[53563] <=  8'h61;        memory[53564] <=  8'h77;        memory[53565] <=  8'h71;        memory[53566] <=  8'h6e;        memory[53567] <=  8'h20;        memory[53568] <=  8'h62;        memory[53569] <=  8'h73;        memory[53570] <=  8'h76;        memory[53571] <=  8'h61;        memory[53572] <=  8'h67;        memory[53573] <=  8'h76;        memory[53574] <=  8'h68;        memory[53575] <=  8'h67;        memory[53576] <=  8'h61;        memory[53577] <=  8'h73;        memory[53578] <=  8'h6a;        memory[53579] <=  8'h6b;        memory[53580] <=  8'h63;        memory[53581] <=  8'h78;        memory[53582] <=  8'h76;        memory[53583] <=  8'h6e;        memory[53584] <=  8'h73;        memory[53585] <=  8'h64;        memory[53586] <=  8'h20;        memory[53587] <=  8'h66;        memory[53588] <=  8'h62;        memory[53589] <=  8'h64;        memory[53590] <=  8'h61;        memory[53591] <=  8'h73;        memory[53592] <=  8'h76;        memory[53593] <=  8'h67;        memory[53594] <=  8'h63;        memory[53595] <=  8'h79;        memory[53596] <=  8'h7a;        memory[53597] <=  8'h78;        memory[53598] <=  8'h79;        memory[53599] <=  8'h75;        memory[53600] <=  8'h20;        memory[53601] <=  8'h69;        memory[53602] <=  8'h6a;        memory[53603] <=  8'h64;        memory[53604] <=  8'h66;        memory[53605] <=  8'h6b;        memory[53606] <=  8'h61;        memory[53607] <=  8'h64;        memory[53608] <=  8'h63;        memory[53609] <=  8'h78;        memory[53610] <=  8'h68;        memory[53611] <=  8'h20;        memory[53612] <=  8'h67;        memory[53613] <=  8'h61;        memory[53614] <=  8'h68;        memory[53615] <=  8'h75;        memory[53616] <=  8'h64;        memory[53617] <=  8'h73;        memory[53618] <=  8'h69;        memory[53619] <=  8'h6a;        memory[53620] <=  8'h61;        memory[53621] <=  8'h6b;        memory[53622] <=  8'h63;        memory[53623] <=  8'h62;        memory[53624] <=  8'h61;        memory[53625] <=  8'h72;        memory[53626] <=  8'h73;        memory[53627] <=  8'h68;        memory[53628] <=  8'h64;        memory[53629] <=  8'h66;        memory[53630] <=  8'h67;        memory[53631] <=  8'h73;        memory[53632] <=  8'h68;        memory[53633] <=  8'h64;        memory[53634] <=  8'h66;        memory[53635] <=  8'h68;        memory[53636] <=  8'h64;        memory[53637] <=  8'h6a;        memory[53638] <=  8'h68;        memory[53639] <=  8'h62;        memory[53640] <=  8'h67;        memory[53641] <=  8'h63;        memory[53642] <=  8'h61;        memory[53643] <=  8'h66;        memory[53644] <=  8'h73;        memory[53645] <=  8'h79;        memory[53646] <=  8'h67;        memory[53647] <=  8'h6b;        memory[53648] <=  8'h75;        memory[53649] <=  8'h64;        memory[53650] <=  8'h68;        memory[53651] <=  8'h62;        memory[53652] <=  8'h77;        memory[53653] <=  8'h76;        memory[53654] <=  8'h67;        memory[53655] <=  8'h61;        memory[53656] <=  8'h66;        memory[53657] <=  8'h64;        memory[53658] <=  8'h74;        memory[53659] <=  8'h75;        memory[53660] <=  8'h66;        memory[53661] <=  8'h79;        memory[53662] <=  8'h67;        memory[53663] <=  8'h69;        memory[53664] <=  8'h75;        memory[53665] <=  8'h68;        memory[53666] <=  8'h6c;        memory[53667] <=  8'h6a;        memory[53668] <=  8'h62;        memory[53669] <=  8'h6b;        memory[53670] <=  8'h68;        memory[53671] <=  8'h76;        memory[53672] <=  8'h67;        memory[53673] <=  8'h63;        memory[53674] <=  8'h66;        memory[53675] <=  8'h78;        memory[53676] <=  8'h64;        memory[53677] <=  8'h74;        memory[53678] <=  8'h75;        memory[53679] <=  8'h79;        memory[53680] <=  8'h69;        memory[53681] <=  8'h75;        memory[53682] <=  8'h68;        memory[53683] <=  8'h6c;        memory[53684] <=  8'h6a;        memory[53685] <=  8'h6b;        memory[53686] <=  8'h67;        memory[53687] <=  8'h6a;        memory[53688] <=  8'h63;        memory[53689] <=  8'h66;        memory[53690] <=  8'h68;        memory[53691] <=  8'h64;        memory[53692] <=  8'h67;        memory[53693] <=  8'h72;        memory[53694] <=  8'h79;        memory[53695] <=  8'h74;        memory[53696] <=  8'h66;        memory[53697] <=  8'h75;        memory[53698] <=  8'h79;        memory[53699] <=  8'h69;        memory[53700] <=  8'h68;        memory[53701] <=  8'h6c;        memory[53702] <=  8'h62;        memory[53703] <=  8'h6d;        memory[53704] <=  8'h76;        memory[53705] <=  8'h6e;        memory[53706] <=  8'h63;        memory[53707] <=  8'h66;        memory[53708] <=  8'h68;        memory[53709] <=  8'h64;        memory[53710] <=  8'h74;        memory[53711] <=  8'h75;        memory[53712] <=  8'h67;        memory[53713] <=  8'h79;        memory[53714] <=  8'h69;        memory[53715] <=  8'h68;        memory[53716] <=  8'h75;        memory[53717] <=  8'h6a;        memory[53718] <=  8'h6c;        memory[53719] <=  8'h62;        memory[53720] <=  8'h6d;        memory[53721] <=  8'h76;        memory[53722] <=  8'h6e;        memory[53723] <=  8'h63;        memory[53724] <=  8'h66;        memory[53725] <=  8'h68;        memory[53726] <=  8'h67;        memory[53727] <=  8'h79;        memory[53728] <=  8'h68;        memory[53729] <=  8'h75;        memory[53730] <=  8'h6a;        memory[53731] <=  8'h6e;        memory[53732] <=  8'h2c;        memory[53733] <=  8'h62;        memory[53734] <=  8'h6e;        memory[53735] <=  8'h6d;        memory[53736] <=  8'h76;        memory[53737] <=  8'h6e;        memory[53738] <=  8'h63;        memory[53739] <=  8'h66;        memory[53740] <=  8'h68;        memory[53741] <=  8'h74;        memory[53742] <=  8'h79;        memory[53743] <=  8'h69;        memory[53744] <=  8'h75;        memory[53745] <=  8'h6c;        memory[53746] <=  8'h6a;        memory[53747] <=  8'h62;        memory[53748] <=  8'h6d;        memory[53749] <=  8'h76;        memory[53750] <=  8'h6e;        memory[53751] <=  8'h63;        memory[53752] <=  8'h66;        memory[53753] <=  8'h74;        memory[53754] <=  8'h75;        memory[53755] <=  8'h79;        memory[53756] <=  8'h69;        memory[53757] <=  8'h68;        memory[53758] <=  8'h6b;        memory[53759] <=  8'h62;        memory[53760] <=  8'h76;        memory[53761] <=  8'h63;        memory[53762] <=  8'h66;        memory[53763] <=  8'h67;        memory[53764] <=  8'h74;        memory[53765] <=  8'h75;        memory[53766] <=  8'h79;        memory[53767] <=  8'h69;        memory[53768] <=  8'h75;        memory[53769] <=  8'h68;        memory[53770] <=  8'h6a;        memory[53771] <=  8'h6b;        memory[53772] <=  8'h62;        memory[53773] <=  8'h76;        memory[53774] <=  8'h63;        memory[53775] <=  8'h66;        memory[53776] <=  8'h74;        memory[53777] <=  8'h75;        memory[53778] <=  8'h79;        memory[53779] <=  8'h69;        memory[53780] <=  8'h75;        memory[53781] <=  8'h6a;        memory[53782] <=  8'h6b;        memory[53783] <=  8'h6e;        memory[53784] <=  8'h62;        memory[53785] <=  8'h76;        memory[53786] <=  8'h67;        memory[53787] <=  8'h66;        memory[53788] <=  8'h74;        memory[53789] <=  8'h79;        memory[53790] <=  8'h75;        memory[53791] <=  8'h75;        memory[53792] <=  8'h69;        memory[53793] <=  8'h6a;        memory[53794] <=  8'h6b;        memory[53795] <=  8'h68;        memory[53796] <=  8'h62;        memory[53797] <=  8'h6a;        memory[53798] <=  8'h67;        memory[53799] <=  8'h68;        memory[53800] <=  8'h66;        memory[53801] <=  8'h79;        memory[53802] <=  8'h74;        memory[53803] <=  8'h79;        memory[53804] <=  8'h69;        memory[53805] <=  8'h75;        memory[53806] <=  8'h64;        memory[53807] <=  8'h6a;        memory[53808] <=  8'h6b;        memory[53809] <=  8'h68;        memory[53810] <=  8'h63;        memory[53811] <=  8'h7a;        memory[53812] <=  8'h67;        memory[53813] <=  8'h68;        memory[53814] <=  8'h74;        memory[53815] <=  8'h75;        memory[53816] <=  8'h79;        memory[53817] <=  8'h69;        memory[53818] <=  8'h61;        memory[53819] <=  8'h73;        memory[53820] <=  8'h75;        memory[53821] <=  8'h6a;        memory[53822] <=  8'h6b;        memory[53823] <=  8'h62;        memory[53824] <=  8'h6e;        memory[53825] <=  8'h61;        memory[53826] <=  8'h76;        memory[53827] <=  8'h63;        memory[53828] <=  8'h66;        memory[53829] <=  8'h68;        memory[53830] <=  8'h75;        memory[53831] <=  8'h61;        memory[53832] <=  8'h73;        memory[53833] <=  8'h79;        memory[53834] <=  8'h64;        memory[53835] <=  8'h75;        memory[53836] <=  8'h69;        memory[53837] <=  8'h6a;        memory[53838] <=  8'h61;        memory[53839] <=  8'h6b;        memory[53840] <=  8'h62;        memory[53841] <=  8'h63;        memory[53842] <=  8'h78;        memory[53843] <=  8'h68;        memory[53844] <=  8'h67;        memory[53845] <=  8'h79;        memory[53846] <=  8'h75;        memory[53847] <=  8'h7a;        memory[53848] <=  8'h63;        memory[53849] <=  8'h61;        memory[53850] <=  8'h73;        memory[53851] <=  8'h69;        memory[53852] <=  8'h75;        memory[53853] <=  8'h6f;        memory[53854] <=  8'h69;        memory[53855] <=  8'h6a;        memory[53856] <=  8'h61;        memory[53857] <=  8'h6c;        memory[53858] <=  8'h63;        memory[53859] <=  8'h78;        memory[53860] <=  8'h62;        memory[53861] <=  8'h63;        memory[53862] <=  8'h20;        memory[53863] <=  8'h6e;        memory[53864] <=  8'h76;        memory[53865] <=  8'h63;        memory[53866] <=  8'h61;        memory[53867] <=  8'h64;        memory[53868] <=  8'h73;        memory[53869] <=  8'h67;        memory[53870] <=  8'h79;        memory[53871] <=  8'h68;        memory[53872] <=  8'h75;        memory[53873] <=  8'h61;        memory[53874] <=  8'h6a;        memory[53875] <=  8'h6b;        memory[53876] <=  8'h78;        memory[53877] <=  8'h62;        memory[53878] <=  8'h20;        memory[53879] <=  8'h6e;        memory[53880] <=  8'h76;        memory[53881] <=  8'h63;        memory[53882] <=  8'h61;        memory[53883] <=  8'h73;        memory[53884] <=  8'h67;        memory[53885] <=  8'h68;        memory[53886] <=  8'h75;        memory[53887] <=  8'h6a;        memory[53888] <=  8'h6c;        memory[53889] <=  8'h6b;        memory[53890] <=  8'h63;        memory[53891] <=  8'h78;        memory[53892] <=  8'h20;        memory[53893] <=  8'h6a;        memory[53894] <=  8'h6b;        memory[53895] <=  8'h68;        memory[53896] <=  8'h61;        memory[53897] <=  8'h73;        memory[53898] <=  8'h76;        memory[53899] <=  8'h64;        memory[53900] <=  8'h6e;        memory[53901] <=  8'h20;        memory[53902] <=  8'h62;        memory[53903] <=  8'h6e;        memory[53904] <=  8'h6d;        memory[53905] <=  8'h6b;        memory[53906] <=  8'h77;        memory[53907] <=  8'h64;        memory[53908] <=  8'h6f;        memory[53909] <=  8'h77;        memory[53910] <=  8'h69;        memory[53911] <=  8'h6f;        memory[53912] <=  8'h75;        memory[53913] <=  8'h69;        memory[53914] <=  8'h68;        memory[53915] <=  8'h62;        memory[53916] <=  8'h6e;        memory[53917] <=  8'h6b;        memory[53918] <=  8'h77;        memory[53919] <=  8'h69;        memory[53920] <=  8'h6f;        memory[53921] <=  8'h75;        memory[53922] <=  8'h71;        memory[53923] <=  8'h69;        memory[53924] <=  8'h79;        memory[53925] <=  8'h67;        memory[53926] <=  8'h6a;        memory[53927] <=  8'h64;        memory[53928] <=  8'h61;        memory[53929] <=  8'h76;        memory[53930] <=  8'h62;        memory[53931] <=  8'h6e;        memory[53932] <=  8'h6b;        memory[53933] <=  8'h6f;        memory[53934] <=  8'h70;        memory[53935] <=  8'h64;        memory[53936] <=  8'h76;        memory[53937] <=  8'h69;        memory[53938] <=  8'h6f;        memory[53939] <=  8'h75;        memory[53940] <=  8'h69;        memory[53941] <=  8'h48;        memory[53942] <=  8'h42;        memory[53943] <=  8'h6b;        memory[53944] <=  8'h64;        memory[53945] <=  8'h6e;        memory[53946] <=  8'h6c;        memory[53947] <=  8'h71;        memory[53948] <=  8'h6b;        memory[53949] <=  8'h6d;        memory[53950] <=  8'h6a;        memory[53951] <=  8'h70;        memory[53952] <=  8'h69;        memory[53953] <=  8'h6f;        memory[53954] <=  8'h68;        memory[53955] <=  8'h65;        memory[53956] <=  8'h66;        memory[53957] <=  8'h75;        memory[53958] <=  8'h67;        memory[53959] <=  8'h69;        memory[53960] <=  8'h73;        memory[53961] <=  8'h61;        memory[53962] <=  8'h62;        memory[53963] <=  8'h64;        memory[53964] <=  8'h6b;        memory[53965] <=  8'h6a;        memory[53966] <=  8'h6b;        memory[53967] <=  8'h6c;        memory[53968] <=  8'h6a;        memory[53969] <=  8'h69;        memory[53970] <=  8'h73;        memory[53971] <=  8'h6f;        memory[53972] <=  8'h71;        memory[53973] <=  8'h68;        memory[53974] <=  8'h77;        memory[53975] <=  8'h67;        memory[53976] <=  8'h69;        memory[53977] <=  8'h79;        memory[53978] <=  8'h6a;        memory[53979] <=  8'h64;        memory[53980] <=  8'h76;        memory[53981] <=  8'h62;        memory[53982] <=  8'h6e;        memory[53983] <=  8'h61;        memory[53984] <=  8'h73;        memory[53985] <=  8'h66;        memory[53986] <=  8'h6c;        memory[53987] <=  8'h6b;        memory[53988] <=  8'h64;        memory[53989] <=  8'h6a;        memory[53990] <=  8'h68;        memory[53991] <=  8'h63;        memory[53992] <=  8'h67;        memory[53993] <=  8'h6a;        memory[53994] <=  8'h76;        memory[53995] <=  8'h73;        memory[53996] <=  8'h64;        memory[53997] <=  8'h62;        memory[53998] <=  8'h62;        memory[53999] <=  8'h61;        memory[54000] <=  8'h72;        memory[54001] <=  8'h62;        memory[54002] <=  8'h62;        memory[54003] <=  8'h73;        memory[54004] <=  8'h62;        memory[54005] <=  8'h67;        memory[54006] <=  8'h73;        memory[54007] <=  8'h66;        memory[54008] <=  8'h67;        memory[54009] <=  8'h61;        memory[54010] <=  8'h68;        memory[54011] <=  8'h66;        memory[54012] <=  8'h73;        memory[54013] <=  8'h68;        memory[54014] <=  8'h61;        memory[54015] <=  8'h66;        memory[54016] <=  8'h73;        memory[54017] <=  8'h66;        memory[54018] <=  8'h68;        memory[54019] <=  8'h61;        memory[54020] <=  8'h69;        memory[54021] <=  8'h64;        memory[54022] <=  8'h75;        memory[54023] <=  8'h67;        memory[54024] <=  8'h64;        memory[54025] <=  8'h77;        memory[54026] <=  8'h62;        memory[54027] <=  8'h61;        memory[54028] <=  8'h62;        memory[54029] <=  8'h72;        memory[54030] <=  8'h62;        memory[54031] <=  8'h61;        memory[54032] <=  8'h62;        memory[54033] <=  8'h62;        memory[54034] <=  8'h74;        memory[54035] <=  8'h62;        memory[54036] <=  8'h62;        memory[54037] <=  8'h62;        memory[54038] <=  8'h62;        memory[54039] <=  8'h62;        memory[54040] <=  8'h62;        memory[54041] <=  8'h62;        memory[54042] <=  8'h62;        memory[54043] <=  8'h61;        memory[54044] <=  8'h62;        memory[54045] <=  8'h62;        memory[54046] <=  8'h72;        memory[54047] <=  8'h74;        memory[54048] <=  8'h62;        memory[54049] <=  8'h62;        memory[54050] <=  8'h61;        memory[54051] <=  8'h62;        memory[54052] <=  8'h72;        memory[54053] <=  8'h62;        memory[54054] <=  8'h74;        memory[54055] <=  8'h62;        memory[54056] <=  8'h62;        memory[54057] <=  8'h62;        memory[54058] <=  8'h63;        memory[54059] <=  8'h61;        memory[54060] <=  8'h72;        memory[54061] <=  8'h74;        memory[54062] <=  8'h73;        memory[54063] <=  8'h62;        memory[54064] <=  8'h61;        memory[54065] <=  8'h72;        memory[54066] <=  8'h74;        memory[54067] <=  8'h74;        memory[54068] <=  8'h62;        memory[54069] <=  8'h61;        memory[54070] <=  8'h72;        memory[54071] <=  8'h74;        memory[54072] <=  8'h78;        memory[54073] <=  8'h61;        memory[54074] <=  8'h74;        memory[54075] <=  8'h6b;        memory[54076] <=  8'h73;        memory[54077] <=  8'h68;        memory[54078] <=  8'h63;        memory[54079] <=  8'h66;        memory[54080] <=  8'h69;        memory[54081] <=  8'h77;        memory[54082] <=  8'h68;        memory[54083] <=  8'h61;        memory[54084] <=  8'h74;        memory[54085] <=  8'h61;        memory[54086] <=  8'h6e;        memory[54087] <=  8'h61;        memory[54088] <=  8'h62;        memory[54089] <=  8'h61;        memory[54090] <=  8'h63;        memory[54091] <=  8'h61;        memory[54092] <=  8'h74;        memory[54093] <=  8'h61;        memory[54094] <=  8'h62;        memory[54095] <=  8'h61;        memory[54096] <=  8'h72;        memory[54097] <=  8'h63;        memory[54098] <=  8'h61;        memory[54099] <=  8'h68;        memory[54100] <=  8'h64;        memory[54101] <=  8'h75;        memory[54102] <=  8'h63;        memory[54103] <=  8'h74;        memory[54104] <=  8'h61;        memory[54105] <=  8'h64;        memory[54106] <=  8'h61;        memory[54107] <=  8'h61;        memory[54108] <=  8'h63;        memory[54109] <=  8'h61;        memory[54110] <=  8'h72;        memory[54111] <=  8'h63;        memory[54112] <=  8'h74;        memory[54113] <=  8'h72;        memory[54114] <=  8'h63;        memory[54115] <=  8'h61;        memory[54116] <=  8'h74;        memory[54117] <=  8'h72;        memory[54118] <=  8'h63;        memory[54119] <=  8'h61;        memory[54120] <=  8'h74;        memory[54121] <=  8'h63;        memory[54122] <=  8'h62;        memory[54123] <=  8'h61;        memory[54124] <=  8'h74;        memory[54125] <=  8'h62;        memory[54126] <=  8'h72;        memory[54127] <=  8'h63;        memory[54128] <=  8'h61;        memory[54129] <=  8'h74;        memory[54130] <=  8'h72;        memory[54131] <=  8'h6e;        memory[54132] <=  8'h62;        memory[54133] <=  8'h61;        memory[54134] <=  8'h63;        memory[54135] <=  8'h61;        memory[54136] <=  8'h74;        memory[54137] <=  8'h79;        memory[54138] <=  8'h73;        memory[54139] <=  8'h6e;        memory[54140] <=  8'h63;        memory[54141] <=  8'h74;        memory[54142] <=  8'h61;        memory[54143] <=  8'h6e;        memory[54144] <=  8'h62;        memory[54145] <=  8'h61;        memory[54146] <=  8'h63;        memory[54147] <=  8'h72;        memory[54148] <=  8'h6e;        memory[54149] <=  8'h74;        memory[54150] <=  8'h61;        memory[54151] <=  8'h62;        memory[54152] <=  8'h74;        memory[54153] <=  8'h6e;        memory[54154] <=  8'h61;        memory[54155] <=  8'h72;        memory[54156] <=  8'h62;        memory[54157] <=  8'h78;        memory[54158] <=  8'h74;        memory[54159] <=  8'h61;        memory[54160] <=  8'h72;        memory[54161] <=  8'h62;        memory[54162] <=  8'h61;        memory[54163] <=  8'h72;        memory[54164] <=  8'h74;        memory[54165] <=  8'h74;        memory[54166] <=  8'h62;        memory[54167] <=  8'h61;        memory[54168] <=  8'h72;        memory[54169] <=  8'h74;        memory[54170] <=  8'h78;        memory[54171] <=  8'h61;        memory[54172] <=  8'h74;        memory[54173] <=  8'h6b;        memory[54174] <=  8'h73;        memory[54175] <=  8'h68;        memory[54176] <=  8'h63;        memory[54177] <=  8'h66;        memory[54178] <=  8'h69;        memory[54179] <=  8'h77;        memory[54180] <=  8'h68;        memory[54181] <=  8'h61;        memory[54182] <=  8'h74;        memory[54183] <=  8'h61;        memory[54184] <=  8'h6e;        memory[54185] <=  8'h61;        memory[54186] <=  8'h62;        memory[54187] <=  8'h61;        memory[54188] <=  8'h63;        memory[54189] <=  8'h61;        memory[54190] <=  8'h74;        memory[54191] <=  8'h61;        memory[54192] <=  8'h62;        memory[54193] <=  8'h61;        memory[54194] <=  8'h72;        memory[54195] <=  8'h63;        memory[54196] <=  8'h61;        memory[54197] <=  8'h68;        memory[54198] <=  8'h64;        memory[54199] <=  8'h75;        memory[54200] <=  8'h63;        memory[54201] <=  8'h74;        memory[54202] <=  8'h61;        memory[54203] <=  8'h64;        memory[54204] <=  8'h61;        memory[54205] <=  8'h61;        memory[54206] <=  8'h63;        memory[54207] <=  8'h61;        memory[54208] <=  8'h72;        memory[54209] <=  8'h63;        memory[54210] <=  8'h74;        memory[54211] <=  8'h72;        memory[54212] <=  8'h63;        memory[54213] <=  8'h61;        memory[54214] <=  8'h74;        memory[54215] <=  8'h72;        memory[54216] <=  8'h63;        memory[54217] <=  8'h61;        memory[54218] <=  8'h74;        memory[54219] <=  8'h63;        memory[54220] <=  8'h62;        memory[54221] <=  8'h61;        memory[54222] <=  8'h74;        memory[54223] <=  8'h62;        memory[54224] <=  8'h72;        memory[54225] <=  8'h63;        memory[54226] <=  8'h61;        memory[54227] <=  8'h74;        memory[54228] <=  8'h72;        memory[54229] <=  8'h6e;        memory[54230] <=  8'h62;        memory[54231] <=  8'h61;        memory[54232] <=  8'h63;        memory[54233] <=  8'h61;        memory[54234] <=  8'h74;        memory[54235] <=  8'h79;        memory[54236] <=  8'h73;        memory[54237] <=  8'h6e;        memory[54238] <=  8'h63;        memory[54239] <=  8'h74;        memory[54240] <=  8'h61;        memory[54241] <=  8'h6e;        memory[54242] <=  8'h62;        memory[54243] <=  8'h61;        memory[54244] <=  8'h63;        memory[54245] <=  8'h72;        memory[54246] <=  8'h6e;        memory[54247] <=  8'h74;        memory[54248] <=  8'h61;        memory[54249] <=  8'h62;        memory[54250] <=  8'h74;        memory[54251] <=  8'h6e;        memory[54252] <=  8'h61;        memory[54253] <=  8'h72;        memory[54254] <=  8'h62;        memory[54255] <=  8'h78;        memory[54256] <=  8'h74;        memory[54257] <=  8'h61;        memory[54258] <=  8'h72;        memory[54259] <=  8'h62;        memory[54260] <=  8'h61;        memory[54261] <=  8'h72;        memory[54262] <=  8'h74;        memory[54263] <=  8'h74;        memory[54264] <=  8'h62;        memory[54265] <=  8'h61;        memory[54266] <=  8'h72;        memory[54267] <=  8'h74;        memory[54268] <=  8'h78;        memory[54269] <=  8'h61;        memory[54270] <=  8'h74;        memory[54271] <=  8'h6b;        memory[54272] <=  8'h73;        memory[54273] <=  8'h68;        memory[54274] <=  8'h63;        memory[54275] <=  8'h66;        memory[54276] <=  8'h69;        memory[54277] <=  8'h77;        memory[54278] <=  8'h68;        memory[54279] <=  8'h61;        memory[54280] <=  8'h74;        memory[54281] <=  8'h61;        memory[54282] <=  8'h6e;        memory[54283] <=  8'h61;        memory[54284] <=  8'h62;        memory[54285] <=  8'h61;        memory[54286] <=  8'h63;        memory[54287] <=  8'h61;        memory[54288] <=  8'h74;        memory[54289] <=  8'h61;        memory[54290] <=  8'h62;        memory[54291] <=  8'h61;        memory[54292] <=  8'h72;        memory[54293] <=  8'h63;        memory[54294] <=  8'h61;        memory[54295] <=  8'h68;        memory[54296] <=  8'h64;        memory[54297] <=  8'h75;        memory[54298] <=  8'h63;        memory[54299] <=  8'h74;        memory[54300] <=  8'h61;        memory[54301] <=  8'h64;        memory[54302] <=  8'h61;        memory[54303] <=  8'h61;        memory[54304] <=  8'h63;        memory[54305] <=  8'h61;        memory[54306] <=  8'h72;        memory[54307] <=  8'h63;        memory[54308] <=  8'h74;        memory[54309] <=  8'h72;        memory[54310] <=  8'h63;        memory[54311] <=  8'h61;        memory[54312] <=  8'h74;        memory[54313] <=  8'h72;        memory[54314] <=  8'h63;        memory[54315] <=  8'h61;        memory[54316] <=  8'h74;        memory[54317] <=  8'h63;        memory[54318] <=  8'h62;        memory[54319] <=  8'h61;        memory[54320] <=  8'h74;        memory[54321] <=  8'h62;        memory[54322] <=  8'h72;        memory[54323] <=  8'h63;        memory[54324] <=  8'h61;        memory[54325] <=  8'h74;        memory[54326] <=  8'h72;        memory[54327] <=  8'h6e;        memory[54328] <=  8'h62;        memory[54329] <=  8'h61;        memory[54330] <=  8'h63;        memory[54331] <=  8'h61;        memory[54332] <=  8'h74;        memory[54333] <=  8'h79;        memory[54334] <=  8'h73;        memory[54335] <=  8'h6e;        memory[54336] <=  8'h63;        memory[54337] <=  8'h74;        memory[54338] <=  8'h61;        memory[54339] <=  8'h6e;        memory[54340] <=  8'h62;        memory[54341] <=  8'h61;        memory[54342] <=  8'h63;        memory[54343] <=  8'h72;        memory[54344] <=  8'h6e;        memory[54345] <=  8'h74;        memory[54346] <=  8'h61;        memory[54347] <=  8'h62;        memory[54348] <=  8'h74;        memory[54349] <=  8'h6e;        memory[54350] <=  8'h61;        memory[54351] <=  8'h72;        memory[54352] <=  8'h62;        memory[54353] <=  8'h78;        memory[54354] <=  8'h74;        memory[54355] <=  8'h61;        memory[54356] <=  8'h72;        memory[54357] <=  8'h5d;        memory[54358] <=  8'h5d;        memory[54359] <=  8'h65;        memory[54360] <=  8'h66;        memory[54361] <=  8'h77;        memory[54362] <=  8'h65;        memory[54363] <=  8'h5d;        memory[54364] <=  8'h65;        memory[54365] <=  8'h67;        memory[54366] <=  8'h73;        memory[54367] <=  8'h67;        memory[54368] <=  8'h66;        memory[54369] <=  8'h62;        memory[54370] <=  8'h61;        memory[54371] <=  8'h72;        memory[54372] <=  8'h74;        memory[54373] <=  8'h74;        memory[54374] <=  8'h62;        memory[54375] <=  8'h61;        memory[54376] <=  8'h72;        memory[54377] <=  8'h74;        memory[54378] <=  8'h78;        memory[54379] <=  8'h61;        memory[54380] <=  8'h74;        memory[54381] <=  8'h6b;        memory[54382] <=  8'h73;        memory[54383] <=  8'h68;        memory[54384] <=  8'h63;        memory[54385] <=  8'h66;        memory[54386] <=  8'h69;        memory[54387] <=  8'h77;        memory[54388] <=  8'h68;        memory[54389] <=  8'h61;        memory[54390] <=  8'h74;        memory[54391] <=  8'h61;        memory[54392] <=  8'h6e;        memory[54393] <=  8'h61;        memory[54394] <=  8'h62;        memory[54395] <=  8'h61;        memory[54396] <=  8'h63;        memory[54397] <=  8'h61;        memory[54398] <=  8'h74;        memory[54399] <=  8'h61;        memory[54400] <=  8'h62;        memory[54401] <=  8'h61;        memory[54402] <=  8'h72;        memory[54403] <=  8'h63;        memory[54404] <=  8'h61;        memory[54405] <=  8'h68;        memory[54406] <=  8'h64;        memory[54407] <=  8'h75;        memory[54408] <=  8'h63;        memory[54409] <=  8'h74;        memory[54410] <=  8'h61;        memory[54411] <=  8'h64;        memory[54412] <=  8'h61;        memory[54413] <=  8'h61;        memory[54414] <=  8'h63;        memory[54415] <=  8'h61;        memory[54416] <=  8'h72;        memory[54417] <=  8'h63;        memory[54418] <=  8'h74;        memory[54419] <=  8'h72;        memory[54420] <=  8'h63;        memory[54421] <=  8'h61;        memory[54422] <=  8'h74;        memory[54423] <=  8'h72;        memory[54424] <=  8'h63;        memory[54425] <=  8'h61;        memory[54426] <=  8'h74;        memory[54427] <=  8'h63;        memory[54428] <=  8'h62;        memory[54429] <=  8'h61;        memory[54430] <=  8'h74;        memory[54431] <=  8'h62;        memory[54432] <=  8'h72;        memory[54433] <=  8'h63;        memory[54434] <=  8'h61;        memory[54435] <=  8'h74;        memory[54436] <=  8'h72;        memory[54437] <=  8'h6e;        memory[54438] <=  8'h62;        memory[54439] <=  8'h61;        memory[54440] <=  8'h63;        memory[54441] <=  8'h61;        memory[54442] <=  8'h74;        memory[54443] <=  8'h79;        memory[54444] <=  8'h73;        memory[54445] <=  8'h6e;        memory[54446] <=  8'h63;        memory[54447] <=  8'h74;        memory[54448] <=  8'h61;        memory[54449] <=  8'h6e;        memory[54450] <=  8'h62;        memory[54451] <=  8'h61;        memory[54452] <=  8'h63;        memory[54453] <=  8'h72;        memory[54454] <=  8'h6e;        memory[54455] <=  8'h74;        memory[54456] <=  8'h61;        memory[54457] <=  8'h62;        memory[54458] <=  8'h74;        memory[54459] <=  8'h6e;        memory[54460] <=  8'h61;        memory[54461] <=  8'h72;        memory[54462] <=  8'h62;        memory[54463] <=  8'h78;        memory[54464] <=  8'h74;        memory[54465] <=  8'h61;        memory[54466] <=  8'h72;        memory[54467] <=  8'h62;        memory[54468] <=  8'h61;        memory[54469] <=  8'h72;        memory[54470] <=  8'h74;        memory[54471] <=  8'h74;        memory[54472] <=  8'h62;        memory[54473] <=  8'h61;        memory[54474] <=  8'h72;        memory[54475] <=  8'h74;        memory[54476] <=  8'h78;        memory[54477] <=  8'h61;        memory[54478] <=  8'h74;        memory[54479] <=  8'h6b;        memory[54480] <=  8'h73;        memory[54481] <=  8'h68;        memory[54482] <=  8'h63;        memory[54483] <=  8'h66;        memory[54484] <=  8'h69;        memory[54485] <=  8'h77;        memory[54486] <=  8'h68;        memory[54487] <=  8'h61;        memory[54488] <=  8'h74;        memory[54489] <=  8'h61;        memory[54490] <=  8'h6e;        memory[54491] <=  8'h61;        memory[54492] <=  8'h62;        memory[54493] <=  8'h61;        memory[54494] <=  8'h63;        memory[54495] <=  8'h61;        memory[54496] <=  8'h74;        memory[54497] <=  8'h61;        memory[54498] <=  8'h62;        memory[54499] <=  8'h61;        memory[54500] <=  8'h72;        memory[54501] <=  8'h63;        memory[54502] <=  8'h61;        memory[54503] <=  8'h68;        memory[54504] <=  8'h64;        memory[54505] <=  8'h75;        memory[54506] <=  8'h63;        memory[54507] <=  8'h74;        memory[54508] <=  8'h61;        memory[54509] <=  8'h64;        memory[54510] <=  8'h61;        memory[54511] <=  8'h61;        memory[54512] <=  8'h63;        memory[54513] <=  8'h61;        memory[54514] <=  8'h72;        memory[54515] <=  8'h63;        memory[54516] <=  8'h74;        memory[54517] <=  8'h72;        memory[54518] <=  8'h63;        memory[54519] <=  8'h61;        memory[54520] <=  8'h74;        memory[54521] <=  8'h72;        memory[54522] <=  8'h63;        memory[54523] <=  8'h61;        memory[54524] <=  8'h74;        memory[54525] <=  8'h63;        memory[54526] <=  8'h62;        memory[54527] <=  8'h61;        memory[54528] <=  8'h74;        memory[54529] <=  8'h62;        memory[54530] <=  8'h72;        memory[54531] <=  8'h63;        memory[54532] <=  8'h61;        memory[54533] <=  8'h74;        memory[54534] <=  8'h72;        memory[54535] <=  8'h6e;        memory[54536] <=  8'h62;        memory[54537] <=  8'h61;        memory[54538] <=  8'h63;        memory[54539] <=  8'h61;        memory[54540] <=  8'h74;        memory[54541] <=  8'h79;        memory[54542] <=  8'h73;        memory[54543] <=  8'h6e;        memory[54544] <=  8'h63;        memory[54545] <=  8'h74;        memory[54546] <=  8'h61;        memory[54547] <=  8'h6e;        memory[54548] <=  8'h62;        memory[54549] <=  8'h61;        memory[54550] <=  8'h63;        memory[54551] <=  8'h72;        memory[54552] <=  8'h6e;        memory[54553] <=  8'h74;        memory[54554] <=  8'h61;        memory[54555] <=  8'h62;        memory[54556] <=  8'h74;        memory[54557] <=  8'h6e;        memory[54558] <=  8'h61;        memory[54559] <=  8'h72;        memory[54560] <=  8'h62;        memory[54561] <=  8'h78;        memory[54562] <=  8'h74;        memory[54563] <=  8'h61;        memory[54564] <=  8'h72;        memory[54565] <=  8'h64;        memory[54566] <=  8'h66;        memory[54567] <=  8'h73;        memory[54568] <=  8'h67;        memory[54569] <=  8'h76;        memory[54570] <=  8'h68;        memory[54571] <=  8'h62;        memory[54572] <=  8'h6b;        memory[54573] <=  8'h6a;        memory[54574] <=  8'h6e;        memory[54575] <=  8'h6d;        memory[54576] <=  8'h62;        memory[54577] <=  8'h76;        memory[54578] <=  8'h78;        memory[54579] <=  8'h63;        memory[54580] <=  8'h73;        memory[54581] <=  8'h66;        memory[54582] <=  8'h72;        memory[54583] <=  8'h74;        memory[54584] <=  8'h79;        memory[54585] <=  8'h75;        memory[54586] <=  8'h6a;        memory[54587] <=  8'h6e;        memory[54588] <=  8'h62;        memory[54589] <=  8'h76;        memory[54590] <=  8'h63;        memory[54591] <=  8'h64;        memory[54592] <=  8'h74;        memory[54593] <=  8'h79;        memory[54594] <=  8'h75;        memory[54595] <=  8'h69;        memory[54596] <=  8'h6b;        memory[54597] <=  8'h6d;        memory[54598] <=  8'h6e;        memory[54599] <=  8'h62;        memory[54600] <=  8'h76;        memory[54601] <=  8'h63;        memory[54602] <=  8'h78;        memory[54603] <=  8'h73;        memory[54604] <=  8'h64;        memory[54605] <=  8'h72;        memory[54606] <=  8'h74;        memory[54607] <=  8'h79;        memory[54608] <=  8'h75;        memory[54609] <=  8'h69;        memory[54610] <=  8'h6b;        memory[54611] <=  8'h6d;        memory[54612] <=  8'h6e;        memory[54613] <=  8'h62;        memory[54614] <=  8'h76;        memory[54615] <=  8'h63;        memory[54616] <=  8'h73;        memory[54617] <=  8'h77;        memory[54618] <=  8'h33;        memory[54619] <=  8'h34;        memory[54620] <=  8'h35;        memory[54621] <=  8'h36;        memory[54622] <=  8'h37;        memory[54623] <=  8'h38;        memory[54624] <=  8'h69;        memory[54625] <=  8'h6b;        memory[54626] <=  8'h6d;        memory[54627] <=  8'h6e;        memory[54628] <=  8'h62;        memory[54629] <=  8'h76;        memory[54630] <=  8'h63;        memory[54631] <=  8'h64;        memory[54632] <=  8'h65;        memory[54633] <=  8'h72;        memory[54634] <=  8'h36;        memory[54635] <=  8'h37;        memory[54636] <=  8'h38;        memory[54637] <=  8'h69;        memory[54638] <=  8'h6f;        memory[54639] <=  8'h6b;        memory[54640] <=  8'h6a;        memory[54641] <=  8'h6e;        memory[54642] <=  8'h62;        memory[54643] <=  8'h76;        memory[54644] <=  8'h63;        memory[54645] <=  8'h64;        memory[54646] <=  8'h72;        memory[54647] <=  8'h74;        memory[54648] <=  8'h79;        memory[54649] <=  8'h75;        memory[54650] <=  8'h73;        memory[54651] <=  8'h6a;        memory[54652] <=  8'h63;        memory[54653] <=  8'h6e;        memory[54654] <=  8'h62;        memory[54655] <=  8'h64;        memory[54656] <=  8'h66;        memory[54657] <=  8'h73;        memory[54658] <=  8'h74;        memory[54659] <=  8'h79;        memory[54660] <=  8'h75;        memory[54661] <=  8'h61;        memory[54662] <=  8'h69;        memory[54663] <=  8'h6b;        memory[54664] <=  8'h78;        memory[54665] <=  8'h6d;        memory[54666] <=  8'h6e;        memory[54667] <=  8'h73;        memory[54668] <=  8'h6a;        memory[54669] <=  8'h6f;        memory[54670] <=  8'h64;        memory[54671] <=  8'h6c;        memory[54672] <=  8'h63;        memory[54673] <=  8'h78;        memory[54674] <=  8'h62;        memory[54675] <=  8'h61;        memory[54676] <=  8'h72;        memory[54677] <=  8'h74;        memory[54678] <=  8'h78;        memory[54679] <=  8'h61;        memory[54680] <=  8'h74;        memory[54681] <=  8'h6b;        memory[54682] <=  8'h73;        memory[54683] <=  8'h68;        memory[54684] <=  8'h63;        memory[54685] <=  8'h66;        memory[54686] <=  8'h69;        memory[54687] <=  8'h77;        memory[54688] <=  8'h68;        memory[54689] <=  8'h61;        memory[54690] <=  8'h74;        memory[54691] <=  8'h61;        memory[54692] <=  8'h6e;        memory[54693] <=  8'h61;        memory[54694] <=  8'h62;        memory[54695] <=  8'h61;        memory[54696] <=  8'h63;        memory[54697] <=  8'h61;        memory[54698] <=  8'h74;        memory[54699] <=  8'h61;        memory[54700] <=  8'h62;        memory[54701] <=  8'h61;        memory[54702] <=  8'h72;        memory[54703] <=  8'h63;        memory[54704] <=  8'h61;        memory[54705] <=  8'h68;        memory[54706] <=  8'h64;        memory[54707] <=  8'h75;        memory[54708] <=  8'h63;        memory[54709] <=  8'h74;        memory[54710] <=  8'h61;        memory[54711] <=  8'h64;        memory[54712] <=  8'h61;        memory[54713] <=  8'h61;        memory[54714] <=  8'h63;        memory[54715] <=  8'h61;        memory[54716] <=  8'h72;        memory[54717] <=  8'h62;        memory[54718] <=  8'h61;        memory[54719] <=  8'h72;        memory[54720] <=  8'h74;        memory[54721] <=  8'h78;        memory[54722] <=  8'h61;        memory[54723] <=  8'h74;        memory[54724] <=  8'h6b;        memory[54725] <=  8'h73;        memory[54726] <=  8'h68;        memory[54727] <=  8'h63;        memory[54728] <=  8'h66;        memory[54729] <=  8'h69;        memory[54730] <=  8'h77;        memory[54731] <=  8'h68;        memory[54732] <=  8'h61;        memory[54733] <=  8'h74;        memory[54734] <=  8'h61;        memory[54735] <=  8'h6e;        memory[54736] <=  8'h61;        memory[54737] <=  8'h62;        memory[54738] <=  8'h61;        memory[54739] <=  8'h63;        memory[54740] <=  8'h61;        memory[54741] <=  8'h74;        memory[54742] <=  8'h61;        memory[54743] <=  8'h62;        memory[54744] <=  8'h61;        memory[54745] <=  8'h72;        memory[54746] <=  8'h63;        memory[54747] <=  8'h61;        memory[54748] <=  8'h68;        memory[54749] <=  8'h64;        memory[54750] <=  8'h75;        memory[54751] <=  8'h63;        memory[54752] <=  8'h74;        memory[54753] <=  8'h61;        memory[54754] <=  8'h64;        memory[54755] <=  8'h61;        memory[54756] <=  8'h61;        memory[54757] <=  8'h63;        memory[54758] <=  8'h61;        memory[54759] <=  8'h72;        memory[54760] <=  8'h62;        memory[54761] <=  8'h61;        memory[54762] <=  8'h72;        memory[54763] <=  8'h74;        memory[54764] <=  8'h78;        memory[54765] <=  8'h61;        memory[54766] <=  8'h74;        memory[54767] <=  8'h6b;        memory[54768] <=  8'h73;        memory[54769] <=  8'h68;        memory[54770] <=  8'h63;        memory[54771] <=  8'h66;        memory[54772] <=  8'h69;        memory[54773] <=  8'h77;        memory[54774] <=  8'h68;        memory[54775] <=  8'h61;        memory[54776] <=  8'h74;        memory[54777] <=  8'h61;        memory[54778] <=  8'h6e;        memory[54779] <=  8'h61;        memory[54780] <=  8'h62;        memory[54781] <=  8'h61;        memory[54782] <=  8'h63;        memory[54783] <=  8'h61;        memory[54784] <=  8'h74;        memory[54785] <=  8'h61;        memory[54786] <=  8'h62;        memory[54787] <=  8'h61;        memory[54788] <=  8'h72;        memory[54789] <=  8'h63;        memory[54790] <=  8'h61;        memory[54791] <=  8'h68;        memory[54792] <=  8'h64;        memory[54793] <=  8'h75;        memory[54794] <=  8'h63;        memory[54795] <=  8'h74;        memory[54796] <=  8'h61;        memory[54797] <=  8'h64;        memory[54798] <=  8'h61;        memory[54799] <=  8'h61;        memory[54800] <=  8'h63;        memory[54801] <=  8'h61;        memory[54802] <=  8'h72;        memory[54803] <=  8'h62;        memory[54804] <=  8'h61;        memory[54805] <=  8'h72;        memory[54806] <=  8'h74;        memory[54807] <=  8'h78;        memory[54808] <=  8'h61;        memory[54809] <=  8'h74;        memory[54810] <=  8'h6b;        memory[54811] <=  8'h73;        memory[54812] <=  8'h68;        memory[54813] <=  8'h63;        memory[54814] <=  8'h66;        memory[54815] <=  8'h69;        memory[54816] <=  8'h77;        memory[54817] <=  8'h68;        memory[54818] <=  8'h61;        memory[54819] <=  8'h74;        memory[54820] <=  8'h61;        memory[54821] <=  8'h6e;        memory[54822] <=  8'h61;        memory[54823] <=  8'h62;        memory[54824] <=  8'h61;        memory[54825] <=  8'h63;        memory[54826] <=  8'h61;        memory[54827] <=  8'h74;        memory[54828] <=  8'h61;        memory[54829] <=  8'h62;        memory[54830] <=  8'h61;        memory[54831] <=  8'h72;        memory[54832] <=  8'h63;        memory[54833] <=  8'h61;        memory[54834] <=  8'h68;        memory[54835] <=  8'h64;        memory[54836] <=  8'h75;        memory[54837] <=  8'h63;        memory[54838] <=  8'h74;        memory[54839] <=  8'h61;        memory[54840] <=  8'h64;        memory[54841] <=  8'h61;        memory[54842] <=  8'h61;        memory[54843] <=  8'h63;        memory[54844] <=  8'h61;        memory[54845] <=  8'h72;        memory[54846] <=  8'h62;        memory[54847] <=  8'h61;        memory[54848] <=  8'h72;        memory[54849] <=  8'h74;        memory[54850] <=  8'h78;        memory[54851] <=  8'h61;        memory[54852] <=  8'h74;        memory[54853] <=  8'h6b;        memory[54854] <=  8'h73;        memory[54855] <=  8'h68;        memory[54856] <=  8'h63;        memory[54857] <=  8'h66;        memory[54858] <=  8'h69;        memory[54859] <=  8'h77;        memory[54860] <=  8'h68;        memory[54861] <=  8'h61;        memory[54862] <=  8'h74;        memory[54863] <=  8'h61;        memory[54864] <=  8'h6e;        memory[54865] <=  8'h61;        memory[54866] <=  8'h62;        memory[54867] <=  8'h61;        memory[54868] <=  8'h63;        memory[54869] <=  8'h61;        memory[54870] <=  8'h74;        memory[54871] <=  8'h61;        memory[54872] <=  8'h62;        memory[54873] <=  8'h61;        memory[54874] <=  8'h72;        memory[54875] <=  8'h63;        memory[54876] <=  8'h61;        memory[54877] <=  8'h68;        memory[54878] <=  8'h64;        memory[54879] <=  8'h75;        memory[54880] <=  8'h63;        memory[54881] <=  8'h74;        memory[54882] <=  8'h61;        memory[54883] <=  8'h64;        memory[54884] <=  8'h61;        memory[54885] <=  8'h61;        memory[54886] <=  8'h63;        memory[54887] <=  8'h61;        memory[54888] <=  8'h72;        memory[54889] <=  8'h62;        memory[54890] <=  8'h61;        memory[54891] <=  8'h72;        memory[54892] <=  8'h74;        memory[54893] <=  8'h78;        memory[54894] <=  8'h61;        memory[54895] <=  8'h74;        memory[54896] <=  8'h6b;        memory[54897] <=  8'h73;        memory[54898] <=  8'h68;        memory[54899] <=  8'h63;        memory[54900] <=  8'h66;        memory[54901] <=  8'h69;        memory[54902] <=  8'h77;        memory[54903] <=  8'h68;        memory[54904] <=  8'h61;        memory[54905] <=  8'h74;        memory[54906] <=  8'h61;        memory[54907] <=  8'h6e;        memory[54908] <=  8'h61;        memory[54909] <=  8'h62;        memory[54910] <=  8'h61;        memory[54911] <=  8'h63;        memory[54912] <=  8'h61;        memory[54913] <=  8'h74;        memory[54914] <=  8'h61;        memory[54915] <=  8'h62;        memory[54916] <=  8'h61;        memory[54917] <=  8'h72;        memory[54918] <=  8'h63;        memory[54919] <=  8'h61;        memory[54920] <=  8'h68;        memory[54921] <=  8'h64;        memory[54922] <=  8'h75;        memory[54923] <=  8'h63;        memory[54924] <=  8'h74;        memory[54925] <=  8'h61;        memory[54926] <=  8'h64;        memory[54927] <=  8'h61;        memory[54928] <=  8'h61;        memory[54929] <=  8'h63;        memory[54930] <=  8'h61;        memory[54931] <=  8'h72;        memory[54932] <=  8'h62;        memory[54933] <=  8'h61;        memory[54934] <=  8'h72;        memory[54935] <=  8'h74;        memory[54936] <=  8'h78;        memory[54937] <=  8'h61;        memory[54938] <=  8'h74;        memory[54939] <=  8'h6b;        memory[54940] <=  8'h73;        memory[54941] <=  8'h68;        memory[54942] <=  8'h63;        memory[54943] <=  8'h66;        memory[54944] <=  8'h69;        memory[54945] <=  8'h77;        memory[54946] <=  8'h68;        memory[54947] <=  8'h61;        memory[54948] <=  8'h74;        memory[54949] <=  8'h61;        memory[54950] <=  8'h6e;        memory[54951] <=  8'h61;        memory[54952] <=  8'h62;        memory[54953] <=  8'h61;        memory[54954] <=  8'h63;        memory[54955] <=  8'h61;        memory[54956] <=  8'h74;        memory[54957] <=  8'h61;        memory[54958] <=  8'h62;        memory[54959] <=  8'h61;        memory[54960] <=  8'h72;        memory[54961] <=  8'h63;        memory[54962] <=  8'h61;        memory[54963] <=  8'h68;        memory[54964] <=  8'h64;        memory[54965] <=  8'h75;        memory[54966] <=  8'h63;        memory[54967] <=  8'h74;        memory[54968] <=  8'h61;        memory[54969] <=  8'h64;        memory[54970] <=  8'h61;        memory[54971] <=  8'h61;        memory[54972] <=  8'h63;        memory[54973] <=  8'h61;        memory[54974] <=  8'h72;        memory[54975] <=  8'h62;        memory[54976] <=  8'h61;        memory[54977] <=  8'h72;        memory[54978] <=  8'h74;        memory[54979] <=  8'h78;        memory[54980] <=  8'h61;        memory[54981] <=  8'h74;        memory[54982] <=  8'h6b;        memory[54983] <=  8'h73;        memory[54984] <=  8'h68;        memory[54985] <=  8'h63;        memory[54986] <=  8'h66;        memory[54987] <=  8'h69;        memory[54988] <=  8'h77;        memory[54989] <=  8'h68;        memory[54990] <=  8'h61;        memory[54991] <=  8'h74;        memory[54992] <=  8'h61;        memory[54993] <=  8'h6e;        memory[54994] <=  8'h61;        memory[54995] <=  8'h62;        memory[54996] <=  8'h61;        memory[54997] <=  8'h63;        memory[54998] <=  8'h61;        memory[54999] <=  8'h74;        memory[55000] <=  8'h61;        memory[55001] <=  8'h62;        memory[55002] <=  8'h61;        memory[55003] <=  8'h72;        memory[55004] <=  8'h63;        memory[55005] <=  8'h61;        memory[55006] <=  8'h68;        memory[55007] <=  8'h64;        memory[55008] <=  8'h75;        memory[55009] <=  8'h63;        memory[55010] <=  8'h74;        memory[55011] <=  8'h61;        memory[55012] <=  8'h64;        memory[55013] <=  8'h61;        memory[55014] <=  8'h61;        memory[55015] <=  8'h63;        memory[55016] <=  8'h61;        memory[55017] <=  8'h72;        memory[55018] <=  8'h62;        memory[55019] <=  8'h61;        memory[55020] <=  8'h72;        memory[55021] <=  8'h74;        memory[55022] <=  8'h78;        memory[55023] <=  8'h61;        memory[55024] <=  8'h74;        memory[55025] <=  8'h6b;        memory[55026] <=  8'h73;        memory[55027] <=  8'h68;        memory[55028] <=  8'h63;        memory[55029] <=  8'h66;        memory[55030] <=  8'h69;        memory[55031] <=  8'h77;        memory[55032] <=  8'h68;        memory[55033] <=  8'h61;        memory[55034] <=  8'h74;        memory[55035] <=  8'h61;        memory[55036] <=  8'h6e;        memory[55037] <=  8'h61;        memory[55038] <=  8'h62;        memory[55039] <=  8'h61;        memory[55040] <=  8'h63;        memory[55041] <=  8'h61;        memory[55042] <=  8'h74;        memory[55043] <=  8'h61;        memory[55044] <=  8'h62;        memory[55045] <=  8'h61;        memory[55046] <=  8'h72;        memory[55047] <=  8'h63;        memory[55048] <=  8'h61;        memory[55049] <=  8'h68;        memory[55050] <=  8'h64;        memory[55051] <=  8'h75;        memory[55052] <=  8'h63;        memory[55053] <=  8'h74;        memory[55054] <=  8'h61;        memory[55055] <=  8'h64;        memory[55056] <=  8'h61;        memory[55057] <=  8'h61;        memory[55058] <=  8'h63;        memory[55059] <=  8'h61;        memory[55060] <=  8'h72;        memory[55061] <=  8'h62;        memory[55062] <=  8'h61;        memory[55063] <=  8'h72;        memory[55064] <=  8'h74;        memory[55065] <=  8'h74;        memory[55066] <=  8'h62;        memory[55067] <=  8'h61;        memory[55068] <=  8'h72;        memory[55069] <=  8'h74;        memory[55070] <=  8'h78;        memory[55071] <=  8'h61;        memory[55072] <=  8'h74;        memory[55073] <=  8'h6b;        memory[55074] <=  8'h73;        memory[55075] <=  8'h68;        memory[55076] <=  8'h63;        memory[55077] <=  8'h66;        memory[55078] <=  8'h69;        memory[55079] <=  8'h77;        memory[55080] <=  8'h68;        memory[55081] <=  8'h61;        memory[55082] <=  8'h74;        memory[55083] <=  8'h61;        memory[55084] <=  8'h6e;        memory[55085] <=  8'h61;        memory[55086] <=  8'h62;        memory[55087] <=  8'h61;        memory[55088] <=  8'h63;        memory[55089] <=  8'h61;        memory[55090] <=  8'h74;        memory[55091] <=  8'h61;        memory[55092] <=  8'h62;        memory[55093] <=  8'h61;        memory[55094] <=  8'h72;        memory[55095] <=  8'h63;        memory[55096] <=  8'h61;        memory[55097] <=  8'h68;        memory[55098] <=  8'h64;        memory[55099] <=  8'h75;        memory[55100] <=  8'h63;        memory[55101] <=  8'h74;        memory[55102] <=  8'h61;        memory[55103] <=  8'h64;        memory[55104] <=  8'h61;        memory[55105] <=  8'h61;        memory[55106] <=  8'h63;        memory[55107] <=  8'h61;        memory[55108] <=  8'h72;        memory[55109] <=  8'h63;        memory[55110] <=  8'h74;        memory[55111] <=  8'h72;        memory[55112] <=  8'h63;        memory[55113] <=  8'h61;        memory[55114] <=  8'h74;        memory[55115] <=  8'h72;        memory[55116] <=  8'h63;        memory[55117] <=  8'h61;        memory[55118] <=  8'h74;        memory[55119] <=  8'h63;        memory[55120] <=  8'h62;        memory[55121] <=  8'h61;        memory[55122] <=  8'h74;        memory[55123] <=  8'h62;        memory[55124] <=  8'h72;        memory[55125] <=  8'h63;        memory[55126] <=  8'h61;        memory[55127] <=  8'h72;        memory[55128] <=  8'h62;        memory[55129] <=  8'h78;        memory[55130] <=  8'h74;        memory[55131] <=  8'h61;        memory[55132] <=  8'h72;        memory[55133] <=  8'h64;        memory[55134] <=  8'h66;        memory[55135] <=  8'h73;        memory[55136] <=  8'h67;        memory[55137] <=  8'h76;        memory[55138] <=  8'h68;        memory[55139] <=  8'h62;        memory[55140] <=  8'h6b;        memory[55141] <=  8'h6a;        memory[55142] <=  8'h6e;        memory[55143] <=  8'h6d;        memory[55144] <=  8'h62;        memory[55145] <=  8'h76;        memory[55146] <=  8'h78;        memory[55147] <=  8'h63;        memory[55148] <=  8'h73;        memory[55149] <=  8'h66;        memory[55150] <=  8'h72;        memory[55151] <=  8'h74;        memory[55152] <=  8'h79;        memory[55153] <=  8'h75;        memory[55154] <=  8'h6a;        memory[55155] <=  8'h6e;        memory[55156] <=  8'h62;        memory[55157] <=  8'h76;        memory[55158] <=  8'h63;        memory[55159] <=  8'h64;        memory[55160] <=  8'h74;        memory[55161] <=  8'h79;        memory[55162] <=  8'h75;        memory[55163] <=  8'h69;        memory[55164] <=  8'h6b;        memory[55165] <=  8'h6d;        memory[55166] <=  8'h6e;        memory[55167] <=  8'h62;        memory[55168] <=  8'h76;        memory[55169] <=  8'h63;        memory[55170] <=  8'h78;        memory[55171] <=  8'h73;        memory[55172] <=  8'h64;        memory[55173] <=  8'h72;        memory[55174] <=  8'h74;        memory[55175] <=  8'h79;        memory[55176] <=  8'h75;        memory[55177] <=  8'h69;        memory[55178] <=  8'h6b;        memory[55179] <=  8'h6d;        memory[55180] <=  8'h6e;        memory[55181] <=  8'h62;        memory[55182] <=  8'h76;        memory[55183] <=  8'h63;        memory[55184] <=  8'h73;        memory[55185] <=  8'h77;        memory[55186] <=  8'h33;        memory[55187] <=  8'h34;        memory[55188] <=  8'h35;        memory[55189] <=  8'h36;        memory[55190] <=  8'h37;        memory[55191] <=  8'h38;        memory[55192] <=  8'h69;        memory[55193] <=  8'h6b;        memory[55194] <=  8'h6d;        memory[55195] <=  8'h6e;        memory[55196] <=  8'h62;        memory[55197] <=  8'h76;        memory[55198] <=  8'h63;        memory[55199] <=  8'h64;        memory[55200] <=  8'h65;        memory[55201] <=  8'h72;        memory[55202] <=  8'h36;        memory[55203] <=  8'h37;        memory[55204] <=  8'h38;        memory[55205] <=  8'h69;        memory[55206] <=  8'h6f;        memory[55207] <=  8'h6b;        memory[55208] <=  8'h6a;        memory[55209] <=  8'h6e;        memory[55210] <=  8'h62;        memory[55211] <=  8'h76;        memory[55212] <=  8'h63;        memory[55213] <=  8'h64;        memory[55214] <=  8'h72;        memory[55215] <=  8'h74;        memory[55216] <=  8'h79;        memory[55217] <=  8'h75;        memory[55218] <=  8'h73;        memory[55219] <=  8'h6a;        memory[55220] <=  8'h63;        memory[55221] <=  8'h6e;        memory[55222] <=  8'h62;        memory[55223] <=  8'h64;        memory[55224] <=  8'h66;        memory[55225] <=  8'h73;        memory[55226] <=  8'h74;        memory[55227] <=  8'h79;        memory[55228] <=  8'h75;        memory[55229] <=  8'h61;        memory[55230] <=  8'h69;        memory[55231] <=  8'h6b;        memory[55232] <=  8'h78;        memory[55233] <=  8'h6d;        memory[55234] <=  8'h6e;        memory[55235] <=  8'h73;        memory[55236] <=  8'h6a;        memory[55237] <=  8'h6f;        memory[55238] <=  8'h64;        memory[55239] <=  8'h6c;        memory[55240] <=  8'h63;        memory[55241] <=  8'h78;        memory[55242] <=  8'h2c;        memory[55243] <=  8'h6d;        memory[55244] <=  8'h73;        memory[55245] <=  8'h6b;        memory[55246] <=  8'h64;        memory[55247] <=  8'h6c;        memory[55248] <=  8'h70;        memory[55249] <=  8'h5b;        memory[55250] <=  8'h3b;        memory[55251] <=  8'h73;        memory[55252] <=  8'h6c;        memory[55253] <=  8'h64;        memory[55254] <=  8'h70;        memory[55255] <=  8'h76;        memory[55256] <=  8'h63;        memory[55257] <=  8'h5b;        memory[55258] <=  8'h78;        memory[55259] <=  8'h76;        memory[55260] <=  8'h63;        memory[55261] <=  8'h5b;        memory[55262] <=  8'h78;        memory[55263] <=  8'h70;        memory[55264] <=  8'h6f;        memory[55265] <=  8'h20;        memory[55266] <=  8'h62;        memory[55267] <=  8'h61;        memory[55268] <=  8'h72;        memory[55269] <=  8'h74;        memory[55270] <=  8'h74;        memory[55271] <=  8'h62;        memory[55272] <=  8'h61;        memory[55273] <=  8'h72;        memory[55274] <=  8'h74;        memory[55275] <=  8'h78;        memory[55276] <=  8'h61;        memory[55277] <=  8'h74;        memory[55278] <=  8'h6b;        memory[55279] <=  8'h73;        memory[55280] <=  8'h68;        memory[55281] <=  8'h63;        memory[55282] <=  8'h66;        memory[55283] <=  8'h69;        memory[55284] <=  8'h77;        memory[55285] <=  8'h68;        memory[55286] <=  8'h61;        memory[55287] <=  8'h69;        memory[55288] <=  8'h6a;        memory[55289] <=  8'h78;        memory[55290] <=  8'h5d;        memory[55291] <=  8'h65;        memory[55292] <=  8'h6b;        memory[55293] <=  8'h6f;        memory[55294] <=  8'h39;        memory[55295] <=  8'h64;        memory[55296] <=  8'h75;        memory[55297] <=  8'h38;        memory[55298] <=  8'h79;        memory[55299] <=  8'h20;        memory[55300] <=  8'h37;        memory[55301] <=  8'h63;        memory[55302] <=  8'h67;        memory[55303] <=  8'h78;        memory[55304] <=  8'h63;        memory[55305] <=  8'h75;        memory[55306] <=  8'h68;        memory[55307] <=  8'h69;        memory[55308] <=  8'h6a;        memory[55309] <=  8'h77;        memory[55310] <=  8'h69;        memory[55311] <=  8'h64;        memory[55312] <=  8'h66;        memory[55313] <=  8'h68;        memory[55314] <=  8'h75;        memory[55315] <=  8'h76;        memory[55316] <=  8'h64;        memory[55317] <=  8'h62;        memory[55318] <=  8'h66;        memory[55319] <=  8'h6a;        memory[55320] <=  8'h6e;        memory[55321] <=  8'h6b;        memory[55322] <=  8'h6a;        memory[55323] <=  8'h65;        memory[55324] <=  8'h38;        memory[55325] <=  8'h66;        memory[55326] <=  8'h37;        memory[55327] <=  8'h67;        memory[55328] <=  8'h79;        memory[55329] <=  8'h76;        memory[55330] <=  8'h63;        memory[55331] <=  8'h68;        memory[55332] <=  8'h69;        memory[55333] <=  8'h6a;        memory[55334] <=  8'h33;        memory[55335] <=  8'h65;        memory[55336] <=  8'h67;        memory[55337] <=  8'h79;        memory[55338] <=  8'h72;        memory[55339] <=  8'h64;        memory[55340] <=  8'h62;        memory[55341] <=  8'h6e;        memory[55342] <=  8'h63;        memory[55343] <=  8'h7a;        memory[55344] <=  8'h6a;        memory[55345] <=  8'h6f;        memory[55346] <=  8'h66;        memory[55347] <=  8'h78;        memory[55348] <=  8'h6a;        memory[55349] <=  8'h69;        memory[55350] <=  8'h63;        memory[55351] <=  8'h68;        memory[55352] <=  8'h62;        memory[55353] <=  8'h6e;        memory[55354] <=  8'h6d;        memory[55355] <=  8'h63;        memory[55356] <=  8'h73;        memory[55357] <=  8'h6c;        memory[55358] <=  8'h6b;        memory[55359] <=  8'h6a;        memory[55360] <=  8'h69;        memory[55361] <=  8'h68;        memory[55362] <=  8'h76;        memory[55363] <=  8'h75;        memory[55364] <=  8'h69;        memory[55365] <=  8'h64;        memory[55366] <=  8'h68;        memory[55367] <=  8'h75;        memory[55368] <=  8'h67;        memory[55369] <=  8'h79;        memory[55370] <=  8'h62;        memory[55371] <=  8'h68;        memory[55372] <=  8'h65;        memory[55373] <=  8'h6a;        memory[55374] <=  8'h72;        memory[55375] <=  8'h6b;        memory[55376] <=  8'h6a;        memory[55377] <=  8'h6f;        memory[55378] <=  8'h64;        memory[55379] <=  8'h67;        memory[55380] <=  8'h69;        memory[55381] <=  8'h75;        memory[55382] <=  8'h69;        memory[55383] <=  8'h67;        memory[55384] <=  8'h76;        memory[55385] <=  8'h79;        memory[55386] <=  8'h75;        memory[55387] <=  8'h67;        memory[55388] <=  8'h78;        memory[55389] <=  8'h68;        memory[55390] <=  8'h63;        memory[55391] <=  8'h20;        memory[55392] <=  8'h20;        memory[55393] <=  8'h20;        memory[55394] <=  8'h78;        memory[55395] <=  8'h76;        memory[55396] <=  8'h20;        memory[55397] <=  8'h63;        memory[55398] <=  8'h78;        memory[55399] <=  8'h67;        memory[55400] <=  8'h79;        memory[55401] <=  8'h63;        memory[55402] <=  8'h75;        memory[55403] <=  8'h68;        memory[55404] <=  8'h6a;        memory[55405] <=  8'h6b;        memory[55406] <=  8'h61;        memory[55407] <=  8'h6c;        memory[55408] <=  8'h78;        memory[55409] <=  8'h76;        memory[55410] <=  8'h70;        memory[55411] <=  8'h6f;        memory[55412] <=  8'h69;        memory[55413] <=  8'h6a;        memory[55414] <=  8'h69;        memory[55415] <=  8'h68;        memory[55416] <=  8'h6a;        memory[55417] <=  8'h62;        memory[55418] <=  8'h77;        memory[55419] <=  8'h65;        memory[55420] <=  8'h6e;        memory[55421] <=  8'h61;        memory[55422] <=  8'h66;        memory[55423] <=  8'h6d;        memory[55424] <=  8'h64;        memory[55425] <=  8'h6b;        memory[55426] <=  8'h6d;        memory[55427] <=  8'h76;        memory[55428] <=  8'h6c;        memory[55429] <=  8'h63;        memory[55430] <=  8'h6f;        memory[55431] <=  8'h64;        memory[55432] <=  8'h69;        memory[55433] <=  8'h75;        memory[55434] <=  8'h68;        memory[55435] <=  8'h73;        memory[55436] <=  8'h66;        memory[55437] <=  8'h65;        memory[55438] <=  8'h62;        memory[55439] <=  8'h6e;        memory[55440] <=  8'h64;        memory[55441] <=  8'h73;        memory[55442] <=  8'h63;        memory[55443] <=  8'h6b;        memory[55444] <=  8'h20;        memory[55445] <=  8'h78;        memory[55446] <=  8'h6a;        memory[55447] <=  8'h78;        memory[55448] <=  8'h63;        memory[55449] <=  8'h73;        memory[55450] <=  8'h64;        memory[55451] <=  8'h66;        memory[55452] <=  8'h6b;        memory[55453] <=  8'h64;        memory[55454] <=  8'h6e;        memory[55455] <=  8'h6d;        memory[55456] <=  8'h64;        memory[55457] <=  8'h73;        memory[55458] <=  8'h63;        memory[55459] <=  8'h6b;        memory[55460] <=  8'h78;        memory[55461] <=  8'h6c;        memory[55462] <=  8'h6f;        memory[55463] <=  8'h66;        memory[55464] <=  8'h6a;        memory[55465] <=  8'h69;        memory[55466] <=  8'h61;        memory[55467] <=  8'h62;        memory[55468] <=  8'h6e;        memory[55469] <=  8'h20;        memory[55470] <=  8'h78;        memory[55471] <=  8'h6b;        memory[55472] <=  8'h6d;        memory[55473] <=  8'h20;        memory[55474] <=  8'h6f;        memory[55475] <=  8'h63;        memory[55476] <=  8'h76;        memory[55477] <=  8'h73;        memory[55478] <=  8'h64;        memory[55479] <=  8'h69;        memory[55480] <=  8'h66;        memory[55481] <=  8'h68;        memory[55482] <=  8'h65;        memory[55483] <=  8'h71;        memory[55484] <=  8'h6a;        memory[55485] <=  8'h77;        memory[55486] <=  8'h62;        memory[55487] <=  8'h65;        memory[55488] <=  8'h6e;        memory[55489] <=  8'h20;        memory[55490] <=  8'h6d;        memory[55491] <=  8'h64;        memory[55492] <=  8'h73;        memory[55493] <=  8'h6c;        memory[55494] <=  8'h76;        memory[55495] <=  8'h6b;        memory[55496] <=  8'h63;        memory[55497] <=  8'h78;        memory[55498] <=  8'h20;        memory[55499] <=  8'h6f;        memory[55500] <=  8'h78;        memory[55501] <=  8'h69;        memory[55502] <=  8'h63;        memory[55503] <=  8'h6a;        memory[55504] <=  8'h76;        memory[55505] <=  8'h64;        memory[55506] <=  8'h66;        memory[55507] <=  8'h65;        memory[55508] <=  8'h71;        memory[55509] <=  8'h6e;        memory[55510] <=  8'h20;        memory[55511] <=  8'h64;        memory[55512] <=  8'h6d;        memory[55513] <=  8'h73;        memory[55514] <=  8'h6c;        memory[55515] <=  8'h63;        memory[55516] <=  8'h78;        memory[55517] <=  8'h6b;        memory[55518] <=  8'h20;        memory[55519] <=  8'h6f;        memory[55520] <=  8'h78;        memory[55521] <=  8'h63;        memory[55522] <=  8'h76;        memory[55523] <=  8'h6a;        memory[55524] <=  8'h64;        memory[55525] <=  8'h62;        memory[55526] <=  8'h71;        memory[55527] <=  8'h77;        memory[55528] <=  8'h65;        memory[55529] <=  8'h6e;        memory[55530] <=  8'h6d;        memory[55531] <=  8'h64;        memory[55532] <=  8'h6c;        memory[55533] <=  8'h73;        memory[55534] <=  8'h2c;        memory[55535] <=  8'h76;        memory[55536] <=  8'h63;        memory[55537] <=  8'h78;        memory[55538] <=  8'h20;        memory[55539] <=  8'h63;        memory[55540] <=  8'h6f;        memory[55541] <=  8'h69;        memory[55542] <=  8'h76;        memory[55543] <=  8'h68;        memory[55544] <=  8'h73;        memory[55545] <=  8'h64;        memory[55546] <=  8'h62;        memory[55547] <=  8'h71;        memory[55548] <=  8'h77;        memory[55549] <=  8'h65;        memory[55550] <=  8'h6e;        memory[55551] <=  8'h64;        memory[55552] <=  8'h6b;        memory[55553] <=  8'h73;        memory[55554] <=  8'h76;        memory[55555] <=  8'h6f;        memory[55556] <=  8'h63;        memory[55557] <=  8'h20;        memory[55558] <=  8'h76;        memory[55559] <=  8'h69;        memory[55560] <=  8'h75;        memory[55561] <=  8'h69;        memory[55562] <=  8'h68;        memory[55563] <=  8'h63;        memory[55564] <=  8'h78;        memory[55565] <=  8'h69;        memory[55566] <=  8'h6f;        memory[55567] <=  8'h76;        memory[55568] <=  8'h73;        memory[55569] <=  8'h64;        memory[55570] <=  8'h61;        memory[55571] <=  8'h64;        memory[55572] <=  8'h6e;        memory[55573] <=  8'h77;        memory[55574] <=  8'h71;        memory[55575] <=  8'h6b;        memory[55576] <=  8'h6c;        memory[55577] <=  8'h73;        memory[55578] <=  8'h76;        memory[55579] <=  8'h6e;        memory[55580] <=  8'h62;        memory[55581] <=  8'h20;        memory[55582] <=  8'h64;        memory[55583] <=  8'h66;        memory[55584] <=  8'h6a;        memory[55585] <=  8'h6b;        memory[55586] <=  8'h71;        memory[55587] <=  8'h64;        memory[55588] <=  8'h77;        memory[55589] <=  8'h65;        memory[55590] <=  8'h6e;        memory[55591] <=  8'h62;        memory[55592] <=  8'h20;        memory[55593] <=  8'h64;        memory[55594] <=  8'h73;        memory[55595] <=  8'h76;        memory[55596] <=  8'h68;        memory[55597] <=  8'h64;        memory[55598] <=  8'h61;        memory[55599] <=  8'h71;        memory[55600] <=  8'h77;        memory[55601] <=  8'h6a;        memory[55602] <=  8'h65;        memory[55603] <=  8'h6e;        memory[55604] <=  8'h64;        memory[55605] <=  8'h20;        memory[55606] <=  8'h61;        memory[55607] <=  8'h63;        memory[55608] <=  8'h62;        memory[55609] <=  8'h68;        memory[55610] <=  8'h64;        memory[55611] <=  8'h61;        memory[55612] <=  8'h77;        memory[55613] <=  8'h71;        memory[55614] <=  8'h6e;        memory[55615] <=  8'h20;        memory[55616] <=  8'h62;        memory[55617] <=  8'h73;        memory[55618] <=  8'h76;        memory[55619] <=  8'h61;        memory[55620] <=  8'h67;        memory[55621] <=  8'h76;        memory[55622] <=  8'h68;        memory[55623] <=  8'h67;        memory[55624] <=  8'h61;        memory[55625] <=  8'h73;        memory[55626] <=  8'h6a;        memory[55627] <=  8'h6b;        memory[55628] <=  8'h63;        memory[55629] <=  8'h78;        memory[55630] <=  8'h76;        memory[55631] <=  8'h6e;        memory[55632] <=  8'h73;        memory[55633] <=  8'h64;        memory[55634] <=  8'h20;        memory[55635] <=  8'h66;        memory[55636] <=  8'h62;        memory[55637] <=  8'h64;        memory[55638] <=  8'h61;        memory[55639] <=  8'h73;        memory[55640] <=  8'h76;        memory[55641] <=  8'h67;        memory[55642] <=  8'h63;        memory[55643] <=  8'h79;        memory[55644] <=  8'h7a;        memory[55645] <=  8'h78;        memory[55646] <=  8'h79;        memory[55647] <=  8'h75;        memory[55648] <=  8'h20;        memory[55649] <=  8'h69;        memory[55650] <=  8'h6a;        memory[55651] <=  8'h64;        memory[55652] <=  8'h66;        memory[55653] <=  8'h6b;        memory[55654] <=  8'h61;        memory[55655] <=  8'h64;        memory[55656] <=  8'h63;        memory[55657] <=  8'h78;        memory[55658] <=  8'h68;        memory[55659] <=  8'h20;        memory[55660] <=  8'h67;        memory[55661] <=  8'h61;        memory[55662] <=  8'h68;        memory[55663] <=  8'h75;        memory[55664] <=  8'h64;        memory[55665] <=  8'h73;        memory[55666] <=  8'h69;        memory[55667] <=  8'h6a;        memory[55668] <=  8'h61;        memory[55669] <=  8'h6b;        memory[55670] <=  8'h63;        memory[55671] <=  8'h62;        memory[55672] <=  8'h61;        memory[55673] <=  8'h72;        memory[55674] <=  8'h73;        memory[55675] <=  8'h68;        memory[55676] <=  8'h64;        memory[55677] <=  8'h66;        memory[55678] <=  8'h67;        memory[55679] <=  8'h73;        memory[55680] <=  8'h68;        memory[55681] <=  8'h64;        memory[55682] <=  8'h66;        memory[55683] <=  8'h68;        memory[55684] <=  8'h64;        memory[55685] <=  8'h6a;        memory[55686] <=  8'h68;        memory[55687] <=  8'h62;        memory[55688] <=  8'h67;        memory[55689] <=  8'h63;        memory[55690] <=  8'h61;        memory[55691] <=  8'h66;        memory[55692] <=  8'h73;        memory[55693] <=  8'h79;        memory[55694] <=  8'h67;        memory[55695] <=  8'h6b;        memory[55696] <=  8'h75;        memory[55697] <=  8'h64;        memory[55698] <=  8'h68;        memory[55699] <=  8'h62;        memory[55700] <=  8'h77;        memory[55701] <=  8'h76;        memory[55702] <=  8'h67;        memory[55703] <=  8'h61;        memory[55704] <=  8'h66;        memory[55705] <=  8'h64;        memory[55706] <=  8'h74;        memory[55707] <=  8'h75;        memory[55708] <=  8'h66;        memory[55709] <=  8'h79;        memory[55710] <=  8'h67;        memory[55711] <=  8'h69;        memory[55712] <=  8'h75;        memory[55713] <=  8'h68;        memory[55714] <=  8'h6c;        memory[55715] <=  8'h6a;        memory[55716] <=  8'h62;        memory[55717] <=  8'h6b;        memory[55718] <=  8'h68;        memory[55719] <=  8'h76;        memory[55720] <=  8'h67;        memory[55721] <=  8'h63;        memory[55722] <=  8'h66;        memory[55723] <=  8'h78;        memory[55724] <=  8'h64;        memory[55725] <=  8'h74;        memory[55726] <=  8'h75;        memory[55727] <=  8'h79;        memory[55728] <=  8'h69;        memory[55729] <=  8'h75;        memory[55730] <=  8'h68;        memory[55731] <=  8'h6c;        memory[55732] <=  8'h6a;        memory[55733] <=  8'h6b;        memory[55734] <=  8'h67;        memory[55735] <=  8'h6a;        memory[55736] <=  8'h63;        memory[55737] <=  8'h66;        memory[55738] <=  8'h68;        memory[55739] <=  8'h64;        memory[55740] <=  8'h67;        memory[55741] <=  8'h72;        memory[55742] <=  8'h79;        memory[55743] <=  8'h74;        memory[55744] <=  8'h66;        memory[55745] <=  8'h75;        memory[55746] <=  8'h79;        memory[55747] <=  8'h69;        memory[55748] <=  8'h68;        memory[55749] <=  8'h6c;        memory[55750] <=  8'h62;        memory[55751] <=  8'h6d;        memory[55752] <=  8'h76;        memory[55753] <=  8'h6e;        memory[55754] <=  8'h63;        memory[55755] <=  8'h66;        memory[55756] <=  8'h68;        memory[55757] <=  8'h64;        memory[55758] <=  8'h74;        memory[55759] <=  8'h75;        memory[55760] <=  8'h67;        memory[55761] <=  8'h79;        memory[55762] <=  8'h69;        memory[55763] <=  8'h68;        memory[55764] <=  8'h75;        memory[55765] <=  8'h6a;        memory[55766] <=  8'h6c;        memory[55767] <=  8'h62;        memory[55768] <=  8'h6d;        memory[55769] <=  8'h76;        memory[55770] <=  8'h6e;        memory[55771] <=  8'h63;        memory[55772] <=  8'h66;        memory[55773] <=  8'h68;        memory[55774] <=  8'h67;        memory[55775] <=  8'h79;        memory[55776] <=  8'h68;        memory[55777] <=  8'h75;        memory[55778] <=  8'h6a;        memory[55779] <=  8'h6e;        memory[55780] <=  8'h2c;        memory[55781] <=  8'h62;        memory[55782] <=  8'h6e;        memory[55783] <=  8'h6d;        memory[55784] <=  8'h76;        memory[55785] <=  8'h6e;        memory[55786] <=  8'h63;        memory[55787] <=  8'h66;        memory[55788] <=  8'h68;        memory[55789] <=  8'h74;        memory[55790] <=  8'h79;        memory[55791] <=  8'h69;        memory[55792] <=  8'h75;        memory[55793] <=  8'h6c;        memory[55794] <=  8'h6a;        memory[55795] <=  8'h62;        memory[55796] <=  8'h6d;        memory[55797] <=  8'h76;        memory[55798] <=  8'h6e;        memory[55799] <=  8'h63;        memory[55800] <=  8'h66;        memory[55801] <=  8'h74;        memory[55802] <=  8'h75;        memory[55803] <=  8'h79;        memory[55804] <=  8'h69;        memory[55805] <=  8'h68;        memory[55806] <=  8'h6b;        memory[55807] <=  8'h62;        memory[55808] <=  8'h76;        memory[55809] <=  8'h63;        memory[55810] <=  8'h66;        memory[55811] <=  8'h67;        memory[55812] <=  8'h74;        memory[55813] <=  8'h75;        memory[55814] <=  8'h79;        memory[55815] <=  8'h69;        memory[55816] <=  8'h75;        memory[55817] <=  8'h68;        memory[55818] <=  8'h6a;        memory[55819] <=  8'h6b;        memory[55820] <=  8'h62;        memory[55821] <=  8'h76;        memory[55822] <=  8'h63;        memory[55823] <=  8'h66;        memory[55824] <=  8'h74;        memory[55825] <=  8'h75;        memory[55826] <=  8'h79;        memory[55827] <=  8'h69;        memory[55828] <=  8'h75;        memory[55829] <=  8'h6a;        memory[55830] <=  8'h6b;        memory[55831] <=  8'h6e;        memory[55832] <=  8'h62;        memory[55833] <=  8'h76;        memory[55834] <=  8'h67;        memory[55835] <=  8'h66;        memory[55836] <=  8'h74;        memory[55837] <=  8'h79;        memory[55838] <=  8'h75;        memory[55839] <=  8'h75;        memory[55840] <=  8'h69;        memory[55841] <=  8'h6a;        memory[55842] <=  8'h6b;        memory[55843] <=  8'h68;        memory[55844] <=  8'h62;        memory[55845] <=  8'h6a;        memory[55846] <=  8'h67;        memory[55847] <=  8'h68;        memory[55848] <=  8'h66;        memory[55849] <=  8'h79;        memory[55850] <=  8'h74;        memory[55851] <=  8'h79;        memory[55852] <=  8'h69;        memory[55853] <=  8'h75;        memory[55854] <=  8'h64;        memory[55855] <=  8'h6a;        memory[55856] <=  8'h6b;        memory[55857] <=  8'h68;        memory[55858] <=  8'h63;        memory[55859] <=  8'h7a;        memory[55860] <=  8'h67;        memory[55861] <=  8'h68;        memory[55862] <=  8'h74;        memory[55863] <=  8'h75;        memory[55864] <=  8'h79;        memory[55865] <=  8'h69;        memory[55866] <=  8'h61;        memory[55867] <=  8'h73;        memory[55868] <=  8'h75;        memory[55869] <=  8'h6a;        memory[55870] <=  8'h6b;        memory[55871] <=  8'h62;        memory[55872] <=  8'h6e;        memory[55873] <=  8'h61;        memory[55874] <=  8'h76;        memory[55875] <=  8'h63;        memory[55876] <=  8'h66;        memory[55877] <=  8'h68;        memory[55878] <=  8'h75;        memory[55879] <=  8'h61;        memory[55880] <=  8'h73;        memory[55881] <=  8'h79;        memory[55882] <=  8'h64;        memory[55883] <=  8'h75;        memory[55884] <=  8'h69;        memory[55885] <=  8'h6a;        memory[55886] <=  8'h61;        memory[55887] <=  8'h6b;        memory[55888] <=  8'h62;        memory[55889] <=  8'h63;        memory[55890] <=  8'h78;        memory[55891] <=  8'h68;        memory[55892] <=  8'h67;        memory[55893] <=  8'h79;        memory[55894] <=  8'h75;        memory[55895] <=  8'h7a;        memory[55896] <=  8'h63;        memory[55897] <=  8'h61;        memory[55898] <=  8'h73;        memory[55899] <=  8'h69;        memory[55900] <=  8'h75;        memory[55901] <=  8'h6f;        memory[55902] <=  8'h69;        memory[55903] <=  8'h6a;        memory[55904] <=  8'h61;        memory[55905] <=  8'h6c;        memory[55906] <=  8'h63;        memory[55907] <=  8'h78;        memory[55908] <=  8'h62;        memory[55909] <=  8'h63;        memory[55910] <=  8'h20;        memory[55911] <=  8'h6e;        memory[55912] <=  8'h76;        memory[55913] <=  8'h63;        memory[55914] <=  8'h61;        memory[55915] <=  8'h64;        memory[55916] <=  8'h73;        memory[55917] <=  8'h67;        memory[55918] <=  8'h79;        memory[55919] <=  8'h68;        memory[55920] <=  8'h75;        memory[55921] <=  8'h61;        memory[55922] <=  8'h6a;        memory[55923] <=  8'h6b;        memory[55924] <=  8'h78;        memory[55925] <=  8'h62;        memory[55926] <=  8'h20;        memory[55927] <=  8'h6e;        memory[55928] <=  8'h76;        memory[55929] <=  8'h63;        memory[55930] <=  8'h61;        memory[55931] <=  8'h73;        memory[55932] <=  8'h67;        memory[55933] <=  8'h68;        memory[55934] <=  8'h75;        memory[55935] <=  8'h6a;        memory[55936] <=  8'h6c;        memory[55937] <=  8'h6b;        memory[55938] <=  8'h63;        memory[55939] <=  8'h78;        memory[55940] <=  8'h20;        memory[55941] <=  8'h6a;        memory[55942] <=  8'h6b;        memory[55943] <=  8'h68;        memory[55944] <=  8'h61;        memory[55945] <=  8'h73;        memory[55946] <=  8'h76;        memory[55947] <=  8'h64;        memory[55948] <=  8'h6e;        memory[55949] <=  8'h20;        memory[55950] <=  8'h62;        memory[55951] <=  8'h6e;        memory[55952] <=  8'h6d;        memory[55953] <=  8'h6b;        memory[55954] <=  8'h77;        memory[55955] <=  8'h64;        memory[55956] <=  8'h6f;        memory[55957] <=  8'h77;        memory[55958] <=  8'h69;        memory[55959] <=  8'h6f;        memory[55960] <=  8'h75;        memory[55961] <=  8'h69;        memory[55962] <=  8'h68;        memory[55963] <=  8'h62;        memory[55964] <=  8'h6e;        memory[55965] <=  8'h6b;        memory[55966] <=  8'h77;        memory[55967] <=  8'h69;        memory[55968] <=  8'h6f;        memory[55969] <=  8'h75;        memory[55970] <=  8'h71;        memory[55971] <=  8'h69;        memory[55972] <=  8'h79;        memory[55973] <=  8'h67;        memory[55974] <=  8'h6a;        memory[55975] <=  8'h64;        memory[55976] <=  8'h61;        memory[55977] <=  8'h76;        memory[55978] <=  8'h62;        memory[55979] <=  8'h6e;        memory[55980] <=  8'h6b;        memory[55981] <=  8'h6f;        memory[55982] <=  8'h70;        memory[55983] <=  8'h64;        memory[55984] <=  8'h76;        memory[55985] <=  8'h69;        memory[55986] <=  8'h6f;        memory[55987] <=  8'h75;        memory[55988] <=  8'h69;        memory[55989] <=  8'h48;        memory[55990] <=  8'h42;        memory[55991] <=  8'h6b;        memory[55992] <=  8'h64;        memory[55993] <=  8'h6e;        memory[55994] <=  8'h6c;        memory[55995] <=  8'h71;        memory[55996] <=  8'h6b;        memory[55997] <=  8'h6d;        memory[55998] <=  8'h6a;        memory[55999] <=  8'h70;        memory[56000] <=  8'h69;        memory[56001] <=  8'h6f;        memory[56002] <=  8'h68;        memory[56003] <=  8'h65;        memory[56004] <=  8'h66;        memory[56005] <=  8'h75;        memory[56006] <=  8'h67;        memory[56007] <=  8'h69;        memory[56008] <=  8'h73;        memory[56009] <=  8'h61;        memory[56010] <=  8'h62;        memory[56011] <=  8'h64;        memory[56012] <=  8'h6b;        memory[56013] <=  8'h6a;        memory[56014] <=  8'h6b;        memory[56015] <=  8'h6c;        memory[56016] <=  8'h6a;        memory[56017] <=  8'h69;        memory[56018] <=  8'h73;        memory[56019] <=  8'h6f;        memory[56020] <=  8'h71;        memory[56021] <=  8'h68;        memory[56022] <=  8'h77;        memory[56023] <=  8'h67;        memory[56024] <=  8'h69;        memory[56025] <=  8'h79;        memory[56026] <=  8'h6a;        memory[56027] <=  8'h64;        memory[56028] <=  8'h76;        memory[56029] <=  8'h62;        memory[56030] <=  8'h6e;        memory[56031] <=  8'h61;        memory[56032] <=  8'h73;        memory[56033] <=  8'h66;        memory[56034] <=  8'h6c;        memory[56035] <=  8'h6b;        memory[56036] <=  8'h64;        memory[56037] <=  8'h6a;        memory[56038] <=  8'h68;        memory[56039] <=  8'h63;        memory[56040] <=  8'h67;        memory[56041] <=  8'h6a;        memory[56042] <=  8'h76;        memory[56043] <=  8'h73;        memory[56044] <=  8'h64;        memory[56045] <=  8'h62;        memory[56046] <=  8'h62;        memory[56047] <=  8'h61;        memory[56048] <=  8'h72;        memory[56049] <=  8'h62;        memory[56050] <=  8'h62;        memory[56051] <=  8'h73;        memory[56052] <=  8'h62;        memory[56053] <=  8'h67;        memory[56054] <=  8'h73;        memory[56055] <=  8'h66;        memory[56056] <=  8'h67;        memory[56057] <=  8'h61;        memory[56058] <=  8'h68;        memory[56059] <=  8'h66;        memory[56060] <=  8'h73;        memory[56061] <=  8'h68;        memory[56062] <=  8'h61;        memory[56063] <=  8'h66;        memory[56064] <=  8'h73;        memory[56065] <=  8'h66;        memory[56066] <=  8'h68;        memory[56067] <=  8'h61;        memory[56068] <=  8'h69;        memory[56069] <=  8'h64;        memory[56070] <=  8'h75;        memory[56071] <=  8'h67;        memory[56072] <=  8'h64;        memory[56073] <=  8'h77;        memory[56074] <=  8'h62;        memory[56075] <=  8'h61;        memory[56076] <=  8'h62;        memory[56077] <=  8'h72;        memory[56078] <=  8'h62;        memory[56079] <=  8'h61;        memory[56080] <=  8'h62;        memory[56081] <=  8'h62;        memory[56082] <=  8'h74;        memory[56083] <=  8'h62;        memory[56084] <=  8'h62;        memory[56085] <=  8'h62;        memory[56086] <=  8'h62;        memory[56087] <=  8'h62;        memory[56088] <=  8'h62;        memory[56089] <=  8'h62;        memory[56090] <=  8'h62;        memory[56091] <=  8'h61;        memory[56092] <=  8'h62;        memory[56093] <=  8'h62;        memory[56094] <=  8'h72;        memory[56095] <=  8'h74;        memory[56096] <=  8'h62;        memory[56097] <=  8'h62;        memory[56098] <=  8'h61;        memory[56099] <=  8'h62;        memory[56100] <=  8'h72;        memory[56101] <=  8'h62;        memory[56102] <=  8'h74;        memory[56103] <=  8'h62;        memory[56104] <=  8'h62;        memory[56105] <=  8'h62;        memory[56106] <=  8'h63;        memory[56107] <=  8'h61;        memory[56108] <=  8'h72;        memory[56109] <=  8'h74;        memory[56110] <=  8'h73;        memory[56111] <=  8'h62;        memory[56112] <=  8'h61;        memory[56113] <=  8'h72;        memory[56114] <=  8'h74;        memory[56115] <=  8'h74;        memory[56116] <=  8'h62;        memory[56117] <=  8'h61;        memory[56118] <=  8'h72;        memory[56119] <=  8'h74;        memory[56120] <=  8'h78;        memory[56121] <=  8'h61;        memory[56122] <=  8'h74;        memory[56123] <=  8'h6b;        memory[56124] <=  8'h73;        memory[56125] <=  8'h68;        memory[56126] <=  8'h63;        memory[56127] <=  8'h66;        memory[56128] <=  8'h69;        memory[56129] <=  8'h77;        memory[56130] <=  8'h68;        memory[56131] <=  8'h61;        memory[56132] <=  8'h74;        memory[56133] <=  8'h61;        memory[56134] <=  8'h6e;        memory[56135] <=  8'h61;        memory[56136] <=  8'h62;        memory[56137] <=  8'h61;        memory[56138] <=  8'h63;        memory[56139] <=  8'h61;        memory[56140] <=  8'h74;        memory[56141] <=  8'h61;        memory[56142] <=  8'h62;        memory[56143] <=  8'h61;        memory[56144] <=  8'h72;        memory[56145] <=  8'h63;        memory[56146] <=  8'h61;        memory[56147] <=  8'h68;        memory[56148] <=  8'h64;        memory[56149] <=  8'h75;        memory[56150] <=  8'h63;        memory[56151] <=  8'h74;        memory[56152] <=  8'h61;        memory[56153] <=  8'h64;        memory[56154] <=  8'h61;        memory[56155] <=  8'h61;        memory[56156] <=  8'h63;        memory[56157] <=  8'h61;        memory[56158] <=  8'h72;        memory[56159] <=  8'h63;        memory[56160] <=  8'h74;        memory[56161] <=  8'h72;        memory[56162] <=  8'h63;        memory[56163] <=  8'h61;        memory[56164] <=  8'h74;        memory[56165] <=  8'h72;        memory[56166] <=  8'h63;        memory[56167] <=  8'h61;        memory[56168] <=  8'h74;        memory[56169] <=  8'h63;        memory[56170] <=  8'h62;        memory[56171] <=  8'h61;        memory[56172] <=  8'h74;        memory[56173] <=  8'h62;        memory[56174] <=  8'h72;        memory[56175] <=  8'h63;        memory[56176] <=  8'h61;        memory[56177] <=  8'h74;        memory[56178] <=  8'h72;        memory[56179] <=  8'h6e;        memory[56180] <=  8'h62;        memory[56181] <=  8'h61;        memory[56182] <=  8'h63;        memory[56183] <=  8'h61;        memory[56184] <=  8'h74;        memory[56185] <=  8'h79;        memory[56186] <=  8'h73;        memory[56187] <=  8'h6e;        memory[56188] <=  8'h63;        memory[56189] <=  8'h74;        memory[56190] <=  8'h61;        memory[56191] <=  8'h6e;        memory[56192] <=  8'h62;        memory[56193] <=  8'h61;        memory[56194] <=  8'h63;        memory[56195] <=  8'h72;        memory[56196] <=  8'h6e;        memory[56197] <=  8'h74;        memory[56198] <=  8'h61;        memory[56199] <=  8'h62;        memory[56200] <=  8'h74;        memory[56201] <=  8'h6e;        memory[56202] <=  8'h61;        memory[56203] <=  8'h72;        memory[56204] <=  8'h62;        memory[56205] <=  8'h78;        memory[56206] <=  8'h74;        memory[56207] <=  8'h61;        memory[56208] <=  8'h72;        memory[56209] <=  8'h62;        memory[56210] <=  8'h61;        memory[56211] <=  8'h72;        memory[56212] <=  8'h74;        memory[56213] <=  8'h74;        memory[56214] <=  8'h62;        memory[56215] <=  8'h61;        memory[56216] <=  8'h72;        memory[56217] <=  8'h74;        memory[56218] <=  8'h78;        memory[56219] <=  8'h61;        memory[56220] <=  8'h74;        memory[56221] <=  8'h6b;        memory[56222] <=  8'h73;        memory[56223] <=  8'h68;        memory[56224] <=  8'h63;        memory[56225] <=  8'h66;        memory[56226] <=  8'h69;        memory[56227] <=  8'h77;        memory[56228] <=  8'h68;        memory[56229] <=  8'h61;        memory[56230] <=  8'h74;        memory[56231] <=  8'h61;        memory[56232] <=  8'h6e;        memory[56233] <=  8'h61;        memory[56234] <=  8'h62;        memory[56235] <=  8'h61;        memory[56236] <=  8'h63;        memory[56237] <=  8'h61;        memory[56238] <=  8'h74;        memory[56239] <=  8'h61;        memory[56240] <=  8'h62;        memory[56241] <=  8'h61;        memory[56242] <=  8'h72;        memory[56243] <=  8'h63;        memory[56244] <=  8'h61;        memory[56245] <=  8'h68;        memory[56246] <=  8'h64;        memory[56247] <=  8'h75;        memory[56248] <=  8'h63;        memory[56249] <=  8'h74;        memory[56250] <=  8'h61;        memory[56251] <=  8'h64;        memory[56252] <=  8'h61;        memory[56253] <=  8'h61;        memory[56254] <=  8'h63;        memory[56255] <=  8'h61;        memory[56256] <=  8'h72;        memory[56257] <=  8'h63;        memory[56258] <=  8'h74;        memory[56259] <=  8'h72;        memory[56260] <=  8'h63;        memory[56261] <=  8'h61;        memory[56262] <=  8'h74;        memory[56263] <=  8'h72;        memory[56264] <=  8'h63;        memory[56265] <=  8'h61;        memory[56266] <=  8'h74;        memory[56267] <=  8'h63;        memory[56268] <=  8'h62;        memory[56269] <=  8'h61;        memory[56270] <=  8'h74;        memory[56271] <=  8'h62;        memory[56272] <=  8'h72;        memory[56273] <=  8'h63;        memory[56274] <=  8'h61;        memory[56275] <=  8'h74;        memory[56276] <=  8'h72;        memory[56277] <=  8'h6e;        memory[56278] <=  8'h62;        memory[56279] <=  8'h61;        memory[56280] <=  8'h63;        memory[56281] <=  8'h61;        memory[56282] <=  8'h74;        memory[56283] <=  8'h79;        memory[56284] <=  8'h73;        memory[56285] <=  8'h6e;        memory[56286] <=  8'h63;        memory[56287] <=  8'h74;        memory[56288] <=  8'h61;        memory[56289] <=  8'h6e;        memory[56290] <=  8'h62;        memory[56291] <=  8'h61;        memory[56292] <=  8'h63;        memory[56293] <=  8'h72;        memory[56294] <=  8'h6e;        memory[56295] <=  8'h74;        memory[56296] <=  8'h61;        memory[56297] <=  8'h62;        memory[56298] <=  8'h74;        memory[56299] <=  8'h6e;        memory[56300] <=  8'h61;        memory[56301] <=  8'h72;        memory[56302] <=  8'h62;        memory[56303] <=  8'h78;        memory[56304] <=  8'h74;        memory[56305] <=  8'h61;        memory[56306] <=  8'h72;        memory[56307] <=  8'h62;        memory[56308] <=  8'h61;        memory[56309] <=  8'h72;        memory[56310] <=  8'h74;        memory[56311] <=  8'h74;        memory[56312] <=  8'h62;        memory[56313] <=  8'h61;        memory[56314] <=  8'h72;        memory[56315] <=  8'h74;        memory[56316] <=  8'h78;        memory[56317] <=  8'h61;        memory[56318] <=  8'h74;        memory[56319] <=  8'h6b;        memory[56320] <=  8'h73;        memory[56321] <=  8'h68;        memory[56322] <=  8'h63;        memory[56323] <=  8'h66;        memory[56324] <=  8'h69;        memory[56325] <=  8'h77;        memory[56326] <=  8'h68;        memory[56327] <=  8'h61;        memory[56328] <=  8'h74;        memory[56329] <=  8'h61;        memory[56330] <=  8'h6e;        memory[56331] <=  8'h61;        memory[56332] <=  8'h62;        memory[56333] <=  8'h61;        memory[56334] <=  8'h63;        memory[56335] <=  8'h61;        memory[56336] <=  8'h74;        memory[56337] <=  8'h61;        memory[56338] <=  8'h62;        memory[56339] <=  8'h61;        memory[56340] <=  8'h72;        memory[56341] <=  8'h63;        memory[56342] <=  8'h61;        memory[56343] <=  8'h68;        memory[56344] <=  8'h64;        memory[56345] <=  8'h75;        memory[56346] <=  8'h63;        memory[56347] <=  8'h74;        memory[56348] <=  8'h61;        memory[56349] <=  8'h64;        memory[56350] <=  8'h61;        memory[56351] <=  8'h61;        memory[56352] <=  8'h63;        memory[56353] <=  8'h61;        memory[56354] <=  8'h72;        memory[56355] <=  8'h63;        memory[56356] <=  8'h74;        memory[56357] <=  8'h72;        memory[56358] <=  8'h63;        memory[56359] <=  8'h61;        memory[56360] <=  8'h74;        memory[56361] <=  8'h72;        memory[56362] <=  8'h63;        memory[56363] <=  8'h61;        memory[56364] <=  8'h74;        memory[56365] <=  8'h63;        memory[56366] <=  8'h62;        memory[56367] <=  8'h61;        memory[56368] <=  8'h74;        memory[56369] <=  8'h62;        memory[56370] <=  8'h72;        memory[56371] <=  8'h63;        memory[56372] <=  8'h61;        memory[56373] <=  8'h74;        memory[56374] <=  8'h72;        memory[56375] <=  8'h6e;        memory[56376] <=  8'h62;        memory[56377] <=  8'h61;        memory[56378] <=  8'h63;        memory[56379] <=  8'h61;        memory[56380] <=  8'h74;        memory[56381] <=  8'h79;        memory[56382] <=  8'h73;        memory[56383] <=  8'h6e;        memory[56384] <=  8'h63;        memory[56385] <=  8'h74;        memory[56386] <=  8'h61;        memory[56387] <=  8'h6e;        memory[56388] <=  8'h62;        memory[56389] <=  8'h61;        memory[56390] <=  8'h63;        memory[56391] <=  8'h72;        memory[56392] <=  8'h6e;        memory[56393] <=  8'h74;        memory[56394] <=  8'h61;        memory[56395] <=  8'h62;        memory[56396] <=  8'h74;        memory[56397] <=  8'h6e;        memory[56398] <=  8'h61;        memory[56399] <=  8'h72;        memory[56400] <=  8'h62;        memory[56401] <=  8'h78;        memory[56402] <=  8'h74;        memory[56403] <=  8'h61;        memory[56404] <=  8'h72;        memory[56405] <=  8'h5d;        memory[56406] <=  8'h5d;        memory[56407] <=  8'h65;        memory[56408] <=  8'h66;        memory[56409] <=  8'h77;        memory[56410] <=  8'h65;        memory[56411] <=  8'h5d;        memory[56412] <=  8'h65;        memory[56413] <=  8'h67;        memory[56414] <=  8'h73;        memory[56415] <=  8'h67;        memory[56416] <=  8'h66;        memory[56417] <=  8'h62;        memory[56418] <=  8'h61;        memory[56419] <=  8'h72;        memory[56420] <=  8'h74;        memory[56421] <=  8'h74;        memory[56422] <=  8'h62;        memory[56423] <=  8'h61;        memory[56424] <=  8'h72;        memory[56425] <=  8'h74;        memory[56426] <=  8'h78;        memory[56427] <=  8'h61;        memory[56428] <=  8'h74;        memory[56429] <=  8'h6b;        memory[56430] <=  8'h73;        memory[56431] <=  8'h68;        memory[56432] <=  8'h63;        memory[56433] <=  8'h66;        memory[56434] <=  8'h69;        memory[56435] <=  8'h77;        memory[56436] <=  8'h68;        memory[56437] <=  8'h61;        memory[56438] <=  8'h74;        memory[56439] <=  8'h61;        memory[56440] <=  8'h6e;        memory[56441] <=  8'h61;        memory[56442] <=  8'h62;        memory[56443] <=  8'h61;        memory[56444] <=  8'h63;        memory[56445] <=  8'h61;        memory[56446] <=  8'h74;        memory[56447] <=  8'h61;        memory[56448] <=  8'h62;        memory[56449] <=  8'h61;        memory[56450] <=  8'h72;        memory[56451] <=  8'h63;        memory[56452] <=  8'h61;        memory[56453] <=  8'h68;        memory[56454] <=  8'h64;        memory[56455] <=  8'h75;        memory[56456] <=  8'h63;        memory[56457] <=  8'h74;        memory[56458] <=  8'h61;        memory[56459] <=  8'h64;        memory[56460] <=  8'h61;        memory[56461] <=  8'h61;        memory[56462] <=  8'h63;        memory[56463] <=  8'h61;        memory[56464] <=  8'h72;        memory[56465] <=  8'h63;        memory[56466] <=  8'h74;        memory[56467] <=  8'h72;        memory[56468] <=  8'h63;        memory[56469] <=  8'h61;        memory[56470] <=  8'h74;        memory[56471] <=  8'h72;        memory[56472] <=  8'h63;        memory[56473] <=  8'h61;        memory[56474] <=  8'h74;        memory[56475] <=  8'h63;        memory[56476] <=  8'h62;        memory[56477] <=  8'h61;        memory[56478] <=  8'h74;        memory[56479] <=  8'h62;        memory[56480] <=  8'h72;        memory[56481] <=  8'h63;        memory[56482] <=  8'h61;        memory[56483] <=  8'h74;        memory[56484] <=  8'h72;        memory[56485] <=  8'h6e;        memory[56486] <=  8'h62;        memory[56487] <=  8'h61;        memory[56488] <=  8'h63;        memory[56489] <=  8'h61;        memory[56490] <=  8'h74;        memory[56491] <=  8'h79;        memory[56492] <=  8'h73;        memory[56493] <=  8'h6e;        memory[56494] <=  8'h63;        memory[56495] <=  8'h74;        memory[56496] <=  8'h61;        memory[56497] <=  8'h6e;        memory[56498] <=  8'h62;        memory[56499] <=  8'h61;        memory[56500] <=  8'h63;        memory[56501] <=  8'h72;        memory[56502] <=  8'h6e;        memory[56503] <=  8'h74;        memory[56504] <=  8'h61;        memory[56505] <=  8'h62;        memory[56506] <=  8'h74;        memory[56507] <=  8'h6e;        memory[56508] <=  8'h61;        memory[56509] <=  8'h72;        memory[56510] <=  8'h62;        memory[56511] <=  8'h78;        memory[56512] <=  8'h74;        memory[56513] <=  8'h61;        memory[56514] <=  8'h72;        memory[56515] <=  8'h62;        memory[56516] <=  8'h61;        memory[56517] <=  8'h72;        memory[56518] <=  8'h74;        memory[56519] <=  8'h74;        memory[56520] <=  8'h62;        memory[56521] <=  8'h61;        memory[56522] <=  8'h72;        memory[56523] <=  8'h74;        memory[56524] <=  8'h78;        memory[56525] <=  8'h61;        memory[56526] <=  8'h74;        memory[56527] <=  8'h6b;        memory[56528] <=  8'h73;        memory[56529] <=  8'h68;        memory[56530] <=  8'h63;        memory[56531] <=  8'h66;        memory[56532] <=  8'h69;        memory[56533] <=  8'h77;        memory[56534] <=  8'h68;        memory[56535] <=  8'h61;        memory[56536] <=  8'h74;        memory[56537] <=  8'h61;        memory[56538] <=  8'h6e;        memory[56539] <=  8'h61;        memory[56540] <=  8'h62;        memory[56541] <=  8'h61;        memory[56542] <=  8'h63;        memory[56543] <=  8'h61;        memory[56544] <=  8'h74;        memory[56545] <=  8'h61;        memory[56546] <=  8'h62;        memory[56547] <=  8'h61;        memory[56548] <=  8'h72;        memory[56549] <=  8'h63;        memory[56550] <=  8'h61;        memory[56551] <=  8'h68;        memory[56552] <=  8'h64;        memory[56553] <=  8'h75;        memory[56554] <=  8'h63;        memory[56555] <=  8'h74;        memory[56556] <=  8'h61;        memory[56557] <=  8'h64;        memory[56558] <=  8'h61;        memory[56559] <=  8'h61;        memory[56560] <=  8'h63;        memory[56561] <=  8'h61;        memory[56562] <=  8'h72;        memory[56563] <=  8'h63;        memory[56564] <=  8'h74;        memory[56565] <=  8'h72;        memory[56566] <=  8'h63;        memory[56567] <=  8'h61;        memory[56568] <=  8'h74;        memory[56569] <=  8'h72;        memory[56570] <=  8'h63;        memory[56571] <=  8'h61;        memory[56572] <=  8'h74;        memory[56573] <=  8'h63;        memory[56574] <=  8'h62;        memory[56575] <=  8'h61;        memory[56576] <=  8'h74;        memory[56577] <=  8'h62;        memory[56578] <=  8'h72;        memory[56579] <=  8'h63;        memory[56580] <=  8'h61;        memory[56581] <=  8'h74;        memory[56582] <=  8'h72;        memory[56583] <=  8'h6e;        memory[56584] <=  8'h62;        memory[56585] <=  8'h61;        memory[56586] <=  8'h63;        memory[56587] <=  8'h61;        memory[56588] <=  8'h74;        memory[56589] <=  8'h79;        memory[56590] <=  8'h73;        memory[56591] <=  8'h6e;        memory[56592] <=  8'h63;        memory[56593] <=  8'h74;        memory[56594] <=  8'h61;        memory[56595] <=  8'h6e;        memory[56596] <=  8'h62;        memory[56597] <=  8'h61;        memory[56598] <=  8'h63;        memory[56599] <=  8'h72;        memory[56600] <=  8'h6e;        memory[56601] <=  8'h74;        memory[56602] <=  8'h61;        memory[56603] <=  8'h62;        memory[56604] <=  8'h74;        memory[56605] <=  8'h6e;        memory[56606] <=  8'h61;        memory[56607] <=  8'h72;        memory[56608] <=  8'h62;        memory[56609] <=  8'h78;        memory[56610] <=  8'h74;        memory[56611] <=  8'h61;        memory[56612] <=  8'h72;        memory[56613] <=  8'h64;        memory[56614] <=  8'h66;        memory[56615] <=  8'h73;        memory[56616] <=  8'h67;        memory[56617] <=  8'h76;        memory[56618] <=  8'h68;        memory[56619] <=  8'h62;        memory[56620] <=  8'h6b;        memory[56621] <=  8'h6a;        memory[56622] <=  8'h6e;        memory[56623] <=  8'h6d;        memory[56624] <=  8'h62;        memory[56625] <=  8'h76;        memory[56626] <=  8'h78;        memory[56627] <=  8'h63;        memory[56628] <=  8'h73;        memory[56629] <=  8'h66;        memory[56630] <=  8'h72;        memory[56631] <=  8'h74;        memory[56632] <=  8'h79;        memory[56633] <=  8'h75;        memory[56634] <=  8'h6a;        memory[56635] <=  8'h6e;        memory[56636] <=  8'h62;        memory[56637] <=  8'h76;        memory[56638] <=  8'h63;        memory[56639] <=  8'h64;        memory[56640] <=  8'h74;        memory[56641] <=  8'h79;        memory[56642] <=  8'h75;        memory[56643] <=  8'h69;        memory[56644] <=  8'h6b;        memory[56645] <=  8'h6d;        memory[56646] <=  8'h6e;        memory[56647] <=  8'h62;        memory[56648] <=  8'h76;        memory[56649] <=  8'h63;        memory[56650] <=  8'h78;        memory[56651] <=  8'h73;        memory[56652] <=  8'h64;        memory[56653] <=  8'h72;        memory[56654] <=  8'h74;        memory[56655] <=  8'h79;        memory[56656] <=  8'h75;        memory[56657] <=  8'h69;        memory[56658] <=  8'h6b;        memory[56659] <=  8'h6d;        memory[56660] <=  8'h6e;        memory[56661] <=  8'h62;        memory[56662] <=  8'h76;        memory[56663] <=  8'h63;        memory[56664] <=  8'h73;        memory[56665] <=  8'h77;        memory[56666] <=  8'h33;        memory[56667] <=  8'h34;        memory[56668] <=  8'h35;        memory[56669] <=  8'h36;        memory[56670] <=  8'h37;        memory[56671] <=  8'h38;        memory[56672] <=  8'h69;        memory[56673] <=  8'h6b;        memory[56674] <=  8'h6d;        memory[56675] <=  8'h6e;        memory[56676] <=  8'h62;        memory[56677] <=  8'h76;        memory[56678] <=  8'h63;        memory[56679] <=  8'h64;        memory[56680] <=  8'h65;        memory[56681] <=  8'h72;        memory[56682] <=  8'h36;        memory[56683] <=  8'h37;        memory[56684] <=  8'h38;        memory[56685] <=  8'h69;        memory[56686] <=  8'h6f;        memory[56687] <=  8'h6b;        memory[56688] <=  8'h6a;        memory[56689] <=  8'h6e;        memory[56690] <=  8'h62;        memory[56691] <=  8'h76;        memory[56692] <=  8'h63;        memory[56693] <=  8'h64;        memory[56694] <=  8'h72;        memory[56695] <=  8'h74;        memory[56696] <=  8'h79;        memory[56697] <=  8'h75;        memory[56698] <=  8'h73;        memory[56699] <=  8'h6a;        memory[56700] <=  8'h63;        memory[56701] <=  8'h6e;        memory[56702] <=  8'h62;        memory[56703] <=  8'h64;        memory[56704] <=  8'h66;        memory[56705] <=  8'h73;        memory[56706] <=  8'h74;        memory[56707] <=  8'h79;        memory[56708] <=  8'h75;        memory[56709] <=  8'h61;        memory[56710] <=  8'h69;        memory[56711] <=  8'h6b;        memory[56712] <=  8'h78;        memory[56713] <=  8'h6d;        memory[56714] <=  8'h6e;        memory[56715] <=  8'h73;        memory[56716] <=  8'h6a;        memory[56717] <=  8'h6f;        memory[56718] <=  8'h64;        memory[56719] <=  8'h6c;        memory[56720] <=  8'h63;        memory[56721] <=  8'h78;        memory[56722] <=  8'h62;        memory[56723] <=  8'h61;        memory[56724] <=  8'h72;        memory[56725] <=  8'h74;        memory[56726] <=  8'h78;        memory[56727] <=  8'h61;        memory[56728] <=  8'h74;        memory[56729] <=  8'h6b;        memory[56730] <=  8'h73;        memory[56731] <=  8'h68;        memory[56732] <=  8'h63;        memory[56733] <=  8'h66;        memory[56734] <=  8'h69;        memory[56735] <=  8'h77;        memory[56736] <=  8'h68;        memory[56737] <=  8'h61;        memory[56738] <=  8'h74;        memory[56739] <=  8'h61;        memory[56740] <=  8'h6e;        memory[56741] <=  8'h61;        memory[56742] <=  8'h62;        memory[56743] <=  8'h61;        memory[56744] <=  8'h63;        memory[56745] <=  8'h61;        memory[56746] <=  8'h74;        memory[56747] <=  8'h61;        memory[56748] <=  8'h62;        memory[56749] <=  8'h61;        memory[56750] <=  8'h72;        memory[56751] <=  8'h63;        memory[56752] <=  8'h61;        memory[56753] <=  8'h68;        memory[56754] <=  8'h64;        memory[56755] <=  8'h75;        memory[56756] <=  8'h63;        memory[56757] <=  8'h74;        memory[56758] <=  8'h61;        memory[56759] <=  8'h64;        memory[56760] <=  8'h61;        memory[56761] <=  8'h61;        memory[56762] <=  8'h63;        memory[56763] <=  8'h61;        memory[56764] <=  8'h72;        memory[56765] <=  8'h62;        memory[56766] <=  8'h61;        memory[56767] <=  8'h72;        memory[56768] <=  8'h74;        memory[56769] <=  8'h78;        memory[56770] <=  8'h61;        memory[56771] <=  8'h74;        memory[56772] <=  8'h6b;        memory[56773] <=  8'h73;        memory[56774] <=  8'h68;        memory[56775] <=  8'h63;        memory[56776] <=  8'h66;        memory[56777] <=  8'h69;        memory[56778] <=  8'h77;        memory[56779] <=  8'h68;        memory[56780] <=  8'h61;        memory[56781] <=  8'h74;        memory[56782] <=  8'h61;        memory[56783] <=  8'h6e;        memory[56784] <=  8'h61;        memory[56785] <=  8'h62;        memory[56786] <=  8'h61;        memory[56787] <=  8'h63;        memory[56788] <=  8'h61;        memory[56789] <=  8'h74;        memory[56790] <=  8'h61;        memory[56791] <=  8'h62;        memory[56792] <=  8'h61;        memory[56793] <=  8'h72;        memory[56794] <=  8'h63;        memory[56795] <=  8'h61;        memory[56796] <=  8'h68;        memory[56797] <=  8'h64;        memory[56798] <=  8'h75;        memory[56799] <=  8'h63;        memory[56800] <=  8'h74;        memory[56801] <=  8'h61;        memory[56802] <=  8'h64;        memory[56803] <=  8'h61;        memory[56804] <=  8'h61;        memory[56805] <=  8'h63;        memory[56806] <=  8'h61;        memory[56807] <=  8'h72;        memory[56808] <=  8'h62;        memory[56809] <=  8'h61;        memory[56810] <=  8'h72;        memory[56811] <=  8'h74;        memory[56812] <=  8'h78;        memory[56813] <=  8'h61;        memory[56814] <=  8'h74;        memory[56815] <=  8'h6b;        memory[56816] <=  8'h73;        memory[56817] <=  8'h68;        memory[56818] <=  8'h63;        memory[56819] <=  8'h66;        memory[56820] <=  8'h69;        memory[56821] <=  8'h77;        memory[56822] <=  8'h68;        memory[56823] <=  8'h61;        memory[56824] <=  8'h74;        memory[56825] <=  8'h61;        memory[56826] <=  8'h6e;        memory[56827] <=  8'h61;        memory[56828] <=  8'h62;        memory[56829] <=  8'h61;        memory[56830] <=  8'h63;        memory[56831] <=  8'h61;        memory[56832] <=  8'h74;        memory[56833] <=  8'h61;        memory[56834] <=  8'h62;        memory[56835] <=  8'h61;        memory[56836] <=  8'h72;        memory[56837] <=  8'h63;        memory[56838] <=  8'h61;        memory[56839] <=  8'h68;        memory[56840] <=  8'h64;        memory[56841] <=  8'h75;        memory[56842] <=  8'h63;        memory[56843] <=  8'h74;        memory[56844] <=  8'h61;        memory[56845] <=  8'h64;        memory[56846] <=  8'h61;        memory[56847] <=  8'h61;        memory[56848] <=  8'h63;        memory[56849] <=  8'h61;        memory[56850] <=  8'h72;        memory[56851] <=  8'h62;        memory[56852] <=  8'h61;        memory[56853] <=  8'h72;        memory[56854] <=  8'h74;        memory[56855] <=  8'h78;        memory[56856] <=  8'h61;        memory[56857] <=  8'h74;        memory[56858] <=  8'h6b;        memory[56859] <=  8'h73;        memory[56860] <=  8'h68;        memory[56861] <=  8'h63;        memory[56862] <=  8'h66;        memory[56863] <=  8'h69;        memory[56864] <=  8'h77;        memory[56865] <=  8'h68;        memory[56866] <=  8'h61;        memory[56867] <=  8'h74;        memory[56868] <=  8'h61;        memory[56869] <=  8'h6e;        memory[56870] <=  8'h61;        memory[56871] <=  8'h62;        memory[56872] <=  8'h61;        memory[56873] <=  8'h63;        memory[56874] <=  8'h61;        memory[56875] <=  8'h74;        memory[56876] <=  8'h61;        memory[56877] <=  8'h62;        memory[56878] <=  8'h61;        memory[56879] <=  8'h72;        memory[56880] <=  8'h63;        memory[56881] <=  8'h61;        memory[56882] <=  8'h68;        memory[56883] <=  8'h64;        memory[56884] <=  8'h75;        memory[56885] <=  8'h63;        memory[56886] <=  8'h74;        memory[56887] <=  8'h61;        memory[56888] <=  8'h64;        memory[56889] <=  8'h61;        memory[56890] <=  8'h61;        memory[56891] <=  8'h63;        memory[56892] <=  8'h61;        memory[56893] <=  8'h72;        memory[56894] <=  8'h62;        memory[56895] <=  8'h61;        memory[56896] <=  8'h72;        memory[56897] <=  8'h74;        memory[56898] <=  8'h78;        memory[56899] <=  8'h61;        memory[56900] <=  8'h74;        memory[56901] <=  8'h6b;        memory[56902] <=  8'h73;        memory[56903] <=  8'h68;        memory[56904] <=  8'h63;        memory[56905] <=  8'h66;        memory[56906] <=  8'h69;        memory[56907] <=  8'h77;        memory[56908] <=  8'h68;        memory[56909] <=  8'h61;        memory[56910] <=  8'h74;        memory[56911] <=  8'h61;        memory[56912] <=  8'h6e;        memory[56913] <=  8'h61;        memory[56914] <=  8'h62;        memory[56915] <=  8'h61;        memory[56916] <=  8'h63;        memory[56917] <=  8'h61;        memory[56918] <=  8'h74;        memory[56919] <=  8'h61;        memory[56920] <=  8'h62;        memory[56921] <=  8'h61;        memory[56922] <=  8'h72;        memory[56923] <=  8'h63;        memory[56924] <=  8'h61;        memory[56925] <=  8'h68;        memory[56926] <=  8'h64;        memory[56927] <=  8'h75;        memory[56928] <=  8'h63;        memory[56929] <=  8'h74;        memory[56930] <=  8'h61;        memory[56931] <=  8'h64;        memory[56932] <=  8'h61;        memory[56933] <=  8'h61;        memory[56934] <=  8'h63;        memory[56935] <=  8'h61;        memory[56936] <=  8'h72;        memory[56937] <=  8'h62;        memory[56938] <=  8'h61;        memory[56939] <=  8'h72;        memory[56940] <=  8'h74;        memory[56941] <=  8'h78;        memory[56942] <=  8'h61;        memory[56943] <=  8'h74;        memory[56944] <=  8'h6b;        memory[56945] <=  8'h73;        memory[56946] <=  8'h68;        memory[56947] <=  8'h63;        memory[56948] <=  8'h66;        memory[56949] <=  8'h69;        memory[56950] <=  8'h77;        memory[56951] <=  8'h68;        memory[56952] <=  8'h61;        memory[56953] <=  8'h74;        memory[56954] <=  8'h61;        memory[56955] <=  8'h6e;        memory[56956] <=  8'h61;        memory[56957] <=  8'h62;        memory[56958] <=  8'h61;        memory[56959] <=  8'h63;        memory[56960] <=  8'h61;        memory[56961] <=  8'h74;        memory[56962] <=  8'h61;        memory[56963] <=  8'h62;        memory[56964] <=  8'h61;        memory[56965] <=  8'h72;        memory[56966] <=  8'h63;        memory[56967] <=  8'h61;        memory[56968] <=  8'h68;        memory[56969] <=  8'h64;        memory[56970] <=  8'h75;        memory[56971] <=  8'h63;        memory[56972] <=  8'h74;        memory[56973] <=  8'h61;        memory[56974] <=  8'h64;        memory[56975] <=  8'h61;        memory[56976] <=  8'h61;        memory[56977] <=  8'h63;        memory[56978] <=  8'h61;        memory[56979] <=  8'h72;        memory[56980] <=  8'h62;        memory[56981] <=  8'h61;        memory[56982] <=  8'h72;        memory[56983] <=  8'h74;        memory[56984] <=  8'h78;        memory[56985] <=  8'h61;        memory[56986] <=  8'h74;        memory[56987] <=  8'h6b;        memory[56988] <=  8'h73;        memory[56989] <=  8'h68;        memory[56990] <=  8'h63;        memory[56991] <=  8'h66;        memory[56992] <=  8'h69;        memory[56993] <=  8'h77;        memory[56994] <=  8'h68;        memory[56995] <=  8'h61;        memory[56996] <=  8'h74;        memory[56997] <=  8'h61;        memory[56998] <=  8'h6e;        memory[56999] <=  8'h61;        memory[57000] <=  8'h62;        memory[57001] <=  8'h61;        memory[57002] <=  8'h63;        memory[57003] <=  8'h61;        memory[57004] <=  8'h74;        memory[57005] <=  8'h61;        memory[57006] <=  8'h62;        memory[57007] <=  8'h61;        memory[57008] <=  8'h72;        memory[57009] <=  8'h63;        memory[57010] <=  8'h61;        memory[57011] <=  8'h68;        memory[57012] <=  8'h64;        memory[57013] <=  8'h75;        memory[57014] <=  8'h63;        memory[57015] <=  8'h74;        memory[57016] <=  8'h61;        memory[57017] <=  8'h64;        memory[57018] <=  8'h61;        memory[57019] <=  8'h61;        memory[57020] <=  8'h63;        memory[57021] <=  8'h61;        memory[57022] <=  8'h72;        memory[57023] <=  8'h62;        memory[57024] <=  8'h61;        memory[57025] <=  8'h72;        memory[57026] <=  8'h74;        memory[57027] <=  8'h78;        memory[57028] <=  8'h61;        memory[57029] <=  8'h74;        memory[57030] <=  8'h6b;        memory[57031] <=  8'h73;        memory[57032] <=  8'h68;        memory[57033] <=  8'h63;        memory[57034] <=  8'h66;        memory[57035] <=  8'h69;        memory[57036] <=  8'h77;        memory[57037] <=  8'h68;        memory[57038] <=  8'h61;        memory[57039] <=  8'h74;        memory[57040] <=  8'h61;        memory[57041] <=  8'h6e;        memory[57042] <=  8'h61;        memory[57043] <=  8'h62;        memory[57044] <=  8'h61;        memory[57045] <=  8'h63;        memory[57046] <=  8'h61;        memory[57047] <=  8'h74;        memory[57048] <=  8'h61;        memory[57049] <=  8'h62;        memory[57050] <=  8'h61;        memory[57051] <=  8'h72;        memory[57052] <=  8'h63;        memory[57053] <=  8'h61;        memory[57054] <=  8'h68;        memory[57055] <=  8'h64;        memory[57056] <=  8'h75;        memory[57057] <=  8'h63;        memory[57058] <=  8'h74;        memory[57059] <=  8'h61;        memory[57060] <=  8'h64;        memory[57061] <=  8'h61;        memory[57062] <=  8'h61;        memory[57063] <=  8'h63;        memory[57064] <=  8'h61;        memory[57065] <=  8'h72;        memory[57066] <=  8'h62;        memory[57067] <=  8'h61;        memory[57068] <=  8'h72;        memory[57069] <=  8'h74;        memory[57070] <=  8'h78;        memory[57071] <=  8'h61;        memory[57072] <=  8'h74;        memory[57073] <=  8'h6b;        memory[57074] <=  8'h73;        memory[57075] <=  8'h68;        memory[57076] <=  8'h63;        memory[57077] <=  8'h66;        memory[57078] <=  8'h69;        memory[57079] <=  8'h77;        memory[57080] <=  8'h68;        memory[57081] <=  8'h61;        memory[57082] <=  8'h74;        memory[57083] <=  8'h61;        memory[57084] <=  8'h6e;        memory[57085] <=  8'h61;        memory[57086] <=  8'h62;        memory[57087] <=  8'h61;        memory[57088] <=  8'h63;        memory[57089] <=  8'h61;        memory[57090] <=  8'h74;        memory[57091] <=  8'h61;        memory[57092] <=  8'h62;        memory[57093] <=  8'h61;        memory[57094] <=  8'h72;        memory[57095] <=  8'h63;        memory[57096] <=  8'h61;        memory[57097] <=  8'h68;        memory[57098] <=  8'h64;        memory[57099] <=  8'h75;        memory[57100] <=  8'h63;        memory[57101] <=  8'h74;        memory[57102] <=  8'h61;        memory[57103] <=  8'h64;        memory[57104] <=  8'h61;        memory[57105] <=  8'h61;        memory[57106] <=  8'h63;        memory[57107] <=  8'h61;        memory[57108] <=  8'h72;        memory[57109] <=  8'h62;        memory[57110] <=  8'h61;        memory[57111] <=  8'h72;        memory[57112] <=  8'h74;        memory[57113] <=  8'h74;        memory[57114] <=  8'h62;        memory[57115] <=  8'h61;        memory[57116] <=  8'h72;        memory[57117] <=  8'h74;        memory[57118] <=  8'h78;        memory[57119] <=  8'h61;        memory[57120] <=  8'h74;        memory[57121] <=  8'h6b;        memory[57122] <=  8'h73;        memory[57123] <=  8'h68;        memory[57124] <=  8'h63;        memory[57125] <=  8'h66;        memory[57126] <=  8'h69;        memory[57127] <=  8'h77;        memory[57128] <=  8'h68;        memory[57129] <=  8'h61;        memory[57130] <=  8'h74;        memory[57131] <=  8'h61;        memory[57132] <=  8'h6e;        memory[57133] <=  8'h61;        memory[57134] <=  8'h62;        memory[57135] <=  8'h61;        memory[57136] <=  8'h63;        memory[57137] <=  8'h61;        memory[57138] <=  8'h74;        memory[57139] <=  8'h61;        memory[57140] <=  8'h62;        memory[57141] <=  8'h61;        memory[57142] <=  8'h72;        memory[57143] <=  8'h63;        memory[57144] <=  8'h61;        memory[57145] <=  8'h68;        memory[57146] <=  8'h64;        memory[57147] <=  8'h75;        memory[57148] <=  8'h63;        memory[57149] <=  8'h74;        memory[57150] <=  8'h61;        memory[57151] <=  8'h64;        memory[57152] <=  8'h61;        memory[57153] <=  8'h61;        memory[57154] <=  8'h63;        memory[57155] <=  8'h61;        memory[57156] <=  8'h72;        memory[57157] <=  8'h63;        memory[57158] <=  8'h74;        memory[57159] <=  8'h72;        memory[57160] <=  8'h63;        memory[57161] <=  8'h61;        memory[57162] <=  8'h74;        memory[57163] <=  8'h72;        memory[57164] <=  8'h63;        memory[57165] <=  8'h61;        memory[57166] <=  8'h74;        memory[57167] <=  8'h63;        memory[57168] <=  8'h62;        memory[57169] <=  8'h61;        memory[57170] <=  8'h74;        memory[57171] <=  8'h62;        memory[57172] <=  8'h72;        memory[57173] <=  8'h63;        memory[57174] <=  8'h61;        memory[57175] <=  8'h72;        memory[57176] <=  8'h62;        memory[57177] <=  8'h78;        memory[57178] <=  8'h74;        memory[57179] <=  8'h61;        memory[57180] <=  8'h72;        memory[57181] <=  8'h64;        memory[57182] <=  8'h66;        memory[57183] <=  8'h73;        memory[57184] <=  8'h67;        memory[57185] <=  8'h76;        memory[57186] <=  8'h68;        memory[57187] <=  8'h62;        memory[57188] <=  8'h6b;        memory[57189] <=  8'h6a;        memory[57190] <=  8'h6e;        memory[57191] <=  8'h6d;        memory[57192] <=  8'h62;        memory[57193] <=  8'h76;        memory[57194] <=  8'h78;        memory[57195] <=  8'h63;        memory[57196] <=  8'h73;        memory[57197] <=  8'h66;        memory[57198] <=  8'h72;        memory[57199] <=  8'h74;        memory[57200] <=  8'h79;        memory[57201] <=  8'h75;        memory[57202] <=  8'h6a;        memory[57203] <=  8'h6e;        memory[57204] <=  8'h62;        memory[57205] <=  8'h76;        memory[57206] <=  8'h63;        memory[57207] <=  8'h64;        memory[57208] <=  8'h74;        memory[57209] <=  8'h79;        memory[57210] <=  8'h75;        memory[57211] <=  8'h69;        memory[57212] <=  8'h6b;        memory[57213] <=  8'h6d;        memory[57214] <=  8'h6e;        memory[57215] <=  8'h62;        memory[57216] <=  8'h76;        memory[57217] <=  8'h63;        memory[57218] <=  8'h78;        memory[57219] <=  8'h73;        memory[57220] <=  8'h64;        memory[57221] <=  8'h72;        memory[57222] <=  8'h74;        memory[57223] <=  8'h79;        memory[57224] <=  8'h75;        memory[57225] <=  8'h69;        memory[57226] <=  8'h6b;        memory[57227] <=  8'h6d;        memory[57228] <=  8'h6e;        memory[57229] <=  8'h62;        memory[57230] <=  8'h76;        memory[57231] <=  8'h63;        memory[57232] <=  8'h73;        memory[57233] <=  8'h77;        memory[57234] <=  8'h33;        memory[57235] <=  8'h34;        memory[57236] <=  8'h35;        memory[57237] <=  8'h36;        memory[57238] <=  8'h37;        memory[57239] <=  8'h38;        memory[57240] <=  8'h69;        memory[57241] <=  8'h6b;        memory[57242] <=  8'h6d;        memory[57243] <=  8'h6e;        memory[57244] <=  8'h62;        memory[57245] <=  8'h76;        memory[57246] <=  8'h63;        memory[57247] <=  8'h64;        memory[57248] <=  8'h65;        memory[57249] <=  8'h72;        memory[57250] <=  8'h36;        memory[57251] <=  8'h37;        memory[57252] <=  8'h38;        memory[57253] <=  8'h69;        memory[57254] <=  8'h6f;        memory[57255] <=  8'h6b;        memory[57256] <=  8'h6a;        memory[57257] <=  8'h6e;        memory[57258] <=  8'h62;        memory[57259] <=  8'h76;        memory[57260] <=  8'h63;        memory[57261] <=  8'h64;        memory[57262] <=  8'h72;        memory[57263] <=  8'h74;        memory[57264] <=  8'h79;        memory[57265] <=  8'h75;        memory[57266] <=  8'h73;        memory[57267] <=  8'h6a;        memory[57268] <=  8'h63;        memory[57269] <=  8'h6e;        memory[57270] <=  8'h62;        memory[57271] <=  8'h64;        memory[57272] <=  8'h66;        memory[57273] <=  8'h73;        memory[57274] <=  8'h74;        memory[57275] <=  8'h79;        memory[57276] <=  8'h75;        memory[57277] <=  8'h61;        memory[57278] <=  8'h69;        memory[57279] <=  8'h6b;        memory[57280] <=  8'h78;        memory[57281] <=  8'h6d;        memory[57282] <=  8'h6e;        memory[57283] <=  8'h73;        memory[57284] <=  8'h6a;        memory[57285] <=  8'h6f;        memory[57286] <=  8'h64;        memory[57287] <=  8'h6c;        memory[57288] <=  8'h63;        memory[57289] <=  8'h78;        memory[57290] <=  8'h2c;        memory[57291] <=  8'h6d;        memory[57292] <=  8'h73;        memory[57293] <=  8'h6b;        memory[57294] <=  8'h64;        memory[57295] <=  8'h6c;        memory[57296] <=  8'h70;        memory[57297] <=  8'h5b;        memory[57298] <=  8'h3b;        memory[57299] <=  8'h73;        memory[57300] <=  8'h6c;        memory[57301] <=  8'h64;        memory[57302] <=  8'h70;        memory[57303] <=  8'h76;        memory[57304] <=  8'h63;        memory[57305] <=  8'h5b;        memory[57306] <=  8'h78;        memory[57307] <=  8'h76;        memory[57308] <=  8'h63;        memory[57309] <=  8'h5b;        memory[57310] <=  8'h78;        memory[57311] <=  8'h70;        memory[57312] <=  8'h6f;        memory[57313] <=  8'h20;        memory[57314] <=  8'h62;        memory[57315] <=  8'h61;        memory[57316] <=  8'h72;        memory[57317] <=  8'h74;        memory[57318] <=  8'h74;        memory[57319] <=  8'h62;        memory[57320] <=  8'h61;        memory[57321] <=  8'h72;        memory[57322] <=  8'h74;        memory[57323] <=  8'h78;        memory[57324] <=  8'h61;        memory[57325] <=  8'h74;        memory[57326] <=  8'h6b;        memory[57327] <=  8'h73;        memory[57328] <=  8'h68;        memory[57329] <=  8'h63;        memory[57330] <=  8'h66;        memory[57331] <=  8'h69;        memory[57332] <=  8'h77;        memory[57333] <=  8'h68;        memory[57334] <=  8'h61;        memory[57335] <=  8'h69;        memory[57336] <=  8'h6a;        memory[57337] <=  8'h78;        memory[57338] <=  8'h5d;        memory[57339] <=  8'h65;        memory[57340] <=  8'h6b;        memory[57341] <=  8'h6f;        memory[57342] <=  8'h39;        memory[57343] <=  8'h64;        memory[57344] <=  8'h75;        memory[57345] <=  8'h38;        memory[57346] <=  8'h79;        memory[57347] <=  8'h20;        memory[57348] <=  8'h37;        memory[57349] <=  8'h63;        memory[57350] <=  8'h67;        memory[57351] <=  8'h78;        memory[57352] <=  8'h63;        memory[57353] <=  8'h75;        memory[57354] <=  8'h68;        memory[57355] <=  8'h69;        memory[57356] <=  8'h6a;        memory[57357] <=  8'h77;        memory[57358] <=  8'h69;        memory[57359] <=  8'h64;        memory[57360] <=  8'h66;        memory[57361] <=  8'h68;        memory[57362] <=  8'h75;        memory[57363] <=  8'h76;        memory[57364] <=  8'h64;        memory[57365] <=  8'h62;        memory[57366] <=  8'h66;        memory[57367] <=  8'h6a;        memory[57368] <=  8'h6e;        memory[57369] <=  8'h6b;        memory[57370] <=  8'h6a;        memory[57371] <=  8'h65;        memory[57372] <=  8'h38;        memory[57373] <=  8'h66;        memory[57374] <=  8'h37;        memory[57375] <=  8'h67;        memory[57376] <=  8'h79;        memory[57377] <=  8'h76;        memory[57378] <=  8'h63;        memory[57379] <=  8'h68;        memory[57380] <=  8'h69;        memory[57381] <=  8'h6a;        memory[57382] <=  8'h33;        memory[57383] <=  8'h65;        memory[57384] <=  8'h67;        memory[57385] <=  8'h79;        memory[57386] <=  8'h72;        memory[57387] <=  8'h64;        memory[57388] <=  8'h62;        memory[57389] <=  8'h6e;        memory[57390] <=  8'h63;        memory[57391] <=  8'h7a;        memory[57392] <=  8'h6a;        memory[57393] <=  8'h6f;        memory[57394] <=  8'h66;        memory[57395] <=  8'h78;        memory[57396] <=  8'h6a;        memory[57397] <=  8'h69;        memory[57398] <=  8'h63;        memory[57399] <=  8'h68;        memory[57400] <=  8'h62;        memory[57401] <=  8'h6e;        memory[57402] <=  8'h6d;        memory[57403] <=  8'h63;        memory[57404] <=  8'h73;        memory[57405] <=  8'h6c;        memory[57406] <=  8'h6b;        memory[57407] <=  8'h6a;        memory[57408] <=  8'h69;        memory[57409] <=  8'h68;        memory[57410] <=  8'h76;        memory[57411] <=  8'h75;        memory[57412] <=  8'h69;        memory[57413] <=  8'h64;        memory[57414] <=  8'h68;        memory[57415] <=  8'h75;        memory[57416] <=  8'h67;        memory[57417] <=  8'h79;        memory[57418] <=  8'h62;        memory[57419] <=  8'h68;        memory[57420] <=  8'h65;        memory[57421] <=  8'h6a;        memory[57422] <=  8'h72;        memory[57423] <=  8'h6b;        memory[57424] <=  8'h6a;        memory[57425] <=  8'h6f;        memory[57426] <=  8'h64;        memory[57427] <=  8'h67;        memory[57428] <=  8'h69;        memory[57429] <=  8'h75;        memory[57430] <=  8'h69;        memory[57431] <=  8'h67;        memory[57432] <=  8'h76;        memory[57433] <=  8'h79;        memory[57434] <=  8'h75;        memory[57435] <=  8'h67;        memory[57436] <=  8'h78;        memory[57437] <=  8'h68;        memory[57438] <=  8'h63;        memory[57439] <=  8'h20;        memory[57440] <=  8'h20;        memory[57441] <=  8'h20;        memory[57442] <=  8'h78;        memory[57443] <=  8'h76;        memory[57444] <=  8'h20;        memory[57445] <=  8'h63;        memory[57446] <=  8'h78;        memory[57447] <=  8'h67;        memory[57448] <=  8'h79;        memory[57449] <=  8'h63;        memory[57450] <=  8'h75;        memory[57451] <=  8'h68;        memory[57452] <=  8'h6a;        memory[57453] <=  8'h6b;        memory[57454] <=  8'h61;        memory[57455] <=  8'h6c;        memory[57456] <=  8'h78;        memory[57457] <=  8'h76;        memory[57458] <=  8'h70;        memory[57459] <=  8'h6f;        memory[57460] <=  8'h69;        memory[57461] <=  8'h6a;        memory[57462] <=  8'h69;        memory[57463] <=  8'h68;        memory[57464] <=  8'h6a;        memory[57465] <=  8'h62;        memory[57466] <=  8'h77;        memory[57467] <=  8'h65;        memory[57468] <=  8'h6e;        memory[57469] <=  8'h61;        memory[57470] <=  8'h66;        memory[57471] <=  8'h6d;        memory[57472] <=  8'h64;        memory[57473] <=  8'h6b;        memory[57474] <=  8'h6d;        memory[57475] <=  8'h76;        memory[57476] <=  8'h6c;        memory[57477] <=  8'h63;        memory[57478] <=  8'h6f;        memory[57479] <=  8'h64;        memory[57480] <=  8'h69;        memory[57481] <=  8'h75;        memory[57482] <=  8'h68;        memory[57483] <=  8'h73;        memory[57484] <=  8'h66;        memory[57485] <=  8'h65;        memory[57486] <=  8'h62;        memory[57487] <=  8'h6e;        memory[57488] <=  8'h64;        memory[57489] <=  8'h73;        memory[57490] <=  8'h63;        memory[57491] <=  8'h6b;        memory[57492] <=  8'h20;        memory[57493] <=  8'h78;        memory[57494] <=  8'h6a;        memory[57495] <=  8'h78;        memory[57496] <=  8'h63;        memory[57497] <=  8'h73;        memory[57498] <=  8'h64;        memory[57499] <=  8'h66;        memory[57500] <=  8'h6b;        memory[57501] <=  8'h64;        memory[57502] <=  8'h6e;        memory[57503] <=  8'h6d;        memory[57504] <=  8'h64;        memory[57505] <=  8'h73;        memory[57506] <=  8'h63;        memory[57507] <=  8'h6b;        memory[57508] <=  8'h78;        memory[57509] <=  8'h6c;        memory[57510] <=  8'h6f;        memory[57511] <=  8'h66;        memory[57512] <=  8'h6a;        memory[57513] <=  8'h69;        memory[57514] <=  8'h61;        memory[57515] <=  8'h62;        memory[57516] <=  8'h6e;        memory[57517] <=  8'h20;        memory[57518] <=  8'h78;        memory[57519] <=  8'h6b;        memory[57520] <=  8'h6d;        memory[57521] <=  8'h20;        memory[57522] <=  8'h6f;        memory[57523] <=  8'h63;        memory[57524] <=  8'h76;        memory[57525] <=  8'h73;        memory[57526] <=  8'h64;        memory[57527] <=  8'h69;        memory[57528] <=  8'h66;        memory[57529] <=  8'h68;        memory[57530] <=  8'h65;        memory[57531] <=  8'h71;        memory[57532] <=  8'h6a;        memory[57533] <=  8'h77;        memory[57534] <=  8'h62;        memory[57535] <=  8'h65;        memory[57536] <=  8'h6e;        memory[57537] <=  8'h20;        memory[57538] <=  8'h6d;        memory[57539] <=  8'h64;        memory[57540] <=  8'h73;        memory[57541] <=  8'h6c;        memory[57542] <=  8'h76;        memory[57543] <=  8'h6b;        memory[57544] <=  8'h63;        memory[57545] <=  8'h78;        memory[57546] <=  8'h20;        memory[57547] <=  8'h6f;        memory[57548] <=  8'h78;        memory[57549] <=  8'h69;        memory[57550] <=  8'h63;        memory[57551] <=  8'h6a;        memory[57552] <=  8'h76;        memory[57553] <=  8'h64;        memory[57554] <=  8'h66;        memory[57555] <=  8'h65;        memory[57556] <=  8'h71;        memory[57557] <=  8'h6e;        memory[57558] <=  8'h20;        memory[57559] <=  8'h64;        memory[57560] <=  8'h6d;        memory[57561] <=  8'h73;        memory[57562] <=  8'h6c;        memory[57563] <=  8'h63;        memory[57564] <=  8'h78;        memory[57565] <=  8'h6b;        memory[57566] <=  8'h20;        memory[57567] <=  8'h6f;        memory[57568] <=  8'h78;        memory[57569] <=  8'h63;        memory[57570] <=  8'h76;        memory[57571] <=  8'h6a;        memory[57572] <=  8'h64;        memory[57573] <=  8'h62;        memory[57574] <=  8'h71;        memory[57575] <=  8'h77;        memory[57576] <=  8'h65;        memory[57577] <=  8'h6e;        memory[57578] <=  8'h6d;        memory[57579] <=  8'h64;        memory[57580] <=  8'h6c;        memory[57581] <=  8'h73;        memory[57582] <=  8'h2c;        memory[57583] <=  8'h76;        memory[57584] <=  8'h63;        memory[57585] <=  8'h78;        memory[57586] <=  8'h20;        memory[57587] <=  8'h63;        memory[57588] <=  8'h6f;        memory[57589] <=  8'h69;        memory[57590] <=  8'h76;        memory[57591] <=  8'h68;        memory[57592] <=  8'h73;        memory[57593] <=  8'h64;        memory[57594] <=  8'h62;        memory[57595] <=  8'h71;        memory[57596] <=  8'h77;        memory[57597] <=  8'h65;        memory[57598] <=  8'h6e;        memory[57599] <=  8'h64;        memory[57600] <=  8'h6b;        memory[57601] <=  8'h73;        memory[57602] <=  8'h76;        memory[57603] <=  8'h6f;        memory[57604] <=  8'h63;        memory[57605] <=  8'h20;        memory[57606] <=  8'h76;        memory[57607] <=  8'h69;        memory[57608] <=  8'h75;        memory[57609] <=  8'h69;        memory[57610] <=  8'h68;        memory[57611] <=  8'h63;        memory[57612] <=  8'h78;        memory[57613] <=  8'h69;        memory[57614] <=  8'h6f;        memory[57615] <=  8'h76;        memory[57616] <=  8'h73;        memory[57617] <=  8'h64;        memory[57618] <=  8'h61;        memory[57619] <=  8'h64;        memory[57620] <=  8'h6e;        memory[57621] <=  8'h77;        memory[57622] <=  8'h71;        memory[57623] <=  8'h6b;        memory[57624] <=  8'h6c;        memory[57625] <=  8'h73;        memory[57626] <=  8'h76;        memory[57627] <=  8'h6e;        memory[57628] <=  8'h62;        memory[57629] <=  8'h20;        memory[57630] <=  8'h64;        memory[57631] <=  8'h66;        memory[57632] <=  8'h6a;        memory[57633] <=  8'h6b;        memory[57634] <=  8'h71;        memory[57635] <=  8'h64;        memory[57636] <=  8'h77;        memory[57637] <=  8'h65;        memory[57638] <=  8'h6e;        memory[57639] <=  8'h62;        memory[57640] <=  8'h20;        memory[57641] <=  8'h64;        memory[57642] <=  8'h73;        memory[57643] <=  8'h76;        memory[57644] <=  8'h68;        memory[57645] <=  8'h64;        memory[57646] <=  8'h61;        memory[57647] <=  8'h71;        memory[57648] <=  8'h77;        memory[57649] <=  8'h6a;        memory[57650] <=  8'h65;        memory[57651] <=  8'h6e;        memory[57652] <=  8'h64;        memory[57653] <=  8'h20;        memory[57654] <=  8'h61;        memory[57655] <=  8'h63;        memory[57656] <=  8'h62;        memory[57657] <=  8'h68;        memory[57658] <=  8'h64;        memory[57659] <=  8'h61;        memory[57660] <=  8'h77;        memory[57661] <=  8'h71;        memory[57662] <=  8'h6e;        memory[57663] <=  8'h20;        memory[57664] <=  8'h62;        memory[57665] <=  8'h73;        memory[57666] <=  8'h76;        memory[57667] <=  8'h61;        memory[57668] <=  8'h67;        memory[57669] <=  8'h76;        memory[57670] <=  8'h68;        memory[57671] <=  8'h67;        memory[57672] <=  8'h61;        memory[57673] <=  8'h73;        memory[57674] <=  8'h6a;        memory[57675] <=  8'h6b;        memory[57676] <=  8'h63;        memory[57677] <=  8'h78;        memory[57678] <=  8'h76;        memory[57679] <=  8'h6e;        memory[57680] <=  8'h73;        memory[57681] <=  8'h64;        memory[57682] <=  8'h20;        memory[57683] <=  8'h66;        memory[57684] <=  8'h62;        memory[57685] <=  8'h64;        memory[57686] <=  8'h61;        memory[57687] <=  8'h73;        memory[57688] <=  8'h76;        memory[57689] <=  8'h67;        memory[57690] <=  8'h63;        memory[57691] <=  8'h79;        memory[57692] <=  8'h7a;        memory[57693] <=  8'h78;        memory[57694] <=  8'h79;        memory[57695] <=  8'h75;        memory[57696] <=  8'h20;        memory[57697] <=  8'h69;        memory[57698] <=  8'h6a;        memory[57699] <=  8'h64;        memory[57700] <=  8'h66;        memory[57701] <=  8'h6b;        memory[57702] <=  8'h61;        memory[57703] <=  8'h64;        memory[57704] <=  8'h63;        memory[57705] <=  8'h78;        memory[57706] <=  8'h68;        memory[57707] <=  8'h20;        memory[57708] <=  8'h67;        memory[57709] <=  8'h61;        memory[57710] <=  8'h68;        memory[57711] <=  8'h75;        memory[57712] <=  8'h64;        memory[57713] <=  8'h73;        memory[57714] <=  8'h69;        memory[57715] <=  8'h6a;        memory[57716] <=  8'h61;        memory[57717] <=  8'h6b;        memory[57718] <=  8'h63;        memory[57719] <=  8'h62;        memory[57720] <=  8'h61;        memory[57721] <=  8'h72;        memory[57722] <=  8'h73;        memory[57723] <=  8'h68;        memory[57724] <=  8'h64;        memory[57725] <=  8'h66;        memory[57726] <=  8'h67;        memory[57727] <=  8'h73;        memory[57728] <=  8'h68;        memory[57729] <=  8'h64;        memory[57730] <=  8'h66;        memory[57731] <=  8'h68;        memory[57732] <=  8'h64;        memory[57733] <=  8'h6a;        memory[57734] <=  8'h68;        memory[57735] <=  8'h62;        memory[57736] <=  8'h67;        memory[57737] <=  8'h63;        memory[57738] <=  8'h61;        memory[57739] <=  8'h66;        memory[57740] <=  8'h73;        memory[57741] <=  8'h79;        memory[57742] <=  8'h67;        memory[57743] <=  8'h6b;        memory[57744] <=  8'h75;        memory[57745] <=  8'h64;        memory[57746] <=  8'h68;        memory[57747] <=  8'h62;        memory[57748] <=  8'h77;        memory[57749] <=  8'h76;        memory[57750] <=  8'h67;        memory[57751] <=  8'h61;        memory[57752] <=  8'h66;        memory[57753] <=  8'h64;        memory[57754] <=  8'h74;        memory[57755] <=  8'h75;        memory[57756] <=  8'h66;        memory[57757] <=  8'h79;        memory[57758] <=  8'h67;        memory[57759] <=  8'h69;        memory[57760] <=  8'h75;        memory[57761] <=  8'h68;        memory[57762] <=  8'h6c;        memory[57763] <=  8'h6a;        memory[57764] <=  8'h62;        memory[57765] <=  8'h6b;        memory[57766] <=  8'h68;        memory[57767] <=  8'h76;        memory[57768] <=  8'h67;        memory[57769] <=  8'h63;        memory[57770] <=  8'h66;        memory[57771] <=  8'h78;        memory[57772] <=  8'h64;        memory[57773] <=  8'h74;        memory[57774] <=  8'h75;        memory[57775] <=  8'h79;        memory[57776] <=  8'h69;        memory[57777] <=  8'h75;        memory[57778] <=  8'h68;        memory[57779] <=  8'h6c;        memory[57780] <=  8'h6a;        memory[57781] <=  8'h6b;        memory[57782] <=  8'h67;        memory[57783] <=  8'h6a;        memory[57784] <=  8'h63;        memory[57785] <=  8'h66;        memory[57786] <=  8'h68;        memory[57787] <=  8'h64;        memory[57788] <=  8'h67;        memory[57789] <=  8'h72;        memory[57790] <=  8'h79;        memory[57791] <=  8'h74;        memory[57792] <=  8'h66;        memory[57793] <=  8'h75;        memory[57794] <=  8'h79;        memory[57795] <=  8'h69;        memory[57796] <=  8'h68;        memory[57797] <=  8'h6c;        memory[57798] <=  8'h62;        memory[57799] <=  8'h6d;        memory[57800] <=  8'h76;        memory[57801] <=  8'h6e;        memory[57802] <=  8'h63;        memory[57803] <=  8'h66;        memory[57804] <=  8'h68;        memory[57805] <=  8'h64;        memory[57806] <=  8'h74;        memory[57807] <=  8'h75;        memory[57808] <=  8'h67;        memory[57809] <=  8'h79;        memory[57810] <=  8'h69;        memory[57811] <=  8'h68;        memory[57812] <=  8'h75;        memory[57813] <=  8'h6a;        memory[57814] <=  8'h6c;        memory[57815] <=  8'h62;        memory[57816] <=  8'h6d;        memory[57817] <=  8'h76;        memory[57818] <=  8'h6e;        memory[57819] <=  8'h63;        memory[57820] <=  8'h66;        memory[57821] <=  8'h68;        memory[57822] <=  8'h67;        memory[57823] <=  8'h79;        memory[57824] <=  8'h68;        memory[57825] <=  8'h75;        memory[57826] <=  8'h6a;        memory[57827] <=  8'h6e;        memory[57828] <=  8'h2c;        memory[57829] <=  8'h62;        memory[57830] <=  8'h6e;        memory[57831] <=  8'h6d;        memory[57832] <=  8'h76;        memory[57833] <=  8'h6e;        memory[57834] <=  8'h63;        memory[57835] <=  8'h66;        memory[57836] <=  8'h68;        memory[57837] <=  8'h74;        memory[57838] <=  8'h79;        memory[57839] <=  8'h69;        memory[57840] <=  8'h75;        memory[57841] <=  8'h6c;        memory[57842] <=  8'h6a;        memory[57843] <=  8'h62;        memory[57844] <=  8'h6d;        memory[57845] <=  8'h76;        memory[57846] <=  8'h6e;        memory[57847] <=  8'h63;        memory[57848] <=  8'h66;        memory[57849] <=  8'h74;        memory[57850] <=  8'h75;        memory[57851] <=  8'h79;        memory[57852] <=  8'h69;        memory[57853] <=  8'h68;        memory[57854] <=  8'h6b;        memory[57855] <=  8'h62;        memory[57856] <=  8'h76;        memory[57857] <=  8'h63;        memory[57858] <=  8'h66;        memory[57859] <=  8'h67;        memory[57860] <=  8'h74;        memory[57861] <=  8'h75;        memory[57862] <=  8'h79;        memory[57863] <=  8'h69;        memory[57864] <=  8'h75;        memory[57865] <=  8'h68;        memory[57866] <=  8'h6a;        memory[57867] <=  8'h6b;        memory[57868] <=  8'h62;        memory[57869] <=  8'h76;        memory[57870] <=  8'h63;        memory[57871] <=  8'h66;        memory[57872] <=  8'h74;        memory[57873] <=  8'h75;        memory[57874] <=  8'h79;        memory[57875] <=  8'h69;        memory[57876] <=  8'h75;        memory[57877] <=  8'h6a;        memory[57878] <=  8'h6b;        memory[57879] <=  8'h6e;        memory[57880] <=  8'h62;        memory[57881] <=  8'h76;        memory[57882] <=  8'h67;        memory[57883] <=  8'h66;        memory[57884] <=  8'h74;        memory[57885] <=  8'h79;        memory[57886] <=  8'h75;        memory[57887] <=  8'h75;        memory[57888] <=  8'h69;        memory[57889] <=  8'h6a;        memory[57890] <=  8'h6b;        memory[57891] <=  8'h68;        memory[57892] <=  8'h62;        memory[57893] <=  8'h6a;        memory[57894] <=  8'h67;        memory[57895] <=  8'h68;        memory[57896] <=  8'h66;        memory[57897] <=  8'h79;        memory[57898] <=  8'h74;        memory[57899] <=  8'h79;        memory[57900] <=  8'h69;        memory[57901] <=  8'h75;        memory[57902] <=  8'h64;        memory[57903] <=  8'h6a;        memory[57904] <=  8'h6b;        memory[57905] <=  8'h68;        memory[57906] <=  8'h63;        memory[57907] <=  8'h7a;        memory[57908] <=  8'h67;        memory[57909] <=  8'h68;        memory[57910] <=  8'h74;        memory[57911] <=  8'h75;        memory[57912] <=  8'h79;        memory[57913] <=  8'h69;        memory[57914] <=  8'h61;        memory[57915] <=  8'h73;        memory[57916] <=  8'h75;        memory[57917] <=  8'h6a;        memory[57918] <=  8'h6b;        memory[57919] <=  8'h62;        memory[57920] <=  8'h6e;        memory[57921] <=  8'h61;        memory[57922] <=  8'h76;        memory[57923] <=  8'h63;        memory[57924] <=  8'h66;        memory[57925] <=  8'h68;        memory[57926] <=  8'h75;        memory[57927] <=  8'h61;        memory[57928] <=  8'h73;        memory[57929] <=  8'h79;        memory[57930] <=  8'h64;        memory[57931] <=  8'h75;        memory[57932] <=  8'h69;        memory[57933] <=  8'h6a;        memory[57934] <=  8'h61;        memory[57935] <=  8'h6b;        memory[57936] <=  8'h62;        memory[57937] <=  8'h63;        memory[57938] <=  8'h78;        memory[57939] <=  8'h68;        memory[57940] <=  8'h67;        memory[57941] <=  8'h79;        memory[57942] <=  8'h75;        memory[57943] <=  8'h7a;        memory[57944] <=  8'h63;        memory[57945] <=  8'h61;        memory[57946] <=  8'h73;        memory[57947] <=  8'h69;        memory[57948] <=  8'h75;        memory[57949] <=  8'h6f;        memory[57950] <=  8'h69;        memory[57951] <=  8'h6a;        memory[57952] <=  8'h61;        memory[57953] <=  8'h6c;        memory[57954] <=  8'h63;        memory[57955] <=  8'h78;        memory[57956] <=  8'h62;        memory[57957] <=  8'h63;        memory[57958] <=  8'h20;        memory[57959] <=  8'h6e;        memory[57960] <=  8'h76;        memory[57961] <=  8'h63;        memory[57962] <=  8'h61;        memory[57963] <=  8'h64;        memory[57964] <=  8'h73;        memory[57965] <=  8'h67;        memory[57966] <=  8'h79;        memory[57967] <=  8'h68;        memory[57968] <=  8'h75;        memory[57969] <=  8'h61;        memory[57970] <=  8'h6a;        memory[57971] <=  8'h6b;        memory[57972] <=  8'h78;        memory[57973] <=  8'h62;        memory[57974] <=  8'h20;        memory[57975] <=  8'h6e;        memory[57976] <=  8'h76;        memory[57977] <=  8'h63;        memory[57978] <=  8'h61;        memory[57979] <=  8'h73;        memory[57980] <=  8'h67;        memory[57981] <=  8'h68;        memory[57982] <=  8'h75;        memory[57983] <=  8'h6a;        memory[57984] <=  8'h6c;        memory[57985] <=  8'h6b;        memory[57986] <=  8'h63;        memory[57987] <=  8'h78;        memory[57988] <=  8'h20;        memory[57989] <=  8'h6a;        memory[57990] <=  8'h6b;        memory[57991] <=  8'h68;        memory[57992] <=  8'h61;        memory[57993] <=  8'h73;        memory[57994] <=  8'h76;        memory[57995] <=  8'h64;        memory[57996] <=  8'h6e;        memory[57997] <=  8'h20;        memory[57998] <=  8'h62;        memory[57999] <=  8'h6e;        memory[58000] <=  8'h6d;        memory[58001] <=  8'h6b;        memory[58002] <=  8'h77;        memory[58003] <=  8'h64;        memory[58004] <=  8'h6f;        memory[58005] <=  8'h77;        memory[58006] <=  8'h69;        memory[58007] <=  8'h6f;        memory[58008] <=  8'h75;        memory[58009] <=  8'h69;        memory[58010] <=  8'h68;        memory[58011] <=  8'h62;        memory[58012] <=  8'h6e;        memory[58013] <=  8'h6b;        memory[58014] <=  8'h77;        memory[58015] <=  8'h69;        memory[58016] <=  8'h6f;        memory[58017] <=  8'h75;        memory[58018] <=  8'h71;        memory[58019] <=  8'h69;        memory[58020] <=  8'h79;        memory[58021] <=  8'h67;        memory[58022] <=  8'h6a;        memory[58023] <=  8'h64;        memory[58024] <=  8'h61;        memory[58025] <=  8'h76;        memory[58026] <=  8'h62;        memory[58027] <=  8'h6e;        memory[58028] <=  8'h6b;        memory[58029] <=  8'h6f;        memory[58030] <=  8'h70;        memory[58031] <=  8'h64;        memory[58032] <=  8'h76;        memory[58033] <=  8'h69;        memory[58034] <=  8'h6f;        memory[58035] <=  8'h75;        memory[58036] <=  8'h69;        memory[58037] <=  8'h48;        memory[58038] <=  8'h42;        memory[58039] <=  8'h6b;        memory[58040] <=  8'h64;        memory[58041] <=  8'h6e;        memory[58042] <=  8'h6c;        memory[58043] <=  8'h71;        memory[58044] <=  8'h6b;        memory[58045] <=  8'h6d;        memory[58046] <=  8'h6a;        memory[58047] <=  8'h70;        memory[58048] <=  8'h69;        memory[58049] <=  8'h6f;        memory[58050] <=  8'h68;        memory[58051] <=  8'h65;        memory[58052] <=  8'h66;        memory[58053] <=  8'h75;        memory[58054] <=  8'h67;        memory[58055] <=  8'h69;        memory[58056] <=  8'h73;        memory[58057] <=  8'h61;        memory[58058] <=  8'h62;        memory[58059] <=  8'h64;        memory[58060] <=  8'h6b;        memory[58061] <=  8'h6a;        memory[58062] <=  8'h6b;        memory[58063] <=  8'h6c;        memory[58064] <=  8'h6a;        memory[58065] <=  8'h69;        memory[58066] <=  8'h73;        memory[58067] <=  8'h6f;        memory[58068] <=  8'h71;        memory[58069] <=  8'h68;        memory[58070] <=  8'h77;        memory[58071] <=  8'h67;        memory[58072] <=  8'h69;        memory[58073] <=  8'h79;        memory[58074] <=  8'h6a;        memory[58075] <=  8'h64;        memory[58076] <=  8'h76;        memory[58077] <=  8'h62;        memory[58078] <=  8'h6e;        memory[58079] <=  8'h61;        memory[58080] <=  8'h73;        memory[58081] <=  8'h66;        memory[58082] <=  8'h6c;        memory[58083] <=  8'h6b;        memory[58084] <=  8'h64;        memory[58085] <=  8'h6a;        memory[58086] <=  8'h68;        memory[58087] <=  8'h63;        memory[58088] <=  8'h67;        memory[58089] <=  8'h6a;        memory[58090] <=  8'h76;        memory[58091] <=  8'h73;        memory[58092] <=  8'h64;        memory[58093] <=  8'h62;        memory[58094] <=  8'h62;        memory[58095] <=  8'h61;        memory[58096] <=  8'h72;        memory[58097] <=  8'h62;        memory[58098] <=  8'h62;        memory[58099] <=  8'h73;        memory[58100] <=  8'h62;        memory[58101] <=  8'h67;        memory[58102] <=  8'h73;        memory[58103] <=  8'h66;        memory[58104] <=  8'h67;        memory[58105] <=  8'h61;        memory[58106] <=  8'h68;        memory[58107] <=  8'h66;        memory[58108] <=  8'h73;        memory[58109] <=  8'h68;        memory[58110] <=  8'h61;        memory[58111] <=  8'h66;        memory[58112] <=  8'h73;        memory[58113] <=  8'h66;        memory[58114] <=  8'h68;        memory[58115] <=  8'h61;        memory[58116] <=  8'h69;        memory[58117] <=  8'h64;        memory[58118] <=  8'h75;        memory[58119] <=  8'h67;        memory[58120] <=  8'h64;        memory[58121] <=  8'h77;        memory[58122] <=  8'h62;        memory[58123] <=  8'h61;        memory[58124] <=  8'h62;        memory[58125] <=  8'h72;        memory[58126] <=  8'h62;        memory[58127] <=  8'h61;        memory[58128] <=  8'h62;        memory[58129] <=  8'h62;        memory[58130] <=  8'h74;        memory[58131] <=  8'h62;        memory[58132] <=  8'h62;        memory[58133] <=  8'h62;        memory[58134] <=  8'h62;        memory[58135] <=  8'h62;        memory[58136] <=  8'h62;        memory[58137] <=  8'h62;        memory[58138] <=  8'h62;        memory[58139] <=  8'h61;        memory[58140] <=  8'h62;        memory[58141] <=  8'h62;        memory[58142] <=  8'h72;        memory[58143] <=  8'h74;        memory[58144] <=  8'h62;        memory[58145] <=  8'h62;        memory[58146] <=  8'h61;        memory[58147] <=  8'h62;        memory[58148] <=  8'h72;        memory[58149] <=  8'h62;        memory[58150] <=  8'h74;        memory[58151] <=  8'h62;        memory[58152] <=  8'h62;        memory[58153] <=  8'h62;        memory[58154] <=  8'h63;        memory[58155] <=  8'h61;        memory[58156] <=  8'h72;        memory[58157] <=  8'h74;        memory[58158] <=  8'h73;        memory[58159] <=  8'h62;        memory[58160] <=  8'h61;        memory[58161] <=  8'h72;        memory[58162] <=  8'h74;        memory[58163] <=  8'h74;        memory[58164] <=  8'h62;        memory[58165] <=  8'h61;        memory[58166] <=  8'h72;        memory[58167] <=  8'h74;        memory[58168] <=  8'h78;        memory[58169] <=  8'h61;        memory[58170] <=  8'h74;        memory[58171] <=  8'h6b;        memory[58172] <=  8'h73;        memory[58173] <=  8'h68;        memory[58174] <=  8'h63;        memory[58175] <=  8'h66;        memory[58176] <=  8'h69;        memory[58177] <=  8'h77;        memory[58178] <=  8'h68;        memory[58179] <=  8'h61;        memory[58180] <=  8'h74;        memory[58181] <=  8'h61;        memory[58182] <=  8'h6e;        memory[58183] <=  8'h61;        memory[58184] <=  8'h62;        memory[58185] <=  8'h61;        memory[58186] <=  8'h63;        memory[58187] <=  8'h61;        memory[58188] <=  8'h74;        memory[58189] <=  8'h61;        memory[58190] <=  8'h62;        memory[58191] <=  8'h61;        memory[58192] <=  8'h72;        memory[58193] <=  8'h63;        memory[58194] <=  8'h61;        memory[58195] <=  8'h68;        memory[58196] <=  8'h64;        memory[58197] <=  8'h75;        memory[58198] <=  8'h63;        memory[58199] <=  8'h74;        memory[58200] <=  8'h61;        memory[58201] <=  8'h64;        memory[58202] <=  8'h61;        memory[58203] <=  8'h61;        memory[58204] <=  8'h63;        memory[58205] <=  8'h61;        memory[58206] <=  8'h72;        memory[58207] <=  8'h63;        memory[58208] <=  8'h74;        memory[58209] <=  8'h72;        memory[58210] <=  8'h63;        memory[58211] <=  8'h61;        memory[58212] <=  8'h74;        memory[58213] <=  8'h72;        memory[58214] <=  8'h63;        memory[58215] <=  8'h61;        memory[58216] <=  8'h74;        memory[58217] <=  8'h63;        memory[58218] <=  8'h62;        memory[58219] <=  8'h61;        memory[58220] <=  8'h74;        memory[58221] <=  8'h62;        memory[58222] <=  8'h72;        memory[58223] <=  8'h63;        memory[58224] <=  8'h61;        memory[58225] <=  8'h74;        memory[58226] <=  8'h72;        memory[58227] <=  8'h6e;        memory[58228] <=  8'h62;        memory[58229] <=  8'h61;        memory[58230] <=  8'h63;        memory[58231] <=  8'h61;        memory[58232] <=  8'h74;        memory[58233] <=  8'h79;        memory[58234] <=  8'h73;        memory[58235] <=  8'h6e;        memory[58236] <=  8'h63;        memory[58237] <=  8'h74;        memory[58238] <=  8'h61;        memory[58239] <=  8'h6e;        memory[58240] <=  8'h62;        memory[58241] <=  8'h61;        memory[58242] <=  8'h63;        memory[58243] <=  8'h72;        memory[58244] <=  8'h6e;        memory[58245] <=  8'h74;        memory[58246] <=  8'h61;        memory[58247] <=  8'h62;        memory[58248] <=  8'h74;        memory[58249] <=  8'h6e;        memory[58250] <=  8'h61;        memory[58251] <=  8'h72;        memory[58252] <=  8'h62;        memory[58253] <=  8'h78;        memory[58254] <=  8'h74;        memory[58255] <=  8'h61;        memory[58256] <=  8'h72;        memory[58257] <=  8'h62;        memory[58258] <=  8'h61;        memory[58259] <=  8'h72;        memory[58260] <=  8'h74;        memory[58261] <=  8'h74;        memory[58262] <=  8'h62;        memory[58263] <=  8'h61;        memory[58264] <=  8'h72;        memory[58265] <=  8'h74;        memory[58266] <=  8'h78;        memory[58267] <=  8'h61;        memory[58268] <=  8'h74;        memory[58269] <=  8'h6b;        memory[58270] <=  8'h73;        memory[58271] <=  8'h68;        memory[58272] <=  8'h63;        memory[58273] <=  8'h66;        memory[58274] <=  8'h69;        memory[58275] <=  8'h77;        memory[58276] <=  8'h68;        memory[58277] <=  8'h61;        memory[58278] <=  8'h74;        memory[58279] <=  8'h61;        memory[58280] <=  8'h6e;        memory[58281] <=  8'h61;        memory[58282] <=  8'h62;        memory[58283] <=  8'h61;        memory[58284] <=  8'h63;        memory[58285] <=  8'h61;        memory[58286] <=  8'h74;        memory[58287] <=  8'h61;        memory[58288] <=  8'h62;        memory[58289] <=  8'h61;        memory[58290] <=  8'h72;        memory[58291] <=  8'h63;        memory[58292] <=  8'h61;        memory[58293] <=  8'h68;        memory[58294] <=  8'h64;        memory[58295] <=  8'h75;        memory[58296] <=  8'h63;        memory[58297] <=  8'h74;        memory[58298] <=  8'h61;        memory[58299] <=  8'h64;        memory[58300] <=  8'h61;        memory[58301] <=  8'h61;        memory[58302] <=  8'h63;        memory[58303] <=  8'h61;        memory[58304] <=  8'h72;        memory[58305] <=  8'h63;        memory[58306] <=  8'h74;        memory[58307] <=  8'h72;        memory[58308] <=  8'h63;        memory[58309] <=  8'h61;        memory[58310] <=  8'h74;        memory[58311] <=  8'h72;        memory[58312] <=  8'h63;        memory[58313] <=  8'h61;        memory[58314] <=  8'h74;        memory[58315] <=  8'h63;        memory[58316] <=  8'h62;        memory[58317] <=  8'h61;        memory[58318] <=  8'h74;        memory[58319] <=  8'h62;        memory[58320] <=  8'h72;        memory[58321] <=  8'h63;        memory[58322] <=  8'h61;        memory[58323] <=  8'h74;        memory[58324] <=  8'h72;        memory[58325] <=  8'h6e;        memory[58326] <=  8'h62;        memory[58327] <=  8'h61;        memory[58328] <=  8'h63;        memory[58329] <=  8'h61;        memory[58330] <=  8'h74;        memory[58331] <=  8'h79;        memory[58332] <=  8'h73;        memory[58333] <=  8'h6e;        memory[58334] <=  8'h63;        memory[58335] <=  8'h74;        memory[58336] <=  8'h61;        memory[58337] <=  8'h6e;        memory[58338] <=  8'h62;        memory[58339] <=  8'h61;        memory[58340] <=  8'h63;        memory[58341] <=  8'h72;        memory[58342] <=  8'h6e;        memory[58343] <=  8'h74;        memory[58344] <=  8'h61;        memory[58345] <=  8'h62;        memory[58346] <=  8'h74;        memory[58347] <=  8'h6e;        memory[58348] <=  8'h61;        memory[58349] <=  8'h72;        memory[58350] <=  8'h62;        memory[58351] <=  8'h78;        memory[58352] <=  8'h74;        memory[58353] <=  8'h61;        memory[58354] <=  8'h72;        memory[58355] <=  8'h62;        memory[58356] <=  8'h61;        memory[58357] <=  8'h72;        memory[58358] <=  8'h74;        memory[58359] <=  8'h74;        memory[58360] <=  8'h62;        memory[58361] <=  8'h61;        memory[58362] <=  8'h72;        memory[58363] <=  8'h74;        memory[58364] <=  8'h78;        memory[58365] <=  8'h61;        memory[58366] <=  8'h74;        memory[58367] <=  8'h6b;        memory[58368] <=  8'h73;        memory[58369] <=  8'h68;        memory[58370] <=  8'h63;        memory[58371] <=  8'h66;        memory[58372] <=  8'h69;        memory[58373] <=  8'h77;        memory[58374] <=  8'h68;        memory[58375] <=  8'h61;        memory[58376] <=  8'h74;        memory[58377] <=  8'h61;        memory[58378] <=  8'h6e;        memory[58379] <=  8'h61;        memory[58380] <=  8'h62;        memory[58381] <=  8'h61;        memory[58382] <=  8'h63;        memory[58383] <=  8'h61;        memory[58384] <=  8'h74;        memory[58385] <=  8'h61;        memory[58386] <=  8'h62;        memory[58387] <=  8'h61;        memory[58388] <=  8'h72;        memory[58389] <=  8'h63;        memory[58390] <=  8'h61;        memory[58391] <=  8'h68;        memory[58392] <=  8'h64;        memory[58393] <=  8'h75;        memory[58394] <=  8'h63;        memory[58395] <=  8'h74;        memory[58396] <=  8'h61;        memory[58397] <=  8'h64;        memory[58398] <=  8'h61;        memory[58399] <=  8'h61;        memory[58400] <=  8'h63;        memory[58401] <=  8'h61;        memory[58402] <=  8'h72;        memory[58403] <=  8'h63;        memory[58404] <=  8'h74;        memory[58405] <=  8'h72;        memory[58406] <=  8'h63;        memory[58407] <=  8'h61;        memory[58408] <=  8'h74;        memory[58409] <=  8'h72;        memory[58410] <=  8'h63;        memory[58411] <=  8'h61;        memory[58412] <=  8'h74;        memory[58413] <=  8'h63;        memory[58414] <=  8'h62;        memory[58415] <=  8'h61;        memory[58416] <=  8'h74;        memory[58417] <=  8'h62;        memory[58418] <=  8'h72;        memory[58419] <=  8'h63;        memory[58420] <=  8'h61;        memory[58421] <=  8'h74;        memory[58422] <=  8'h72;        memory[58423] <=  8'h6e;        memory[58424] <=  8'h62;        memory[58425] <=  8'h61;        memory[58426] <=  8'h63;        memory[58427] <=  8'h61;        memory[58428] <=  8'h74;        memory[58429] <=  8'h79;        memory[58430] <=  8'h73;        memory[58431] <=  8'h6e;        memory[58432] <=  8'h63;        memory[58433] <=  8'h74;        memory[58434] <=  8'h61;        memory[58435] <=  8'h6e;        memory[58436] <=  8'h62;        memory[58437] <=  8'h61;        memory[58438] <=  8'h63;        memory[58439] <=  8'h72;        memory[58440] <=  8'h6e;        memory[58441] <=  8'h74;        memory[58442] <=  8'h61;        memory[58443] <=  8'h62;        memory[58444] <=  8'h74;        memory[58445] <=  8'h6e;        memory[58446] <=  8'h61;        memory[58447] <=  8'h72;        memory[58448] <=  8'h62;        memory[58449] <=  8'h78;        memory[58450] <=  8'h74;        memory[58451] <=  8'h61;        memory[58452] <=  8'h72;        memory[58453] <=  8'h5d;        memory[58454] <=  8'h5d;        memory[58455] <=  8'h65;        memory[58456] <=  8'h66;        memory[58457] <=  8'h77;        memory[58458] <=  8'h65;        memory[58459] <=  8'h5d;        memory[58460] <=  8'h65;        memory[58461] <=  8'h67;        memory[58462] <=  8'h73;        memory[58463] <=  8'h67;        memory[58464] <=  8'h66;        memory[58465] <=  8'h62;        memory[58466] <=  8'h61;        memory[58467] <=  8'h72;        memory[58468] <=  8'h74;        memory[58469] <=  8'h74;        memory[58470] <=  8'h62;        memory[58471] <=  8'h61;        memory[58472] <=  8'h72;        memory[58473] <=  8'h74;        memory[58474] <=  8'h78;        memory[58475] <=  8'h61;        memory[58476] <=  8'h74;        memory[58477] <=  8'h6b;        memory[58478] <=  8'h73;        memory[58479] <=  8'h68;        memory[58480] <=  8'h63;        memory[58481] <=  8'h66;        memory[58482] <=  8'h69;        memory[58483] <=  8'h77;        memory[58484] <=  8'h68;        memory[58485] <=  8'h61;        memory[58486] <=  8'h74;        memory[58487] <=  8'h61;        memory[58488] <=  8'h6e;        memory[58489] <=  8'h61;        memory[58490] <=  8'h62;        memory[58491] <=  8'h61;        memory[58492] <=  8'h63;        memory[58493] <=  8'h61;        memory[58494] <=  8'h74;        memory[58495] <=  8'h61;        memory[58496] <=  8'h62;        memory[58497] <=  8'h61;        memory[58498] <=  8'h72;        memory[58499] <=  8'h63;        memory[58500] <=  8'h61;        memory[58501] <=  8'h68;        memory[58502] <=  8'h64;        memory[58503] <=  8'h75;        memory[58504] <=  8'h63;        memory[58505] <=  8'h74;        memory[58506] <=  8'h61;        memory[58507] <=  8'h64;        memory[58508] <=  8'h61;        memory[58509] <=  8'h61;        memory[58510] <=  8'h63;        memory[58511] <=  8'h61;        memory[58512] <=  8'h72;        memory[58513] <=  8'h63;        memory[58514] <=  8'h74;        memory[58515] <=  8'h72;        memory[58516] <=  8'h63;        memory[58517] <=  8'h61;        memory[58518] <=  8'h74;        memory[58519] <=  8'h72;        memory[58520] <=  8'h63;        memory[58521] <=  8'h61;        memory[58522] <=  8'h74;        memory[58523] <=  8'h63;        memory[58524] <=  8'h62;        memory[58525] <=  8'h61;        memory[58526] <=  8'h74;        memory[58527] <=  8'h62;        memory[58528] <=  8'h72;        memory[58529] <=  8'h63;        memory[58530] <=  8'h61;        memory[58531] <=  8'h74;        memory[58532] <=  8'h72;        memory[58533] <=  8'h6e;        memory[58534] <=  8'h62;        memory[58535] <=  8'h61;        memory[58536] <=  8'h63;        memory[58537] <=  8'h61;        memory[58538] <=  8'h74;        memory[58539] <=  8'h79;        memory[58540] <=  8'h73;        memory[58541] <=  8'h6e;        memory[58542] <=  8'h63;        memory[58543] <=  8'h74;        memory[58544] <=  8'h61;        memory[58545] <=  8'h6e;        memory[58546] <=  8'h62;        memory[58547] <=  8'h61;        memory[58548] <=  8'h63;        memory[58549] <=  8'h72;        memory[58550] <=  8'h6e;        memory[58551] <=  8'h74;        memory[58552] <=  8'h61;        memory[58553] <=  8'h62;        memory[58554] <=  8'h74;        memory[58555] <=  8'h6e;        memory[58556] <=  8'h61;        memory[58557] <=  8'h72;        memory[58558] <=  8'h62;        memory[58559] <=  8'h78;        memory[58560] <=  8'h74;        memory[58561] <=  8'h61;        memory[58562] <=  8'h72;        memory[58563] <=  8'h62;        memory[58564] <=  8'h61;        memory[58565] <=  8'h72;        memory[58566] <=  8'h74;        memory[58567] <=  8'h74;        memory[58568] <=  8'h62;        memory[58569] <=  8'h61;        memory[58570] <=  8'h72;        memory[58571] <=  8'h74;        memory[58572] <=  8'h78;        memory[58573] <=  8'h61;        memory[58574] <=  8'h74;        memory[58575] <=  8'h6b;        memory[58576] <=  8'h73;        memory[58577] <=  8'h68;        memory[58578] <=  8'h63;        memory[58579] <=  8'h66;        memory[58580] <=  8'h69;        memory[58581] <=  8'h77;        memory[58582] <=  8'h68;        memory[58583] <=  8'h61;        memory[58584] <=  8'h74;        memory[58585] <=  8'h61;        memory[58586] <=  8'h6e;        memory[58587] <=  8'h61;        memory[58588] <=  8'h62;        memory[58589] <=  8'h61;        memory[58590] <=  8'h63;        memory[58591] <=  8'h61;        memory[58592] <=  8'h74;        memory[58593] <=  8'h61;        memory[58594] <=  8'h62;        memory[58595] <=  8'h61;        memory[58596] <=  8'h72;        memory[58597] <=  8'h63;        memory[58598] <=  8'h61;        memory[58599] <=  8'h68;        memory[58600] <=  8'h64;        memory[58601] <=  8'h75;        memory[58602] <=  8'h63;        memory[58603] <=  8'h74;        memory[58604] <=  8'h61;        memory[58605] <=  8'h64;        memory[58606] <=  8'h61;        memory[58607] <=  8'h61;        memory[58608] <=  8'h63;        memory[58609] <=  8'h61;        memory[58610] <=  8'h72;        memory[58611] <=  8'h63;        memory[58612] <=  8'h74;        memory[58613] <=  8'h72;        memory[58614] <=  8'h63;        memory[58615] <=  8'h61;        memory[58616] <=  8'h74;        memory[58617] <=  8'h72;        memory[58618] <=  8'h63;        memory[58619] <=  8'h61;        memory[58620] <=  8'h74;        memory[58621] <=  8'h63;        memory[58622] <=  8'h62;        memory[58623] <=  8'h61;        memory[58624] <=  8'h74;        memory[58625] <=  8'h62;        memory[58626] <=  8'h72;        memory[58627] <=  8'h63;        memory[58628] <=  8'h61;        memory[58629] <=  8'h74;        memory[58630] <=  8'h72;        memory[58631] <=  8'h6e;        memory[58632] <=  8'h62;        memory[58633] <=  8'h61;        memory[58634] <=  8'h63;        memory[58635] <=  8'h61;        memory[58636] <=  8'h74;        memory[58637] <=  8'h79;        memory[58638] <=  8'h73;        memory[58639] <=  8'h6e;        memory[58640] <=  8'h63;        memory[58641] <=  8'h74;        memory[58642] <=  8'h61;        memory[58643] <=  8'h6e;        memory[58644] <=  8'h62;        memory[58645] <=  8'h61;        memory[58646] <=  8'h63;        memory[58647] <=  8'h72;        memory[58648] <=  8'h6e;        memory[58649] <=  8'h74;        memory[58650] <=  8'h61;        memory[58651] <=  8'h62;        memory[58652] <=  8'h74;        memory[58653] <=  8'h6e;        memory[58654] <=  8'h61;        memory[58655] <=  8'h72;        memory[58656] <=  8'h62;        memory[58657] <=  8'h78;        memory[58658] <=  8'h74;        memory[58659] <=  8'h61;        memory[58660] <=  8'h72;        memory[58661] <=  8'h64;        memory[58662] <=  8'h66;        memory[58663] <=  8'h73;        memory[58664] <=  8'h67;        memory[58665] <=  8'h76;        memory[58666] <=  8'h68;        memory[58667] <=  8'h62;        memory[58668] <=  8'h6b;        memory[58669] <=  8'h6a;        memory[58670] <=  8'h6e;        memory[58671] <=  8'h6d;        memory[58672] <=  8'h62;        memory[58673] <=  8'h76;        memory[58674] <=  8'h78;        memory[58675] <=  8'h63;        memory[58676] <=  8'h73;        memory[58677] <=  8'h66;        memory[58678] <=  8'h72;        memory[58679] <=  8'h74;        memory[58680] <=  8'h79;        memory[58681] <=  8'h75;        memory[58682] <=  8'h6a;        memory[58683] <=  8'h6e;        memory[58684] <=  8'h62;        memory[58685] <=  8'h76;        memory[58686] <=  8'h63;        memory[58687] <=  8'h64;        memory[58688] <=  8'h74;        memory[58689] <=  8'h79;        memory[58690] <=  8'h75;        memory[58691] <=  8'h69;        memory[58692] <=  8'h6b;        memory[58693] <=  8'h6d;        memory[58694] <=  8'h6e;        memory[58695] <=  8'h62;        memory[58696] <=  8'h76;        memory[58697] <=  8'h63;        memory[58698] <=  8'h78;        memory[58699] <=  8'h73;        memory[58700] <=  8'h64;        memory[58701] <=  8'h72;        memory[58702] <=  8'h74;        memory[58703] <=  8'h79;        memory[58704] <=  8'h75;        memory[58705] <=  8'h69;        memory[58706] <=  8'h6b;        memory[58707] <=  8'h6d;        memory[58708] <=  8'h6e;        memory[58709] <=  8'h62;        memory[58710] <=  8'h76;        memory[58711] <=  8'h63;        memory[58712] <=  8'h73;        memory[58713] <=  8'h77;        memory[58714] <=  8'h33;        memory[58715] <=  8'h34;        memory[58716] <=  8'h35;        memory[58717] <=  8'h36;        memory[58718] <=  8'h37;        memory[58719] <=  8'h38;        memory[58720] <=  8'h69;        memory[58721] <=  8'h6b;        memory[58722] <=  8'h6d;        memory[58723] <=  8'h6e;        memory[58724] <=  8'h62;        memory[58725] <=  8'h76;        memory[58726] <=  8'h63;        memory[58727] <=  8'h64;        memory[58728] <=  8'h65;        memory[58729] <=  8'h72;        memory[58730] <=  8'h36;        memory[58731] <=  8'h37;        memory[58732] <=  8'h38;        memory[58733] <=  8'h69;        memory[58734] <=  8'h6f;        memory[58735] <=  8'h6b;        memory[58736] <=  8'h6a;        memory[58737] <=  8'h6e;        memory[58738] <=  8'h62;        memory[58739] <=  8'h76;        memory[58740] <=  8'h63;        memory[58741] <=  8'h64;        memory[58742] <=  8'h72;        memory[58743] <=  8'h74;        memory[58744] <=  8'h79;        memory[58745] <=  8'h75;        memory[58746] <=  8'h73;        memory[58747] <=  8'h6a;        memory[58748] <=  8'h63;        memory[58749] <=  8'h6e;        memory[58750] <=  8'h62;        memory[58751] <=  8'h64;        memory[58752] <=  8'h66;        memory[58753] <=  8'h73;        memory[58754] <=  8'h74;        memory[58755] <=  8'h79;        memory[58756] <=  8'h75;        memory[58757] <=  8'h61;        memory[58758] <=  8'h69;        memory[58759] <=  8'h6b;        memory[58760] <=  8'h78;        memory[58761] <=  8'h6d;        memory[58762] <=  8'h6e;        memory[58763] <=  8'h73;        memory[58764] <=  8'h6a;        memory[58765] <=  8'h6f;        memory[58766] <=  8'h64;        memory[58767] <=  8'h6c;        memory[58768] <=  8'h63;        memory[58769] <=  8'h78;        memory[58770] <=  8'h62;        memory[58771] <=  8'h61;        memory[58772] <=  8'h72;        memory[58773] <=  8'h74;        memory[58774] <=  8'h78;        memory[58775] <=  8'h61;        memory[58776] <=  8'h74;        memory[58777] <=  8'h6b;        memory[58778] <=  8'h73;        memory[58779] <=  8'h68;        memory[58780] <=  8'h63;        memory[58781] <=  8'h66;        memory[58782] <=  8'h69;        memory[58783] <=  8'h77;        memory[58784] <=  8'h68;        memory[58785] <=  8'h61;        memory[58786] <=  8'h74;        memory[58787] <=  8'h61;        memory[58788] <=  8'h6e;        memory[58789] <=  8'h61;        memory[58790] <=  8'h62;        memory[58791] <=  8'h61;        memory[58792] <=  8'h63;        memory[58793] <=  8'h61;        memory[58794] <=  8'h74;        memory[58795] <=  8'h61;        memory[58796] <=  8'h62;        memory[58797] <=  8'h61;        memory[58798] <=  8'h72;        memory[58799] <=  8'h63;        memory[58800] <=  8'h61;        memory[58801] <=  8'h68;        memory[58802] <=  8'h64;        memory[58803] <=  8'h75;        memory[58804] <=  8'h63;        memory[58805] <=  8'h74;        memory[58806] <=  8'h61;        memory[58807] <=  8'h64;        memory[58808] <=  8'h61;        memory[58809] <=  8'h61;        memory[58810] <=  8'h63;        memory[58811] <=  8'h61;        memory[58812] <=  8'h72;        memory[58813] <=  8'h62;        memory[58814] <=  8'h61;        memory[58815] <=  8'h72;        memory[58816] <=  8'h74;        memory[58817] <=  8'h78;        memory[58818] <=  8'h61;        memory[58819] <=  8'h74;        memory[58820] <=  8'h6b;        memory[58821] <=  8'h73;        memory[58822] <=  8'h68;        memory[58823] <=  8'h63;        memory[58824] <=  8'h66;        memory[58825] <=  8'h69;        memory[58826] <=  8'h77;        memory[58827] <=  8'h68;        memory[58828] <=  8'h61;        memory[58829] <=  8'h74;        memory[58830] <=  8'h61;        memory[58831] <=  8'h6e;        memory[58832] <=  8'h61;        memory[58833] <=  8'h62;        memory[58834] <=  8'h61;        memory[58835] <=  8'h63;        memory[58836] <=  8'h61;        memory[58837] <=  8'h74;        memory[58838] <=  8'h61;        memory[58839] <=  8'h62;        memory[58840] <=  8'h61;        memory[58841] <=  8'h72;        memory[58842] <=  8'h63;        memory[58843] <=  8'h61;        memory[58844] <=  8'h68;        memory[58845] <=  8'h64;        memory[58846] <=  8'h75;        memory[58847] <=  8'h63;        memory[58848] <=  8'h74;        memory[58849] <=  8'h61;        memory[58850] <=  8'h64;        memory[58851] <=  8'h61;        memory[58852] <=  8'h61;        memory[58853] <=  8'h63;        memory[58854] <=  8'h61;        memory[58855] <=  8'h72;        memory[58856] <=  8'h62;        memory[58857] <=  8'h61;        memory[58858] <=  8'h72;        memory[58859] <=  8'h74;        memory[58860] <=  8'h78;        memory[58861] <=  8'h61;        memory[58862] <=  8'h74;        memory[58863] <=  8'h6b;        memory[58864] <=  8'h73;        memory[58865] <=  8'h68;        memory[58866] <=  8'h63;        memory[58867] <=  8'h66;        memory[58868] <=  8'h69;        memory[58869] <=  8'h77;        memory[58870] <=  8'h68;        memory[58871] <=  8'h61;        memory[58872] <=  8'h74;        memory[58873] <=  8'h61;        memory[58874] <=  8'h6e;        memory[58875] <=  8'h61;        memory[58876] <=  8'h62;        memory[58877] <=  8'h61;        memory[58878] <=  8'h63;        memory[58879] <=  8'h61;        memory[58880] <=  8'h74;        memory[58881] <=  8'h61;        memory[58882] <=  8'h62;        memory[58883] <=  8'h61;        memory[58884] <=  8'h72;        memory[58885] <=  8'h63;        memory[58886] <=  8'h61;        memory[58887] <=  8'h68;        memory[58888] <=  8'h64;        memory[58889] <=  8'h75;        memory[58890] <=  8'h63;        memory[58891] <=  8'h74;        memory[58892] <=  8'h61;        memory[58893] <=  8'h64;        memory[58894] <=  8'h61;        memory[58895] <=  8'h61;        memory[58896] <=  8'h63;        memory[58897] <=  8'h61;        memory[58898] <=  8'h72;        memory[58899] <=  8'h62;        memory[58900] <=  8'h61;        memory[58901] <=  8'h72;        memory[58902] <=  8'h74;        memory[58903] <=  8'h78;        memory[58904] <=  8'h61;        memory[58905] <=  8'h74;        memory[58906] <=  8'h6b;        memory[58907] <=  8'h73;        memory[58908] <=  8'h68;        memory[58909] <=  8'h63;        memory[58910] <=  8'h66;        memory[58911] <=  8'h69;        memory[58912] <=  8'h77;        memory[58913] <=  8'h68;        memory[58914] <=  8'h61;        memory[58915] <=  8'h74;        memory[58916] <=  8'h61;        memory[58917] <=  8'h6e;        memory[58918] <=  8'h61;        memory[58919] <=  8'h62;        memory[58920] <=  8'h61;        memory[58921] <=  8'h63;        memory[58922] <=  8'h61;        memory[58923] <=  8'h74;        memory[58924] <=  8'h61;        memory[58925] <=  8'h62;        memory[58926] <=  8'h61;        memory[58927] <=  8'h72;        memory[58928] <=  8'h63;        memory[58929] <=  8'h61;        memory[58930] <=  8'h68;        memory[58931] <=  8'h64;        memory[58932] <=  8'h75;        memory[58933] <=  8'h63;        memory[58934] <=  8'h74;        memory[58935] <=  8'h61;        memory[58936] <=  8'h64;        memory[58937] <=  8'h61;        memory[58938] <=  8'h61;        memory[58939] <=  8'h63;        memory[58940] <=  8'h61;        memory[58941] <=  8'h72;        memory[58942] <=  8'h62;        memory[58943] <=  8'h61;        memory[58944] <=  8'h72;        memory[58945] <=  8'h74;        memory[58946] <=  8'h78;        memory[58947] <=  8'h61;        memory[58948] <=  8'h74;        memory[58949] <=  8'h6b;        memory[58950] <=  8'h73;        memory[58951] <=  8'h68;        memory[58952] <=  8'h63;        memory[58953] <=  8'h66;        memory[58954] <=  8'h69;        memory[58955] <=  8'h77;        memory[58956] <=  8'h68;        memory[58957] <=  8'h61;        memory[58958] <=  8'h74;        memory[58959] <=  8'h61;        memory[58960] <=  8'h6e;        memory[58961] <=  8'h61;        memory[58962] <=  8'h62;        memory[58963] <=  8'h61;        memory[58964] <=  8'h63;        memory[58965] <=  8'h61;        memory[58966] <=  8'h74;        memory[58967] <=  8'h61;        memory[58968] <=  8'h62;        memory[58969] <=  8'h61;        memory[58970] <=  8'h72;        memory[58971] <=  8'h63;        memory[58972] <=  8'h61;        memory[58973] <=  8'h68;        memory[58974] <=  8'h64;        memory[58975] <=  8'h75;        memory[58976] <=  8'h63;        memory[58977] <=  8'h74;        memory[58978] <=  8'h61;        memory[58979] <=  8'h64;        memory[58980] <=  8'h61;        memory[58981] <=  8'h61;        memory[58982] <=  8'h63;        memory[58983] <=  8'h61;        memory[58984] <=  8'h72;        memory[58985] <=  8'h62;        memory[58986] <=  8'h61;        memory[58987] <=  8'h72;        memory[58988] <=  8'h74;        memory[58989] <=  8'h78;        memory[58990] <=  8'h61;        memory[58991] <=  8'h74;        memory[58992] <=  8'h6b;        memory[58993] <=  8'h73;        memory[58994] <=  8'h68;        memory[58995] <=  8'h63;        memory[58996] <=  8'h66;        memory[58997] <=  8'h69;        memory[58998] <=  8'h77;        memory[58999] <=  8'h68;        memory[59000] <=  8'h61;        memory[59001] <=  8'h74;        memory[59002] <=  8'h61;        memory[59003] <=  8'h6e;        memory[59004] <=  8'h61;        memory[59005] <=  8'h62;        memory[59006] <=  8'h61;        memory[59007] <=  8'h63;        memory[59008] <=  8'h61;        memory[59009] <=  8'h74;        memory[59010] <=  8'h61;        memory[59011] <=  8'h62;        memory[59012] <=  8'h61;        memory[59013] <=  8'h72;        memory[59014] <=  8'h63;        memory[59015] <=  8'h61;        memory[59016] <=  8'h68;        memory[59017] <=  8'h64;        memory[59018] <=  8'h75;        memory[59019] <=  8'h63;        memory[59020] <=  8'h74;        memory[59021] <=  8'h61;        memory[59022] <=  8'h64;        memory[59023] <=  8'h61;        memory[59024] <=  8'h61;        memory[59025] <=  8'h63;        memory[59026] <=  8'h61;        memory[59027] <=  8'h72;        memory[59028] <=  8'h62;        memory[59029] <=  8'h61;        memory[59030] <=  8'h72;        memory[59031] <=  8'h74;        memory[59032] <=  8'h78;        memory[59033] <=  8'h61;        memory[59034] <=  8'h74;        memory[59035] <=  8'h6b;        memory[59036] <=  8'h73;        memory[59037] <=  8'h68;        memory[59038] <=  8'h63;        memory[59039] <=  8'h66;        memory[59040] <=  8'h69;        memory[59041] <=  8'h77;        memory[59042] <=  8'h68;        memory[59043] <=  8'h61;        memory[59044] <=  8'h74;        memory[59045] <=  8'h61;        memory[59046] <=  8'h6e;        memory[59047] <=  8'h61;        memory[59048] <=  8'h62;        memory[59049] <=  8'h61;        memory[59050] <=  8'h63;        memory[59051] <=  8'h61;        memory[59052] <=  8'h74;        memory[59053] <=  8'h61;        memory[59054] <=  8'h62;        memory[59055] <=  8'h61;        memory[59056] <=  8'h72;        memory[59057] <=  8'h63;        memory[59058] <=  8'h61;        memory[59059] <=  8'h68;        memory[59060] <=  8'h64;        memory[59061] <=  8'h75;        memory[59062] <=  8'h63;        memory[59063] <=  8'h74;        memory[59064] <=  8'h61;        memory[59065] <=  8'h64;        memory[59066] <=  8'h61;        memory[59067] <=  8'h61;        memory[59068] <=  8'h63;        memory[59069] <=  8'h61;        memory[59070] <=  8'h72;        memory[59071] <=  8'h62;        memory[59072] <=  8'h61;        memory[59073] <=  8'h72;        memory[59074] <=  8'h74;        memory[59075] <=  8'h78;        memory[59076] <=  8'h61;        memory[59077] <=  8'h74;        memory[59078] <=  8'h6b;        memory[59079] <=  8'h73;        memory[59080] <=  8'h68;        memory[59081] <=  8'h63;        memory[59082] <=  8'h66;        memory[59083] <=  8'h69;        memory[59084] <=  8'h77;        memory[59085] <=  8'h68;        memory[59086] <=  8'h61;        memory[59087] <=  8'h74;        memory[59088] <=  8'h61;        memory[59089] <=  8'h6e;        memory[59090] <=  8'h61;        memory[59091] <=  8'h62;        memory[59092] <=  8'h61;        memory[59093] <=  8'h63;        memory[59094] <=  8'h61;        memory[59095] <=  8'h74;        memory[59096] <=  8'h61;        memory[59097] <=  8'h62;        memory[59098] <=  8'h61;        memory[59099] <=  8'h72;        memory[59100] <=  8'h63;        memory[59101] <=  8'h61;        memory[59102] <=  8'h68;        memory[59103] <=  8'h64;        memory[59104] <=  8'h75;        memory[59105] <=  8'h63;        memory[59106] <=  8'h74;        memory[59107] <=  8'h61;        memory[59108] <=  8'h64;        memory[59109] <=  8'h61;        memory[59110] <=  8'h61;        memory[59111] <=  8'h63;        memory[59112] <=  8'h61;        memory[59113] <=  8'h72;        memory[59114] <=  8'h62;        memory[59115] <=  8'h61;        memory[59116] <=  8'h72;        memory[59117] <=  8'h74;        memory[59118] <=  8'h78;        memory[59119] <=  8'h61;        memory[59120] <=  8'h74;        memory[59121] <=  8'h6b;        memory[59122] <=  8'h73;        memory[59123] <=  8'h68;        memory[59124] <=  8'h63;        memory[59125] <=  8'h66;        memory[59126] <=  8'h69;        memory[59127] <=  8'h77;        memory[59128] <=  8'h68;        memory[59129] <=  8'h61;        memory[59130] <=  8'h74;        memory[59131] <=  8'h61;        memory[59132] <=  8'h6e;        memory[59133] <=  8'h61;        memory[59134] <=  8'h62;        memory[59135] <=  8'h61;        memory[59136] <=  8'h63;        memory[59137] <=  8'h61;        memory[59138] <=  8'h74;        memory[59139] <=  8'h61;        memory[59140] <=  8'h62;        memory[59141] <=  8'h61;        memory[59142] <=  8'h72;        memory[59143] <=  8'h63;        memory[59144] <=  8'h61;        memory[59145] <=  8'h68;        memory[59146] <=  8'h64;        memory[59147] <=  8'h75;        memory[59148] <=  8'h63;        memory[59149] <=  8'h74;        memory[59150] <=  8'h61;        memory[59151] <=  8'h64;        memory[59152] <=  8'h61;        memory[59153] <=  8'h61;        memory[59154] <=  8'h63;        memory[59155] <=  8'h61;        memory[59156] <=  8'h72;        memory[59157] <=  8'h62;        memory[59158] <=  8'h61;        memory[59159] <=  8'h72;        memory[59160] <=  8'h74;        memory[59161] <=  8'h74;        memory[59162] <=  8'h62;        memory[59163] <=  8'h61;        memory[59164] <=  8'h72;        memory[59165] <=  8'h74;        memory[59166] <=  8'h78;        memory[59167] <=  8'h61;        memory[59168] <=  8'h74;        memory[59169] <=  8'h6b;        memory[59170] <=  8'h73;        memory[59171] <=  8'h68;        memory[59172] <=  8'h63;        memory[59173] <=  8'h66;        memory[59174] <=  8'h69;        memory[59175] <=  8'h77;        memory[59176] <=  8'h68;        memory[59177] <=  8'h61;        memory[59178] <=  8'h74;        memory[59179] <=  8'h61;        memory[59180] <=  8'h6e;        memory[59181] <=  8'h61;        memory[59182] <=  8'h62;        memory[59183] <=  8'h61;        memory[59184] <=  8'h63;        memory[59185] <=  8'h61;        memory[59186] <=  8'h74;        memory[59187] <=  8'h61;        memory[59188] <=  8'h62;        memory[59189] <=  8'h61;        memory[59190] <=  8'h72;        memory[59191] <=  8'h63;        memory[59192] <=  8'h61;        memory[59193] <=  8'h68;        memory[59194] <=  8'h64;        memory[59195] <=  8'h75;        memory[59196] <=  8'h63;        memory[59197] <=  8'h74;        memory[59198] <=  8'h61;        memory[59199] <=  8'h64;        memory[59200] <=  8'h61;        memory[59201] <=  8'h61;        memory[59202] <=  8'h63;        memory[59203] <=  8'h61;        memory[59204] <=  8'h72;        memory[59205] <=  8'h63;        memory[59206] <=  8'h74;        memory[59207] <=  8'h72;        memory[59208] <=  8'h63;        memory[59209] <=  8'h61;        memory[59210] <=  8'h74;        memory[59211] <=  8'h72;        memory[59212] <=  8'h63;        memory[59213] <=  8'h61;        memory[59214] <=  8'h74;        memory[59215] <=  8'h63;        memory[59216] <=  8'h62;        memory[59217] <=  8'h61;        memory[59218] <=  8'h74;        memory[59219] <=  8'h62;        memory[59220] <=  8'h72;        memory[59221] <=  8'h63;        memory[59222] <=  8'h61;        memory[59223] <=  8'h72;        memory[59224] <=  8'h62;        memory[59225] <=  8'h78;        memory[59226] <=  8'h74;        memory[59227] <=  8'h61;        memory[59228] <=  8'h72;        memory[59229] <=  8'h64;        memory[59230] <=  8'h66;        memory[59231] <=  8'h73;        memory[59232] <=  8'h67;        memory[59233] <=  8'h76;        memory[59234] <=  8'h68;        memory[59235] <=  8'h62;        memory[59236] <=  8'h6b;        memory[59237] <=  8'h6a;        memory[59238] <=  8'h6e;        memory[59239] <=  8'h6d;        memory[59240] <=  8'h62;        memory[59241] <=  8'h76;        memory[59242] <=  8'h78;        memory[59243] <=  8'h63;        memory[59244] <=  8'h73;        memory[59245] <=  8'h66;        memory[59246] <=  8'h72;        memory[59247] <=  8'h74;        memory[59248] <=  8'h79;        memory[59249] <=  8'h75;        memory[59250] <=  8'h6a;        memory[59251] <=  8'h6e;        memory[59252] <=  8'h62;        memory[59253] <=  8'h76;        memory[59254] <=  8'h63;        memory[59255] <=  8'h64;        memory[59256] <=  8'h74;        memory[59257] <=  8'h79;        memory[59258] <=  8'h75;        memory[59259] <=  8'h69;        memory[59260] <=  8'h6b;        memory[59261] <=  8'h6d;        memory[59262] <=  8'h6e;        memory[59263] <=  8'h62;        memory[59264] <=  8'h76;        memory[59265] <=  8'h63;        memory[59266] <=  8'h78;        memory[59267] <=  8'h73;        memory[59268] <=  8'h64;        memory[59269] <=  8'h72;        memory[59270] <=  8'h74;        memory[59271] <=  8'h79;        memory[59272] <=  8'h75;        memory[59273] <=  8'h69;        memory[59274] <=  8'h6b;        memory[59275] <=  8'h6d;        memory[59276] <=  8'h6e;        memory[59277] <=  8'h62;        memory[59278] <=  8'h76;        memory[59279] <=  8'h63;        memory[59280] <=  8'h73;        memory[59281] <=  8'h77;        memory[59282] <=  8'h33;        memory[59283] <=  8'h34;        memory[59284] <=  8'h35;        memory[59285] <=  8'h36;        memory[59286] <=  8'h37;        memory[59287] <=  8'h38;        memory[59288] <=  8'h69;        memory[59289] <=  8'h6b;        memory[59290] <=  8'h6d;        memory[59291] <=  8'h6e;        memory[59292] <=  8'h62;        memory[59293] <=  8'h76;        memory[59294] <=  8'h63;        memory[59295] <=  8'h64;        memory[59296] <=  8'h65;        memory[59297] <=  8'h72;        memory[59298] <=  8'h36;        memory[59299] <=  8'h37;        memory[59300] <=  8'h38;        memory[59301] <=  8'h69;        memory[59302] <=  8'h6f;        memory[59303] <=  8'h6b;        memory[59304] <=  8'h6a;        memory[59305] <=  8'h6e;        memory[59306] <=  8'h62;        memory[59307] <=  8'h76;        memory[59308] <=  8'h63;        memory[59309] <=  8'h64;        memory[59310] <=  8'h72;        memory[59311] <=  8'h74;        memory[59312] <=  8'h79;        memory[59313] <=  8'h75;        memory[59314] <=  8'h73;        memory[59315] <=  8'h6a;        memory[59316] <=  8'h63;        memory[59317] <=  8'h6e;        memory[59318] <=  8'h62;        memory[59319] <=  8'h64;        memory[59320] <=  8'h66;        memory[59321] <=  8'h73;        memory[59322] <=  8'h74;        memory[59323] <=  8'h79;        memory[59324] <=  8'h75;        memory[59325] <=  8'h61;        memory[59326] <=  8'h69;        memory[59327] <=  8'h6b;        memory[59328] <=  8'h78;        memory[59329] <=  8'h6d;        memory[59330] <=  8'h6e;        memory[59331] <=  8'h73;        memory[59332] <=  8'h6a;        memory[59333] <=  8'h6f;        memory[59334] <=  8'h64;        memory[59335] <=  8'h6c;        memory[59336] <=  8'h63;        memory[59337] <=  8'h78;        memory[59338] <=  8'h2c;        memory[59339] <=  8'h6d;        memory[59340] <=  8'h73;        memory[59341] <=  8'h6b;        memory[59342] <=  8'h64;        memory[59343] <=  8'h6c;        memory[59344] <=  8'h70;        memory[59345] <=  8'h5b;        memory[59346] <=  8'h3b;        memory[59347] <=  8'h73;        memory[59348] <=  8'h6c;        memory[59349] <=  8'h64;        memory[59350] <=  8'h70;        memory[59351] <=  8'h76;        memory[59352] <=  8'h63;        memory[59353] <=  8'h5b;        memory[59354] <=  8'h78;        memory[59355] <=  8'h76;        memory[59356] <=  8'h63;        memory[59357] <=  8'h5b;        memory[59358] <=  8'h78;        memory[59359] <=  8'h70;        memory[59360] <=  8'h6f;        memory[59361] <=  8'h20;        memory[59362] <=  8'h62;        memory[59363] <=  8'h61;        memory[59364] <=  8'h72;        memory[59365] <=  8'h74;        memory[59366] <=  8'h74;        memory[59367] <=  8'h62;        memory[59368] <=  8'h61;        memory[59369] <=  8'h72;        memory[59370] <=  8'h74;        memory[59371] <=  8'h78;        memory[59372] <=  8'h61;        memory[59373] <=  8'h74;        memory[59374] <=  8'h6b;        memory[59375] <=  8'h73;        memory[59376] <=  8'h68;        memory[59377] <=  8'h63;        memory[59378] <=  8'h66;        memory[59379] <=  8'h69;        memory[59380] <=  8'h77;        memory[59381] <=  8'h68;        memory[59382] <=  8'h61;        memory[59383] <=  8'h69;        memory[59384] <=  8'h6a;        memory[59385] <=  8'h78;        memory[59386] <=  8'h5d;        memory[59387] <=  8'h65;        memory[59388] <=  8'h6b;        memory[59389] <=  8'h6f;        memory[59390] <=  8'h39;        memory[59391] <=  8'h64;        memory[59392] <=  8'h75;        memory[59393] <=  8'h38;        memory[59394] <=  8'h79;        memory[59395] <=  8'h20;        memory[59396] <=  8'h37;        memory[59397] <=  8'h63;        memory[59398] <=  8'h67;        memory[59399] <=  8'h78;        memory[59400] <=  8'h63;        memory[59401] <=  8'h75;        memory[59402] <=  8'h68;        memory[59403] <=  8'h69;        memory[59404] <=  8'h6a;        memory[59405] <=  8'h77;        memory[59406] <=  8'h69;        memory[59407] <=  8'h64;        memory[59408] <=  8'h66;        memory[59409] <=  8'h68;        memory[59410] <=  8'h75;        memory[59411] <=  8'h76;        memory[59412] <=  8'h64;        memory[59413] <=  8'h62;        memory[59414] <=  8'h66;        memory[59415] <=  8'h6a;        memory[59416] <=  8'h6e;        memory[59417] <=  8'h6b;        memory[59418] <=  8'h6a;        memory[59419] <=  8'h65;        memory[59420] <=  8'h38;        memory[59421] <=  8'h66;        memory[59422] <=  8'h37;        memory[59423] <=  8'h67;        memory[59424] <=  8'h79;        memory[59425] <=  8'h76;        memory[59426] <=  8'h63;        memory[59427] <=  8'h68;        memory[59428] <=  8'h69;        memory[59429] <=  8'h6a;        memory[59430] <=  8'h33;        memory[59431] <=  8'h65;        memory[59432] <=  8'h67;        memory[59433] <=  8'h79;        memory[59434] <=  8'h72;        memory[59435] <=  8'h64;        memory[59436] <=  8'h62;        memory[59437] <=  8'h6e;        memory[59438] <=  8'h63;        memory[59439] <=  8'h7a;        memory[59440] <=  8'h6a;        memory[59441] <=  8'h6f;        memory[59442] <=  8'h66;        memory[59443] <=  8'h78;        memory[59444] <=  8'h6a;        memory[59445] <=  8'h69;        memory[59446] <=  8'h63;        memory[59447] <=  8'h68;        memory[59448] <=  8'h62;        memory[59449] <=  8'h6e;        memory[59450] <=  8'h6d;        memory[59451] <=  8'h63;        memory[59452] <=  8'h73;        memory[59453] <=  8'h6c;        memory[59454] <=  8'h6b;        memory[59455] <=  8'h6a;        memory[59456] <=  8'h69;        memory[59457] <=  8'h68;        memory[59458] <=  8'h76;        memory[59459] <=  8'h75;        memory[59460] <=  8'h69;        memory[59461] <=  8'h64;        memory[59462] <=  8'h68;        memory[59463] <=  8'h75;        memory[59464] <=  8'h67;        memory[59465] <=  8'h79;        memory[59466] <=  8'h62;        memory[59467] <=  8'h68;        memory[59468] <=  8'h65;        memory[59469] <=  8'h6a;        memory[59470] <=  8'h72;        memory[59471] <=  8'h6b;        memory[59472] <=  8'h6a;        memory[59473] <=  8'h6f;        memory[59474] <=  8'h64;        memory[59475] <=  8'h67;        memory[59476] <=  8'h69;        memory[59477] <=  8'h75;        memory[59478] <=  8'h69;        memory[59479] <=  8'h67;        memory[59480] <=  8'h76;        memory[59481] <=  8'h79;        memory[59482] <=  8'h75;        memory[59483] <=  8'h67;        memory[59484] <=  8'h78;        memory[59485] <=  8'h68;        memory[59486] <=  8'h63;        memory[59487] <=  8'h20;        memory[59488] <=  8'h20;        memory[59489] <=  8'h20;        memory[59490] <=  8'h78;        memory[59491] <=  8'h76;        memory[59492] <=  8'h20;        memory[59493] <=  8'h63;        memory[59494] <=  8'h78;        memory[59495] <=  8'h67;        memory[59496] <=  8'h79;        memory[59497] <=  8'h63;        memory[59498] <=  8'h75;        memory[59499] <=  8'h68;        memory[59500] <=  8'h6a;        memory[59501] <=  8'h6b;        memory[59502] <=  8'h61;        memory[59503] <=  8'h6c;        memory[59504] <=  8'h78;        memory[59505] <=  8'h76;        memory[59506] <=  8'h70;        memory[59507] <=  8'h6f;        memory[59508] <=  8'h69;        memory[59509] <=  8'h6a;        memory[59510] <=  8'h69;        memory[59511] <=  8'h68;        memory[59512] <=  8'h6a;        memory[59513] <=  8'h62;        memory[59514] <=  8'h77;        memory[59515] <=  8'h65;        memory[59516] <=  8'h6e;        memory[59517] <=  8'h61;        memory[59518] <=  8'h66;        memory[59519] <=  8'h6d;        memory[59520] <=  8'h64;        memory[59521] <=  8'h6b;        memory[59522] <=  8'h6d;        memory[59523] <=  8'h76;        memory[59524] <=  8'h6c;        memory[59525] <=  8'h63;        memory[59526] <=  8'h6f;        memory[59527] <=  8'h64;        memory[59528] <=  8'h69;        memory[59529] <=  8'h75;        memory[59530] <=  8'h68;        memory[59531] <=  8'h73;        memory[59532] <=  8'h66;        memory[59533] <=  8'h65;        memory[59534] <=  8'h62;        memory[59535] <=  8'h6e;        memory[59536] <=  8'h64;        memory[59537] <=  8'h73;        memory[59538] <=  8'h63;        memory[59539] <=  8'h6b;        memory[59540] <=  8'h20;        memory[59541] <=  8'h78;        memory[59542] <=  8'h6a;        memory[59543] <=  8'h78;        memory[59544] <=  8'h63;        memory[59545] <=  8'h73;        memory[59546] <=  8'h64;        memory[59547] <=  8'h66;        memory[59548] <=  8'h6b;        memory[59549] <=  8'h64;        memory[59550] <=  8'h6e;        memory[59551] <=  8'h6d;        memory[59552] <=  8'h64;        memory[59553] <=  8'h73;        memory[59554] <=  8'h63;        memory[59555] <=  8'h6b;        memory[59556] <=  8'h78;        memory[59557] <=  8'h6c;        memory[59558] <=  8'h6f;        memory[59559] <=  8'h66;        memory[59560] <=  8'h6a;        memory[59561] <=  8'h69;        memory[59562] <=  8'h61;        memory[59563] <=  8'h62;        memory[59564] <=  8'h6e;        memory[59565] <=  8'h20;        memory[59566] <=  8'h78;        memory[59567] <=  8'h6b;        memory[59568] <=  8'h6d;        memory[59569] <=  8'h20;        memory[59570] <=  8'h6f;        memory[59571] <=  8'h63;        memory[59572] <=  8'h76;        memory[59573] <=  8'h73;        memory[59574] <=  8'h64;        memory[59575] <=  8'h69;        memory[59576] <=  8'h66;        memory[59577] <=  8'h68;        memory[59578] <=  8'h65;        memory[59579] <=  8'h71;        memory[59580] <=  8'h6a;        memory[59581] <=  8'h77;        memory[59582] <=  8'h62;        memory[59583] <=  8'h65;        memory[59584] <=  8'h6e;        memory[59585] <=  8'h20;        memory[59586] <=  8'h6d;        memory[59587] <=  8'h64;        memory[59588] <=  8'h73;        memory[59589] <=  8'h6c;        memory[59590] <=  8'h76;        memory[59591] <=  8'h6b;        memory[59592] <=  8'h63;        memory[59593] <=  8'h78;        memory[59594] <=  8'h20;        memory[59595] <=  8'h6f;        memory[59596] <=  8'h78;        memory[59597] <=  8'h69;        memory[59598] <=  8'h63;        memory[59599] <=  8'h6a;        memory[59600] <=  8'h76;        memory[59601] <=  8'h64;        memory[59602] <=  8'h66;        memory[59603] <=  8'h65;        memory[59604] <=  8'h71;        memory[59605] <=  8'h6e;        memory[59606] <=  8'h20;        memory[59607] <=  8'h64;        memory[59608] <=  8'h6d;        memory[59609] <=  8'h73;        memory[59610] <=  8'h6c;        memory[59611] <=  8'h63;        memory[59612] <=  8'h78;        memory[59613] <=  8'h6b;        memory[59614] <=  8'h20;        memory[59615] <=  8'h6f;        memory[59616] <=  8'h78;        memory[59617] <=  8'h63;        memory[59618] <=  8'h76;        memory[59619] <=  8'h6a;        memory[59620] <=  8'h64;        memory[59621] <=  8'h62;        memory[59622] <=  8'h71;        memory[59623] <=  8'h77;        memory[59624] <=  8'h65;        memory[59625] <=  8'h6e;        memory[59626] <=  8'h6d;        memory[59627] <=  8'h64;        memory[59628] <=  8'h6c;        memory[59629] <=  8'h73;        memory[59630] <=  8'h2c;        memory[59631] <=  8'h76;        memory[59632] <=  8'h63;        memory[59633] <=  8'h78;        memory[59634] <=  8'h20;        memory[59635] <=  8'h63;        memory[59636] <=  8'h6f;        memory[59637] <=  8'h69;        memory[59638] <=  8'h76;        memory[59639] <=  8'h68;        memory[59640] <=  8'h73;        memory[59641] <=  8'h64;        memory[59642] <=  8'h62;        memory[59643] <=  8'h71;        memory[59644] <=  8'h77;        memory[59645] <=  8'h65;        memory[59646] <=  8'h6e;        memory[59647] <=  8'h64;        memory[59648] <=  8'h6b;        memory[59649] <=  8'h73;        memory[59650] <=  8'h76;        memory[59651] <=  8'h6f;        memory[59652] <=  8'h63;        memory[59653] <=  8'h20;        memory[59654] <=  8'h76;        memory[59655] <=  8'h69;        memory[59656] <=  8'h75;        memory[59657] <=  8'h69;        memory[59658] <=  8'h68;        memory[59659] <=  8'h63;        memory[59660] <=  8'h78;        memory[59661] <=  8'h69;        memory[59662] <=  8'h6f;        memory[59663] <=  8'h76;        memory[59664] <=  8'h73;        memory[59665] <=  8'h64;        memory[59666] <=  8'h61;        memory[59667] <=  8'h64;        memory[59668] <=  8'h6e;        memory[59669] <=  8'h77;        memory[59670] <=  8'h71;        memory[59671] <=  8'h6b;        memory[59672] <=  8'h6c;        memory[59673] <=  8'h73;        memory[59674] <=  8'h76;        memory[59675] <=  8'h6e;        memory[59676] <=  8'h62;        memory[59677] <=  8'h20;        memory[59678] <=  8'h64;        memory[59679] <=  8'h66;        memory[59680] <=  8'h6a;        memory[59681] <=  8'h6b;        memory[59682] <=  8'h71;        memory[59683] <=  8'h64;        memory[59684] <=  8'h77;        memory[59685] <=  8'h65;        memory[59686] <=  8'h6e;        memory[59687] <=  8'h62;        memory[59688] <=  8'h20;        memory[59689] <=  8'h64;        memory[59690] <=  8'h73;        memory[59691] <=  8'h76;        memory[59692] <=  8'h68;        memory[59693] <=  8'h64;        memory[59694] <=  8'h61;        memory[59695] <=  8'h71;        memory[59696] <=  8'h77;        memory[59697] <=  8'h6a;        memory[59698] <=  8'h65;        memory[59699] <=  8'h6e;        memory[59700] <=  8'h64;        memory[59701] <=  8'h20;        memory[59702] <=  8'h61;        memory[59703] <=  8'h63;        memory[59704] <=  8'h62;        memory[59705] <=  8'h68;        memory[59706] <=  8'h64;        memory[59707] <=  8'h61;        memory[59708] <=  8'h77;        memory[59709] <=  8'h71;        memory[59710] <=  8'h6e;        memory[59711] <=  8'h20;        memory[59712] <=  8'h62;        memory[59713] <=  8'h73;        memory[59714] <=  8'h76;        memory[59715] <=  8'h61;        memory[59716] <=  8'h67;        memory[59717] <=  8'h76;        memory[59718] <=  8'h68;        memory[59719] <=  8'h67;        memory[59720] <=  8'h61;        memory[59721] <=  8'h73;        memory[59722] <=  8'h6a;        memory[59723] <=  8'h6b;        memory[59724] <=  8'h63;        memory[59725] <=  8'h78;        memory[59726] <=  8'h76;        memory[59727] <=  8'h6e;        memory[59728] <=  8'h73;        memory[59729] <=  8'h64;        memory[59730] <=  8'h20;        memory[59731] <=  8'h66;        memory[59732] <=  8'h62;        memory[59733] <=  8'h64;        memory[59734] <=  8'h61;        memory[59735] <=  8'h73;        memory[59736] <=  8'h76;        memory[59737] <=  8'h67;        memory[59738] <=  8'h63;        memory[59739] <=  8'h79;        memory[59740] <=  8'h7a;        memory[59741] <=  8'h78;        memory[59742] <=  8'h79;        memory[59743] <=  8'h75;        memory[59744] <=  8'h20;        memory[59745] <=  8'h69;        memory[59746] <=  8'h6a;        memory[59747] <=  8'h64;        memory[59748] <=  8'h66;        memory[59749] <=  8'h6b;        memory[59750] <=  8'h61;        memory[59751] <=  8'h64;        memory[59752] <=  8'h63;        memory[59753] <=  8'h78;        memory[59754] <=  8'h68;        memory[59755] <=  8'h20;        memory[59756] <=  8'h67;        memory[59757] <=  8'h61;        memory[59758] <=  8'h68;        memory[59759] <=  8'h75;        memory[59760] <=  8'h64;        memory[59761] <=  8'h73;        memory[59762] <=  8'h69;        memory[59763] <=  8'h6a;        memory[59764] <=  8'h61;        memory[59765] <=  8'h6b;        memory[59766] <=  8'h63;        memory[59767] <=  8'h62;        memory[59768] <=  8'h61;        memory[59769] <=  8'h72;        memory[59770] <=  8'h73;        memory[59771] <=  8'h68;        memory[59772] <=  8'h64;        memory[59773] <=  8'h66;        memory[59774] <=  8'h67;        memory[59775] <=  8'h73;        memory[59776] <=  8'h68;        memory[59777] <=  8'h64;        memory[59778] <=  8'h66;        memory[59779] <=  8'h68;        memory[59780] <=  8'h64;        memory[59781] <=  8'h6a;        memory[59782] <=  8'h68;        memory[59783] <=  8'h62;        memory[59784] <=  8'h67;        memory[59785] <=  8'h63;        memory[59786] <=  8'h61;        memory[59787] <=  8'h66;        memory[59788] <=  8'h73;        memory[59789] <=  8'h79;        memory[59790] <=  8'h67;        memory[59791] <=  8'h6b;        memory[59792] <=  8'h75;        memory[59793] <=  8'h64;        memory[59794] <=  8'h68;        memory[59795] <=  8'h62;        memory[59796] <=  8'h77;        memory[59797] <=  8'h76;        memory[59798] <=  8'h67;        memory[59799] <=  8'h61;        memory[59800] <=  8'h66;        memory[59801] <=  8'h64;        memory[59802] <=  8'h74;        memory[59803] <=  8'h75;        memory[59804] <=  8'h66;        memory[59805] <=  8'h79;        memory[59806] <=  8'h67;        memory[59807] <=  8'h69;        memory[59808] <=  8'h75;        memory[59809] <=  8'h68;        memory[59810] <=  8'h6c;        memory[59811] <=  8'h6a;        memory[59812] <=  8'h62;        memory[59813] <=  8'h6b;        memory[59814] <=  8'h68;        memory[59815] <=  8'h76;        memory[59816] <=  8'h67;        memory[59817] <=  8'h63;        memory[59818] <=  8'h66;        memory[59819] <=  8'h78;        memory[59820] <=  8'h64;        memory[59821] <=  8'h74;        memory[59822] <=  8'h75;        memory[59823] <=  8'h79;        memory[59824] <=  8'h69;        memory[59825] <=  8'h75;        memory[59826] <=  8'h68;        memory[59827] <=  8'h6c;        memory[59828] <=  8'h6a;        memory[59829] <=  8'h6b;        memory[59830] <=  8'h67;        memory[59831] <=  8'h6a;        memory[59832] <=  8'h63;        memory[59833] <=  8'h66;        memory[59834] <=  8'h68;        memory[59835] <=  8'h64;        memory[59836] <=  8'h67;        memory[59837] <=  8'h72;        memory[59838] <=  8'h79;        memory[59839] <=  8'h74;        memory[59840] <=  8'h66;        memory[59841] <=  8'h75;        memory[59842] <=  8'h79;        memory[59843] <=  8'h69;        memory[59844] <=  8'h68;        memory[59845] <=  8'h6c;        memory[59846] <=  8'h62;        memory[59847] <=  8'h6d;        memory[59848] <=  8'h76;        memory[59849] <=  8'h6e;        memory[59850] <=  8'h63;        memory[59851] <=  8'h66;        memory[59852] <=  8'h68;        memory[59853] <=  8'h64;        memory[59854] <=  8'h74;        memory[59855] <=  8'h75;        memory[59856] <=  8'h67;        memory[59857] <=  8'h79;        memory[59858] <=  8'h69;        memory[59859] <=  8'h68;        memory[59860] <=  8'h75;        memory[59861] <=  8'h6a;        memory[59862] <=  8'h6c;        memory[59863] <=  8'h62;        memory[59864] <=  8'h6d;        memory[59865] <=  8'h76;        memory[59866] <=  8'h6e;        memory[59867] <=  8'h63;        memory[59868] <=  8'h66;        memory[59869] <=  8'h68;        memory[59870] <=  8'h67;        memory[59871] <=  8'h79;        memory[59872] <=  8'h68;        memory[59873] <=  8'h75;        memory[59874] <=  8'h6a;        memory[59875] <=  8'h6e;        memory[59876] <=  8'h2c;        memory[59877] <=  8'h62;        memory[59878] <=  8'h6e;        memory[59879] <=  8'h6d;        memory[59880] <=  8'h76;        memory[59881] <=  8'h6e;        memory[59882] <=  8'h63;        memory[59883] <=  8'h66;        memory[59884] <=  8'h68;        memory[59885] <=  8'h74;        memory[59886] <=  8'h79;        memory[59887] <=  8'h69;        memory[59888] <=  8'h75;        memory[59889] <=  8'h6c;        memory[59890] <=  8'h6a;        memory[59891] <=  8'h62;        memory[59892] <=  8'h6d;        memory[59893] <=  8'h76;        memory[59894] <=  8'h6e;        memory[59895] <=  8'h63;        memory[59896] <=  8'h66;        memory[59897] <=  8'h74;        memory[59898] <=  8'h75;        memory[59899] <=  8'h79;        memory[59900] <=  8'h69;        memory[59901] <=  8'h68;        memory[59902] <=  8'h6b;        memory[59903] <=  8'h62;        memory[59904] <=  8'h76;        memory[59905] <=  8'h63;        memory[59906] <=  8'h66;        memory[59907] <=  8'h67;        memory[59908] <=  8'h74;        memory[59909] <=  8'h75;        memory[59910] <=  8'h79;        memory[59911] <=  8'h69;        memory[59912] <=  8'h75;        memory[59913] <=  8'h68;        memory[59914] <=  8'h6a;        memory[59915] <=  8'h6b;        memory[59916] <=  8'h62;        memory[59917] <=  8'h76;        memory[59918] <=  8'h63;        memory[59919] <=  8'h66;        memory[59920] <=  8'h74;        memory[59921] <=  8'h75;        memory[59922] <=  8'h79;        memory[59923] <=  8'h69;        memory[59924] <=  8'h75;        memory[59925] <=  8'h6a;        memory[59926] <=  8'h6b;        memory[59927] <=  8'h6e;        memory[59928] <=  8'h62;        memory[59929] <=  8'h76;        memory[59930] <=  8'h67;        memory[59931] <=  8'h66;        memory[59932] <=  8'h74;        memory[59933] <=  8'h79;        memory[59934] <=  8'h75;        memory[59935] <=  8'h75;        memory[59936] <=  8'h69;        memory[59937] <=  8'h6a;        memory[59938] <=  8'h6b;        memory[59939] <=  8'h68;        memory[59940] <=  8'h62;        memory[59941] <=  8'h6a;        memory[59942] <=  8'h67;        memory[59943] <=  8'h68;        memory[59944] <=  8'h66;        memory[59945] <=  8'h79;        memory[59946] <=  8'h74;        memory[59947] <=  8'h79;        memory[59948] <=  8'h69;        memory[59949] <=  8'h75;        memory[59950] <=  8'h64;        memory[59951] <=  8'h6a;        memory[59952] <=  8'h6b;        memory[59953] <=  8'h68;        memory[59954] <=  8'h63;        memory[59955] <=  8'h7a;        memory[59956] <=  8'h67;        memory[59957] <=  8'h68;        memory[59958] <=  8'h74;        memory[59959] <=  8'h75;        memory[59960] <=  8'h79;        memory[59961] <=  8'h69;        memory[59962] <=  8'h61;        memory[59963] <=  8'h73;        memory[59964] <=  8'h75;        memory[59965] <=  8'h6a;        memory[59966] <=  8'h6b;        memory[59967] <=  8'h62;        memory[59968] <=  8'h6e;        memory[59969] <=  8'h61;        memory[59970] <=  8'h76;        memory[59971] <=  8'h63;        memory[59972] <=  8'h66;        memory[59973] <=  8'h68;        memory[59974] <=  8'h75;        memory[59975] <=  8'h61;        memory[59976] <=  8'h73;        memory[59977] <=  8'h79;        memory[59978] <=  8'h64;        memory[59979] <=  8'h75;        memory[59980] <=  8'h69;        memory[59981] <=  8'h6a;        memory[59982] <=  8'h61;        memory[59983] <=  8'h6b;        memory[59984] <=  8'h62;        memory[59985] <=  8'h63;        memory[59986] <=  8'h78;        memory[59987] <=  8'h68;        memory[59988] <=  8'h67;        memory[59989] <=  8'h79;        memory[59990] <=  8'h75;        memory[59991] <=  8'h7a;        memory[59992] <=  8'h63;        memory[59993] <=  8'h61;        memory[59994] <=  8'h73;        memory[59995] <=  8'h69;        memory[59996] <=  8'h75;        memory[59997] <=  8'h6f;        memory[59998] <=  8'h69;        memory[59999] <=  8'h6a;        memory[60000] <=  8'h61;        memory[60001] <=  8'h6c;        memory[60002] <=  8'h63;        memory[60003] <=  8'h78;        memory[60004] <=  8'h62;        memory[60005] <=  8'h63;        memory[60006] <=  8'h20;        memory[60007] <=  8'h6e;        memory[60008] <=  8'h76;        memory[60009] <=  8'h63;        memory[60010] <=  8'h61;        memory[60011] <=  8'h64;        memory[60012] <=  8'h73;        memory[60013] <=  8'h67;        memory[60014] <=  8'h79;        memory[60015] <=  8'h68;        memory[60016] <=  8'h75;        memory[60017] <=  8'h61;        memory[60018] <=  8'h6a;        memory[60019] <=  8'h6b;        memory[60020] <=  8'h78;        memory[60021] <=  8'h62;        memory[60022] <=  8'h20;        memory[60023] <=  8'h6e;        memory[60024] <=  8'h76;        memory[60025] <=  8'h63;        memory[60026] <=  8'h61;        memory[60027] <=  8'h73;        memory[60028] <=  8'h67;        memory[60029] <=  8'h68;        memory[60030] <=  8'h75;        memory[60031] <=  8'h6a;        memory[60032] <=  8'h6c;        memory[60033] <=  8'h6b;        memory[60034] <=  8'h63;        memory[60035] <=  8'h78;        memory[60036] <=  8'h20;        memory[60037] <=  8'h6a;        memory[60038] <=  8'h6b;        memory[60039] <=  8'h68;        memory[60040] <=  8'h61;        memory[60041] <=  8'h73;        memory[60042] <=  8'h76;        memory[60043] <=  8'h64;        memory[60044] <=  8'h6e;        memory[60045] <=  8'h20;        memory[60046] <=  8'h62;        memory[60047] <=  8'h6e;        memory[60048] <=  8'h6d;        memory[60049] <=  8'h6b;        memory[60050] <=  8'h77;        memory[60051] <=  8'h64;        memory[60052] <=  8'h6f;        memory[60053] <=  8'h77;        memory[60054] <=  8'h69;        memory[60055] <=  8'h6f;        memory[60056] <=  8'h75;        memory[60057] <=  8'h69;        memory[60058] <=  8'h68;        memory[60059] <=  8'h62;        memory[60060] <=  8'h6e;        memory[60061] <=  8'h6b;        memory[60062] <=  8'h77;        memory[60063] <=  8'h69;        memory[60064] <=  8'h6f;        memory[60065] <=  8'h75;        memory[60066] <=  8'h71;        memory[60067] <=  8'h69;        memory[60068] <=  8'h79;        memory[60069] <=  8'h67;        memory[60070] <=  8'h6a;        memory[60071] <=  8'h64;        memory[60072] <=  8'h61;        memory[60073] <=  8'h76;        memory[60074] <=  8'h62;        memory[60075] <=  8'h6e;        memory[60076] <=  8'h6b;        memory[60077] <=  8'h6f;        memory[60078] <=  8'h70;        memory[60079] <=  8'h64;        memory[60080] <=  8'h76;        memory[60081] <=  8'h69;        memory[60082] <=  8'h6f;        memory[60083] <=  8'h75;        memory[60084] <=  8'h69;        memory[60085] <=  8'h48;        memory[60086] <=  8'h42;        memory[60087] <=  8'h6b;        memory[60088] <=  8'h64;        memory[60089] <=  8'h6e;        memory[60090] <=  8'h6c;        memory[60091] <=  8'h71;        memory[60092] <=  8'h6b;        memory[60093] <=  8'h6d;        memory[60094] <=  8'h6a;        memory[60095] <=  8'h70;        memory[60096] <=  8'h69;        memory[60097] <=  8'h6f;        memory[60098] <=  8'h68;        memory[60099] <=  8'h65;        memory[60100] <=  8'h66;        memory[60101] <=  8'h75;        memory[60102] <=  8'h67;        memory[60103] <=  8'h69;        memory[60104] <=  8'h73;        memory[60105] <=  8'h61;        memory[60106] <=  8'h62;        memory[60107] <=  8'h64;        memory[60108] <=  8'h6b;        memory[60109] <=  8'h6a;        memory[60110] <=  8'h6b;        memory[60111] <=  8'h6c;        memory[60112] <=  8'h6a;        memory[60113] <=  8'h69;        memory[60114] <=  8'h73;        memory[60115] <=  8'h6f;        memory[60116] <=  8'h71;        memory[60117] <=  8'h68;        memory[60118] <=  8'h77;        memory[60119] <=  8'h67;        memory[60120] <=  8'h69;        memory[60121] <=  8'h79;        memory[60122] <=  8'h6a;        memory[60123] <=  8'h64;        memory[60124] <=  8'h76;        memory[60125] <=  8'h62;        memory[60126] <=  8'h6e;        memory[60127] <=  8'h61;        memory[60128] <=  8'h73;        memory[60129] <=  8'h66;        memory[60130] <=  8'h6c;        memory[60131] <=  8'h6b;        memory[60132] <=  8'h64;        memory[60133] <=  8'h6a;        memory[60134] <=  8'h68;        memory[60135] <=  8'h63;        memory[60136] <=  8'h67;        memory[60137] <=  8'h6a;        memory[60138] <=  8'h76;        memory[60139] <=  8'h73;        memory[60140] <=  8'h64;        memory[60141] <=  8'h62;        memory[60142] <=  8'h62;        memory[60143] <=  8'h61;        memory[60144] <=  8'h72;        memory[60145] <=  8'h62;        memory[60146] <=  8'h62;        memory[60147] <=  8'h73;        memory[60148] <=  8'h62;        memory[60149] <=  8'h67;        memory[60150] <=  8'h73;        memory[60151] <=  8'h66;        memory[60152] <=  8'h67;        memory[60153] <=  8'h61;        memory[60154] <=  8'h68;        memory[60155] <=  8'h66;        memory[60156] <=  8'h73;        memory[60157] <=  8'h68;        memory[60158] <=  8'h61;        memory[60159] <=  8'h66;        memory[60160] <=  8'h73;        memory[60161] <=  8'h66;        memory[60162] <=  8'h68;        memory[60163] <=  8'h61;        memory[60164] <=  8'h69;        memory[60165] <=  8'h64;        memory[60166] <=  8'h75;        memory[60167] <=  8'h67;        memory[60168] <=  8'h64;        memory[60169] <=  8'h77;        memory[60170] <=  8'h62;        memory[60171] <=  8'h61;        memory[60172] <=  8'h62;        memory[60173] <=  8'h72;        memory[60174] <=  8'h62;        memory[60175] <=  8'h61;        memory[60176] <=  8'h62;        memory[60177] <=  8'h62;        memory[60178] <=  8'h74;        memory[60179] <=  8'h62;        memory[60180] <=  8'h62;        memory[60181] <=  8'h62;        memory[60182] <=  8'h62;        memory[60183] <=  8'h62;        memory[60184] <=  8'h62;        memory[60185] <=  8'h62;        memory[60186] <=  8'h62;        memory[60187] <=  8'h61;        memory[60188] <=  8'h62;        memory[60189] <=  8'h62;        memory[60190] <=  8'h72;        memory[60191] <=  8'h74;        memory[60192] <=  8'h62;        memory[60193] <=  8'h62;        memory[60194] <=  8'h61;        memory[60195] <=  8'h62;        memory[60196] <=  8'h72;        memory[60197] <=  8'h62;        memory[60198] <=  8'h74;        memory[60199] <=  8'h62;        memory[60200] <=  8'h62;        memory[60201] <=  8'h62;        memory[60202] <=  8'h63;        memory[60203] <=  8'h61;        memory[60204] <=  8'h72;        memory[60205] <=  8'h74;        memory[60206] <=  8'h73;        memory[60207] <=  8'h62;        memory[60208] <=  8'h61;        memory[60209] <=  8'h72;        memory[60210] <=  8'h74;        memory[60211] <=  8'h74;        memory[60212] <=  8'h62;        memory[60213] <=  8'h61;        memory[60214] <=  8'h72;        memory[60215] <=  8'h74;        memory[60216] <=  8'h78;        memory[60217] <=  8'h61;        memory[60218] <=  8'h74;        memory[60219] <=  8'h6b;        memory[60220] <=  8'h73;        memory[60221] <=  8'h68;        memory[60222] <=  8'h63;        memory[60223] <=  8'h66;        memory[60224] <=  8'h69;        memory[60225] <=  8'h77;        memory[60226] <=  8'h68;        memory[60227] <=  8'h61;        memory[60228] <=  8'h74;        memory[60229] <=  8'h61;        memory[60230] <=  8'h6e;        memory[60231] <=  8'h61;        memory[60232] <=  8'h62;        memory[60233] <=  8'h61;        memory[60234] <=  8'h63;        memory[60235] <=  8'h61;        memory[60236] <=  8'h74;        memory[60237] <=  8'h61;        memory[60238] <=  8'h62;        memory[60239] <=  8'h61;        memory[60240] <=  8'h72;        memory[60241] <=  8'h63;        memory[60242] <=  8'h61;        memory[60243] <=  8'h68;        memory[60244] <=  8'h64;        memory[60245] <=  8'h75;        memory[60246] <=  8'h63;        memory[60247] <=  8'h74;        memory[60248] <=  8'h61;        memory[60249] <=  8'h64;        memory[60250] <=  8'h61;        memory[60251] <=  8'h61;        memory[60252] <=  8'h63;        memory[60253] <=  8'h61;        memory[60254] <=  8'h72;        memory[60255] <=  8'h63;        memory[60256] <=  8'h74;        memory[60257] <=  8'h72;        memory[60258] <=  8'h63;        memory[60259] <=  8'h61;        memory[60260] <=  8'h74;        memory[60261] <=  8'h72;        memory[60262] <=  8'h63;        memory[60263] <=  8'h61;        memory[60264] <=  8'h74;        memory[60265] <=  8'h63;        memory[60266] <=  8'h62;        memory[60267] <=  8'h61;        memory[60268] <=  8'h74;        memory[60269] <=  8'h62;        memory[60270] <=  8'h72;        memory[60271] <=  8'h63;        memory[60272] <=  8'h61;        memory[60273] <=  8'h74;        memory[60274] <=  8'h72;        memory[60275] <=  8'h6e;        memory[60276] <=  8'h62;        memory[60277] <=  8'h61;        memory[60278] <=  8'h63;        memory[60279] <=  8'h61;        memory[60280] <=  8'h74;        memory[60281] <=  8'h79;        memory[60282] <=  8'h73;        memory[60283] <=  8'h6e;        memory[60284] <=  8'h63;        memory[60285] <=  8'h74;        memory[60286] <=  8'h61;        memory[60287] <=  8'h6e;        memory[60288] <=  8'h62;        memory[60289] <=  8'h61;        memory[60290] <=  8'h63;        memory[60291] <=  8'h72;        memory[60292] <=  8'h6e;        memory[60293] <=  8'h74;        memory[60294] <=  8'h61;        memory[60295] <=  8'h62;        memory[60296] <=  8'h74;        memory[60297] <=  8'h6e;        memory[60298] <=  8'h61;        memory[60299] <=  8'h72;        memory[60300] <=  8'h62;        memory[60301] <=  8'h78;        memory[60302] <=  8'h74;        memory[60303] <=  8'h61;        memory[60304] <=  8'h72;        memory[60305] <=  8'h62;        memory[60306] <=  8'h61;        memory[60307] <=  8'h72;        memory[60308] <=  8'h74;        memory[60309] <=  8'h74;        memory[60310] <=  8'h62;        memory[60311] <=  8'h61;        memory[60312] <=  8'h72;        memory[60313] <=  8'h74;        memory[60314] <=  8'h78;        memory[60315] <=  8'h61;        memory[60316] <=  8'h74;        memory[60317] <=  8'h6b;        memory[60318] <=  8'h73;        memory[60319] <=  8'h68;        memory[60320] <=  8'h63;        memory[60321] <=  8'h66;        memory[60322] <=  8'h69;        memory[60323] <=  8'h77;        memory[60324] <=  8'h68;        memory[60325] <=  8'h61;        memory[60326] <=  8'h74;        memory[60327] <=  8'h61;        memory[60328] <=  8'h6e;        memory[60329] <=  8'h61;        memory[60330] <=  8'h62;        memory[60331] <=  8'h61;        memory[60332] <=  8'h63;        memory[60333] <=  8'h61;        memory[60334] <=  8'h74;        memory[60335] <=  8'h61;        memory[60336] <=  8'h62;        memory[60337] <=  8'h61;        memory[60338] <=  8'h72;        memory[60339] <=  8'h63;        memory[60340] <=  8'h61;        memory[60341] <=  8'h68;        memory[60342] <=  8'h64;        memory[60343] <=  8'h75;        memory[60344] <=  8'h63;        memory[60345] <=  8'h74;        memory[60346] <=  8'h61;        memory[60347] <=  8'h64;        memory[60348] <=  8'h61;        memory[60349] <=  8'h61;        memory[60350] <=  8'h63;        memory[60351] <=  8'h61;        memory[60352] <=  8'h72;        memory[60353] <=  8'h63;        memory[60354] <=  8'h74;        memory[60355] <=  8'h72;        memory[60356] <=  8'h63;        memory[60357] <=  8'h61;        memory[60358] <=  8'h74;        memory[60359] <=  8'h72;        memory[60360] <=  8'h63;        memory[60361] <=  8'h61;        memory[60362] <=  8'h74;        memory[60363] <=  8'h63;        memory[60364] <=  8'h62;        memory[60365] <=  8'h61;        memory[60366] <=  8'h74;        memory[60367] <=  8'h62;        memory[60368] <=  8'h72;        memory[60369] <=  8'h63;        memory[60370] <=  8'h61;        memory[60371] <=  8'h74;        memory[60372] <=  8'h72;        memory[60373] <=  8'h6e;        memory[60374] <=  8'h62;        memory[60375] <=  8'h61;        memory[60376] <=  8'h63;        memory[60377] <=  8'h61;        memory[60378] <=  8'h74;        memory[60379] <=  8'h79;        memory[60380] <=  8'h73;        memory[60381] <=  8'h6e;        memory[60382] <=  8'h63;        memory[60383] <=  8'h74;        memory[60384] <=  8'h61;        memory[60385] <=  8'h6e;        memory[60386] <=  8'h62;        memory[60387] <=  8'h61;        memory[60388] <=  8'h63;        memory[60389] <=  8'h72;        memory[60390] <=  8'h6e;        memory[60391] <=  8'h74;        memory[60392] <=  8'h61;        memory[60393] <=  8'h62;        memory[60394] <=  8'h74;        memory[60395] <=  8'h6e;        memory[60396] <=  8'h61;        memory[60397] <=  8'h72;        memory[60398] <=  8'h62;        memory[60399] <=  8'h78;        memory[60400] <=  8'h74;        memory[60401] <=  8'h61;        memory[60402] <=  8'h72;        memory[60403] <=  8'h62;        memory[60404] <=  8'h61;        memory[60405] <=  8'h72;        memory[60406] <=  8'h74;        memory[60407] <=  8'h74;        memory[60408] <=  8'h62;        memory[60409] <=  8'h61;        memory[60410] <=  8'h72;        memory[60411] <=  8'h74;        memory[60412] <=  8'h78;        memory[60413] <=  8'h61;        memory[60414] <=  8'h74;        memory[60415] <=  8'h6b;        memory[60416] <=  8'h73;        memory[60417] <=  8'h68;        memory[60418] <=  8'h63;        memory[60419] <=  8'h66;        memory[60420] <=  8'h69;        memory[60421] <=  8'h77;        memory[60422] <=  8'h68;        memory[60423] <=  8'h61;        memory[60424] <=  8'h74;        memory[60425] <=  8'h61;        memory[60426] <=  8'h6e;        memory[60427] <=  8'h61;        memory[60428] <=  8'h62;        memory[60429] <=  8'h61;        memory[60430] <=  8'h63;        memory[60431] <=  8'h61;        memory[60432] <=  8'h74;        memory[60433] <=  8'h61;        memory[60434] <=  8'h62;        memory[60435] <=  8'h61;        memory[60436] <=  8'h72;        memory[60437] <=  8'h63;        memory[60438] <=  8'h61;        memory[60439] <=  8'h68;        memory[60440] <=  8'h64;        memory[60441] <=  8'h75;        memory[60442] <=  8'h63;        memory[60443] <=  8'h74;        memory[60444] <=  8'h61;        memory[60445] <=  8'h64;        memory[60446] <=  8'h61;        memory[60447] <=  8'h61;        memory[60448] <=  8'h63;        memory[60449] <=  8'h61;        memory[60450] <=  8'h72;        memory[60451] <=  8'h63;        memory[60452] <=  8'h74;        memory[60453] <=  8'h72;        memory[60454] <=  8'h63;        memory[60455] <=  8'h61;        memory[60456] <=  8'h74;        memory[60457] <=  8'h72;        memory[60458] <=  8'h63;        memory[60459] <=  8'h61;        memory[60460] <=  8'h74;        memory[60461] <=  8'h63;        memory[60462] <=  8'h62;        memory[60463] <=  8'h61;        memory[60464] <=  8'h74;        memory[60465] <=  8'h62;        memory[60466] <=  8'h72;        memory[60467] <=  8'h63;        memory[60468] <=  8'h61;        memory[60469] <=  8'h74;        memory[60470] <=  8'h72;        memory[60471] <=  8'h6e;        memory[60472] <=  8'h62;        memory[60473] <=  8'h61;        memory[60474] <=  8'h63;        memory[60475] <=  8'h61;        memory[60476] <=  8'h74;        memory[60477] <=  8'h79;        memory[60478] <=  8'h73;        memory[60479] <=  8'h6e;        memory[60480] <=  8'h63;        memory[60481] <=  8'h74;        memory[60482] <=  8'h61;        memory[60483] <=  8'h6e;        memory[60484] <=  8'h62;        memory[60485] <=  8'h61;        memory[60486] <=  8'h63;        memory[60487] <=  8'h72;        memory[60488] <=  8'h6e;        memory[60489] <=  8'h74;        memory[60490] <=  8'h61;        memory[60491] <=  8'h62;        memory[60492] <=  8'h74;        memory[60493] <=  8'h6e;        memory[60494] <=  8'h61;        memory[60495] <=  8'h72;        memory[60496] <=  8'h62;        memory[60497] <=  8'h78;        memory[60498] <=  8'h74;        memory[60499] <=  8'h61;        memory[60500] <=  8'h72;        memory[60501] <=  8'h5d;        memory[60502] <=  8'h5d;        memory[60503] <=  8'h65;        memory[60504] <=  8'h66;        memory[60505] <=  8'h77;        memory[60506] <=  8'h65;        memory[60507] <=  8'h5d;        memory[60508] <=  8'h65;        memory[60509] <=  8'h67;        memory[60510] <=  8'h73;        memory[60511] <=  8'h67;        memory[60512] <=  8'h66;        memory[60513] <=  8'h62;        memory[60514] <=  8'h61;        memory[60515] <=  8'h72;        memory[60516] <=  8'h74;        memory[60517] <=  8'h74;        memory[60518] <=  8'h62;        memory[60519] <=  8'h61;        memory[60520] <=  8'h72;        memory[60521] <=  8'h74;        memory[60522] <=  8'h78;        memory[60523] <=  8'h61;        memory[60524] <=  8'h74;        memory[60525] <=  8'h6b;        memory[60526] <=  8'h73;        memory[60527] <=  8'h68;        memory[60528] <=  8'h63;        memory[60529] <=  8'h66;        memory[60530] <=  8'h69;        memory[60531] <=  8'h77;        memory[60532] <=  8'h68;        memory[60533] <=  8'h61;        memory[60534] <=  8'h74;        memory[60535] <=  8'h61;        memory[60536] <=  8'h6e;        memory[60537] <=  8'h61;        memory[60538] <=  8'h62;        memory[60539] <=  8'h61;        memory[60540] <=  8'h63;        memory[60541] <=  8'h61;        memory[60542] <=  8'h74;        memory[60543] <=  8'h61;        memory[60544] <=  8'h62;        memory[60545] <=  8'h61;        memory[60546] <=  8'h72;        memory[60547] <=  8'h63;        memory[60548] <=  8'h61;        memory[60549] <=  8'h68;        memory[60550] <=  8'h64;        memory[60551] <=  8'h75;        memory[60552] <=  8'h63;        memory[60553] <=  8'h74;        memory[60554] <=  8'h61;        memory[60555] <=  8'h64;        memory[60556] <=  8'h61;        memory[60557] <=  8'h61;        memory[60558] <=  8'h63;        memory[60559] <=  8'h61;        memory[60560] <=  8'h72;        memory[60561] <=  8'h63;        memory[60562] <=  8'h74;        memory[60563] <=  8'h72;        memory[60564] <=  8'h63;        memory[60565] <=  8'h61;        memory[60566] <=  8'h74;        memory[60567] <=  8'h72;        memory[60568] <=  8'h63;        memory[60569] <=  8'h61;        memory[60570] <=  8'h74;        memory[60571] <=  8'h63;        memory[60572] <=  8'h62;        memory[60573] <=  8'h61;        memory[60574] <=  8'h74;        memory[60575] <=  8'h62;        memory[60576] <=  8'h72;        memory[60577] <=  8'h63;        memory[60578] <=  8'h61;        memory[60579] <=  8'h74;        memory[60580] <=  8'h72;        memory[60581] <=  8'h6e;        memory[60582] <=  8'h62;        memory[60583] <=  8'h61;        memory[60584] <=  8'h63;        memory[60585] <=  8'h61;        memory[60586] <=  8'h74;        memory[60587] <=  8'h79;        memory[60588] <=  8'h73;        memory[60589] <=  8'h6e;        memory[60590] <=  8'h63;        memory[60591] <=  8'h74;        memory[60592] <=  8'h61;        memory[60593] <=  8'h6e;        memory[60594] <=  8'h62;        memory[60595] <=  8'h61;        memory[60596] <=  8'h63;        memory[60597] <=  8'h72;        memory[60598] <=  8'h6e;        memory[60599] <=  8'h74;        memory[60600] <=  8'h61;        memory[60601] <=  8'h62;        memory[60602] <=  8'h74;        memory[60603] <=  8'h6e;        memory[60604] <=  8'h61;        memory[60605] <=  8'h72;        memory[60606] <=  8'h62;        memory[60607] <=  8'h78;        memory[60608] <=  8'h74;        memory[60609] <=  8'h61;        memory[60610] <=  8'h72;        memory[60611] <=  8'h62;        memory[60612] <=  8'h61;        memory[60613] <=  8'h72;        memory[60614] <=  8'h74;        memory[60615] <=  8'h74;        memory[60616] <=  8'h62;        memory[60617] <=  8'h61;        memory[60618] <=  8'h72;        memory[60619] <=  8'h74;        memory[60620] <=  8'h78;        memory[60621] <=  8'h61;        memory[60622] <=  8'h74;        memory[60623] <=  8'h6b;        memory[60624] <=  8'h73;        memory[60625] <=  8'h68;        memory[60626] <=  8'h63;        memory[60627] <=  8'h66;        memory[60628] <=  8'h69;        memory[60629] <=  8'h77;        memory[60630] <=  8'h68;        memory[60631] <=  8'h61;        memory[60632] <=  8'h74;        memory[60633] <=  8'h61;        memory[60634] <=  8'h6e;        memory[60635] <=  8'h61;        memory[60636] <=  8'h62;        memory[60637] <=  8'h61;        memory[60638] <=  8'h63;        memory[60639] <=  8'h61;        memory[60640] <=  8'h74;        memory[60641] <=  8'h61;        memory[60642] <=  8'h62;        memory[60643] <=  8'h61;        memory[60644] <=  8'h72;        memory[60645] <=  8'h63;        memory[60646] <=  8'h61;        memory[60647] <=  8'h68;        memory[60648] <=  8'h64;        memory[60649] <=  8'h75;        memory[60650] <=  8'h63;        memory[60651] <=  8'h74;        memory[60652] <=  8'h61;        memory[60653] <=  8'h64;        memory[60654] <=  8'h61;        memory[60655] <=  8'h61;        memory[60656] <=  8'h63;        memory[60657] <=  8'h61;        memory[60658] <=  8'h72;        memory[60659] <=  8'h63;        memory[60660] <=  8'h74;        memory[60661] <=  8'h72;        memory[60662] <=  8'h63;        memory[60663] <=  8'h61;        memory[60664] <=  8'h74;        memory[60665] <=  8'h72;        memory[60666] <=  8'h63;        memory[60667] <=  8'h61;        memory[60668] <=  8'h74;        memory[60669] <=  8'h63;        memory[60670] <=  8'h62;        memory[60671] <=  8'h61;        memory[60672] <=  8'h74;        memory[60673] <=  8'h62;        memory[60674] <=  8'h72;        memory[60675] <=  8'h63;        memory[60676] <=  8'h61;        memory[60677] <=  8'h74;        memory[60678] <=  8'h72;        memory[60679] <=  8'h6e;        memory[60680] <=  8'h62;        memory[60681] <=  8'h61;        memory[60682] <=  8'h63;        memory[60683] <=  8'h61;        memory[60684] <=  8'h74;        memory[60685] <=  8'h79;        memory[60686] <=  8'h73;        memory[60687] <=  8'h6e;        memory[60688] <=  8'h63;        memory[60689] <=  8'h74;        memory[60690] <=  8'h61;        memory[60691] <=  8'h6e;        memory[60692] <=  8'h62;        memory[60693] <=  8'h61;        memory[60694] <=  8'h63;        memory[60695] <=  8'h72;        memory[60696] <=  8'h6e;        memory[60697] <=  8'h74;        memory[60698] <=  8'h61;        memory[60699] <=  8'h62;        memory[60700] <=  8'h74;        memory[60701] <=  8'h6e;        memory[60702] <=  8'h61;        memory[60703] <=  8'h72;        memory[60704] <=  8'h62;        memory[60705] <=  8'h78;        memory[60706] <=  8'h74;        memory[60707] <=  8'h61;        memory[60708] <=  8'h72;        memory[60709] <=  8'h64;        memory[60710] <=  8'h66;        memory[60711] <=  8'h73;        memory[60712] <=  8'h67;        memory[60713] <=  8'h76;        memory[60714] <=  8'h68;        memory[60715] <=  8'h62;        memory[60716] <=  8'h6b;        memory[60717] <=  8'h6a;        memory[60718] <=  8'h6e;        memory[60719] <=  8'h6d;        memory[60720] <=  8'h62;        memory[60721] <=  8'h76;        memory[60722] <=  8'h78;        memory[60723] <=  8'h63;        memory[60724] <=  8'h73;        memory[60725] <=  8'h66;        memory[60726] <=  8'h72;        memory[60727] <=  8'h74;        memory[60728] <=  8'h79;        memory[60729] <=  8'h75;        memory[60730] <=  8'h6a;        memory[60731] <=  8'h6e;        memory[60732] <=  8'h62;        memory[60733] <=  8'h76;        memory[60734] <=  8'h63;        memory[60735] <=  8'h64;        memory[60736] <=  8'h74;        memory[60737] <=  8'h79;        memory[60738] <=  8'h75;        memory[60739] <=  8'h69;        memory[60740] <=  8'h6b;        memory[60741] <=  8'h6d;        memory[60742] <=  8'h6e;        memory[60743] <=  8'h62;        memory[60744] <=  8'h76;        memory[60745] <=  8'h63;        memory[60746] <=  8'h78;        memory[60747] <=  8'h73;        memory[60748] <=  8'h64;        memory[60749] <=  8'h72;        memory[60750] <=  8'h74;        memory[60751] <=  8'h79;        memory[60752] <=  8'h75;        memory[60753] <=  8'h69;        memory[60754] <=  8'h6b;        memory[60755] <=  8'h6d;        memory[60756] <=  8'h6e;        memory[60757] <=  8'h62;        memory[60758] <=  8'h76;        memory[60759] <=  8'h63;        memory[60760] <=  8'h73;        memory[60761] <=  8'h77;        memory[60762] <=  8'h33;        memory[60763] <=  8'h34;        memory[60764] <=  8'h35;        memory[60765] <=  8'h36;        memory[60766] <=  8'h37;        memory[60767] <=  8'h38;        memory[60768] <=  8'h69;        memory[60769] <=  8'h6b;        memory[60770] <=  8'h6d;        memory[60771] <=  8'h6e;        memory[60772] <=  8'h62;        memory[60773] <=  8'h76;        memory[60774] <=  8'h63;        memory[60775] <=  8'h64;        memory[60776] <=  8'h65;        memory[60777] <=  8'h72;        memory[60778] <=  8'h36;        memory[60779] <=  8'h37;        memory[60780] <=  8'h38;        memory[60781] <=  8'h69;        memory[60782] <=  8'h6f;        memory[60783] <=  8'h6b;        memory[60784] <=  8'h6a;        memory[60785] <=  8'h6e;        memory[60786] <=  8'h62;        memory[60787] <=  8'h76;        memory[60788] <=  8'h63;        memory[60789] <=  8'h64;        memory[60790] <=  8'h72;        memory[60791] <=  8'h74;        memory[60792] <=  8'h79;        memory[60793] <=  8'h75;        memory[60794] <=  8'h73;        memory[60795] <=  8'h6a;        memory[60796] <=  8'h63;        memory[60797] <=  8'h6e;        memory[60798] <=  8'h62;        memory[60799] <=  8'h64;        memory[60800] <=  8'h66;        memory[60801] <=  8'h73;        memory[60802] <=  8'h74;        memory[60803] <=  8'h79;        memory[60804] <=  8'h75;        memory[60805] <=  8'h61;        memory[60806] <=  8'h69;        memory[60807] <=  8'h6b;        memory[60808] <=  8'h78;        memory[60809] <=  8'h6d;        memory[60810] <=  8'h6e;        memory[60811] <=  8'h73;        memory[60812] <=  8'h6a;        memory[60813] <=  8'h6f;        memory[60814] <=  8'h64;        memory[60815] <=  8'h6c;        memory[60816] <=  8'h63;        memory[60817] <=  8'h78;        memory[60818] <=  8'h62;        memory[60819] <=  8'h61;        memory[60820] <=  8'h72;        memory[60821] <=  8'h74;        memory[60822] <=  8'h78;        memory[60823] <=  8'h61;        memory[60824] <=  8'h74;        memory[60825] <=  8'h6b;        memory[60826] <=  8'h73;        memory[60827] <=  8'h68;        memory[60828] <=  8'h63;        memory[60829] <=  8'h66;        memory[60830] <=  8'h69;        memory[60831] <=  8'h77;        memory[60832] <=  8'h68;        memory[60833] <=  8'h61;        memory[60834] <=  8'h74;        memory[60835] <=  8'h61;        memory[60836] <=  8'h6e;        memory[60837] <=  8'h61;        memory[60838] <=  8'h62;        memory[60839] <=  8'h61;        memory[60840] <=  8'h63;        memory[60841] <=  8'h61;        memory[60842] <=  8'h74;        memory[60843] <=  8'h61;        memory[60844] <=  8'h62;        memory[60845] <=  8'h61;        memory[60846] <=  8'h72;        memory[60847] <=  8'h63;        memory[60848] <=  8'h61;        memory[60849] <=  8'h68;        memory[60850] <=  8'h64;        memory[60851] <=  8'h75;        memory[60852] <=  8'h63;        memory[60853] <=  8'h74;        memory[60854] <=  8'h61;        memory[60855] <=  8'h64;        memory[60856] <=  8'h61;        memory[60857] <=  8'h61;        memory[60858] <=  8'h63;        memory[60859] <=  8'h61;        memory[60860] <=  8'h72;        memory[60861] <=  8'h62;        memory[60862] <=  8'h61;        memory[60863] <=  8'h72;        memory[60864] <=  8'h74;        memory[60865] <=  8'h78;        memory[60866] <=  8'h61;        memory[60867] <=  8'h74;        memory[60868] <=  8'h6b;        memory[60869] <=  8'h73;        memory[60870] <=  8'h68;        memory[60871] <=  8'h63;        memory[60872] <=  8'h66;        memory[60873] <=  8'h69;        memory[60874] <=  8'h77;        memory[60875] <=  8'h68;        memory[60876] <=  8'h61;        memory[60877] <=  8'h74;        memory[60878] <=  8'h61;        memory[60879] <=  8'h6e;        memory[60880] <=  8'h61;        memory[60881] <=  8'h62;        memory[60882] <=  8'h61;        memory[60883] <=  8'h63;        memory[60884] <=  8'h61;        memory[60885] <=  8'h74;        memory[60886] <=  8'h61;        memory[60887] <=  8'h62;        memory[60888] <=  8'h61;        memory[60889] <=  8'h72;        memory[60890] <=  8'h63;        memory[60891] <=  8'h61;        memory[60892] <=  8'h68;        memory[60893] <=  8'h64;        memory[60894] <=  8'h75;        memory[60895] <=  8'h63;        memory[60896] <=  8'h74;        memory[60897] <=  8'h61;        memory[60898] <=  8'h64;        memory[60899] <=  8'h61;        memory[60900] <=  8'h61;        memory[60901] <=  8'h63;        memory[60902] <=  8'h61;        memory[60903] <=  8'h72;        memory[60904] <=  8'h62;        memory[60905] <=  8'h61;        memory[60906] <=  8'h72;        memory[60907] <=  8'h74;        memory[60908] <=  8'h78;        memory[60909] <=  8'h61;        memory[60910] <=  8'h74;        memory[60911] <=  8'h6b;        memory[60912] <=  8'h73;        memory[60913] <=  8'h68;        memory[60914] <=  8'h63;        memory[60915] <=  8'h66;        memory[60916] <=  8'h69;        memory[60917] <=  8'h77;        memory[60918] <=  8'h68;        memory[60919] <=  8'h61;        memory[60920] <=  8'h74;        memory[60921] <=  8'h61;        memory[60922] <=  8'h6e;        memory[60923] <=  8'h61;        memory[60924] <=  8'h62;        memory[60925] <=  8'h61;        memory[60926] <=  8'h63;        memory[60927] <=  8'h61;        memory[60928] <=  8'h74;        memory[60929] <=  8'h61;        memory[60930] <=  8'h62;        memory[60931] <=  8'h61;        memory[60932] <=  8'h72;        memory[60933] <=  8'h63;        memory[60934] <=  8'h61;        memory[60935] <=  8'h68;        memory[60936] <=  8'h64;        memory[60937] <=  8'h75;        memory[60938] <=  8'h63;        memory[60939] <=  8'h74;        memory[60940] <=  8'h61;        memory[60941] <=  8'h64;        memory[60942] <=  8'h61;        memory[60943] <=  8'h61;        memory[60944] <=  8'h63;        memory[60945] <=  8'h61;        memory[60946] <=  8'h72;        memory[60947] <=  8'h62;        memory[60948] <=  8'h61;        memory[60949] <=  8'h72;        memory[60950] <=  8'h74;        memory[60951] <=  8'h78;        memory[60952] <=  8'h61;        memory[60953] <=  8'h74;        memory[60954] <=  8'h6b;        memory[60955] <=  8'h73;        memory[60956] <=  8'h68;        memory[60957] <=  8'h63;        memory[60958] <=  8'h66;        memory[60959] <=  8'h69;        memory[60960] <=  8'h77;        memory[60961] <=  8'h68;        memory[60962] <=  8'h61;        memory[60963] <=  8'h74;        memory[60964] <=  8'h61;        memory[60965] <=  8'h6e;        memory[60966] <=  8'h61;        memory[60967] <=  8'h62;        memory[60968] <=  8'h61;        memory[60969] <=  8'h63;        memory[60970] <=  8'h61;        memory[60971] <=  8'h74;        memory[60972] <=  8'h61;        memory[60973] <=  8'h62;        memory[60974] <=  8'h61;        memory[60975] <=  8'h72;        memory[60976] <=  8'h63;        memory[60977] <=  8'h61;        memory[60978] <=  8'h68;        memory[60979] <=  8'h64;        memory[60980] <=  8'h75;        memory[60981] <=  8'h63;        memory[60982] <=  8'h74;        memory[60983] <=  8'h61;        memory[60984] <=  8'h64;        memory[60985] <=  8'h61;        memory[60986] <=  8'h61;        memory[60987] <=  8'h63;        memory[60988] <=  8'h61;        memory[60989] <=  8'h72;        memory[60990] <=  8'h62;        memory[60991] <=  8'h61;        memory[60992] <=  8'h72;        memory[60993] <=  8'h74;        memory[60994] <=  8'h78;        memory[60995] <=  8'h61;        memory[60996] <=  8'h74;        memory[60997] <=  8'h6b;        memory[60998] <=  8'h73;        memory[60999] <=  8'h68;        memory[61000] <=  8'h63;        memory[61001] <=  8'h66;        memory[61002] <=  8'h69;        memory[61003] <=  8'h77;        memory[61004] <=  8'h68;        memory[61005] <=  8'h61;        memory[61006] <=  8'h74;        memory[61007] <=  8'h61;        memory[61008] <=  8'h6e;        memory[61009] <=  8'h61;        memory[61010] <=  8'h62;        memory[61011] <=  8'h61;        memory[61012] <=  8'h63;        memory[61013] <=  8'h61;        memory[61014] <=  8'h74;        memory[61015] <=  8'h61;        memory[61016] <=  8'h62;        memory[61017] <=  8'h61;        memory[61018] <=  8'h72;        memory[61019] <=  8'h63;        memory[61020] <=  8'h61;        memory[61021] <=  8'h68;        memory[61022] <=  8'h64;        memory[61023] <=  8'h75;        memory[61024] <=  8'h63;        memory[61025] <=  8'h74;        memory[61026] <=  8'h61;        memory[61027] <=  8'h64;        memory[61028] <=  8'h61;        memory[61029] <=  8'h61;        memory[61030] <=  8'h63;        memory[61031] <=  8'h61;        memory[61032] <=  8'h72;        memory[61033] <=  8'h62;        memory[61034] <=  8'h61;        memory[61035] <=  8'h72;        memory[61036] <=  8'h74;        memory[61037] <=  8'h78;        memory[61038] <=  8'h61;        memory[61039] <=  8'h74;        memory[61040] <=  8'h6b;        memory[61041] <=  8'h73;        memory[61042] <=  8'h68;        memory[61043] <=  8'h63;        memory[61044] <=  8'h66;        memory[61045] <=  8'h69;        memory[61046] <=  8'h77;        memory[61047] <=  8'h68;        memory[61048] <=  8'h61;        memory[61049] <=  8'h74;        memory[61050] <=  8'h61;        memory[61051] <=  8'h6e;        memory[61052] <=  8'h61;        memory[61053] <=  8'h62;        memory[61054] <=  8'h61;        memory[61055] <=  8'h63;        memory[61056] <=  8'h61;        memory[61057] <=  8'h74;        memory[61058] <=  8'h61;        memory[61059] <=  8'h62;        memory[61060] <=  8'h61;        memory[61061] <=  8'h72;        memory[61062] <=  8'h63;        memory[61063] <=  8'h61;        memory[61064] <=  8'h68;        memory[61065] <=  8'h64;        memory[61066] <=  8'h75;        memory[61067] <=  8'h63;        memory[61068] <=  8'h74;        memory[61069] <=  8'h61;        memory[61070] <=  8'h64;        memory[61071] <=  8'h61;        memory[61072] <=  8'h61;        memory[61073] <=  8'h63;        memory[61074] <=  8'h61;        memory[61075] <=  8'h72;        memory[61076] <=  8'h62;        memory[61077] <=  8'h61;        memory[61078] <=  8'h72;        memory[61079] <=  8'h74;        memory[61080] <=  8'h78;        memory[61081] <=  8'h61;        memory[61082] <=  8'h74;        memory[61083] <=  8'h6b;        memory[61084] <=  8'h73;        memory[61085] <=  8'h68;        memory[61086] <=  8'h63;        memory[61087] <=  8'h66;        memory[61088] <=  8'h69;        memory[61089] <=  8'h77;        memory[61090] <=  8'h68;        memory[61091] <=  8'h61;        memory[61092] <=  8'h74;        memory[61093] <=  8'h61;        memory[61094] <=  8'h6e;        memory[61095] <=  8'h61;        memory[61096] <=  8'h62;        memory[61097] <=  8'h61;        memory[61098] <=  8'h63;        memory[61099] <=  8'h61;        memory[61100] <=  8'h74;        memory[61101] <=  8'h61;        memory[61102] <=  8'h62;        memory[61103] <=  8'h61;        memory[61104] <=  8'h72;        memory[61105] <=  8'h63;        memory[61106] <=  8'h61;        memory[61107] <=  8'h68;        memory[61108] <=  8'h64;        memory[61109] <=  8'h75;        memory[61110] <=  8'h63;        memory[61111] <=  8'h74;        memory[61112] <=  8'h61;        memory[61113] <=  8'h64;        memory[61114] <=  8'h61;        memory[61115] <=  8'h61;        memory[61116] <=  8'h63;        memory[61117] <=  8'h61;        memory[61118] <=  8'h72;        memory[61119] <=  8'h62;        memory[61120] <=  8'h61;        memory[61121] <=  8'h72;        memory[61122] <=  8'h74;        memory[61123] <=  8'h78;        memory[61124] <=  8'h61;        memory[61125] <=  8'h74;        memory[61126] <=  8'h6b;        memory[61127] <=  8'h73;        memory[61128] <=  8'h68;        memory[61129] <=  8'h63;        memory[61130] <=  8'h66;        memory[61131] <=  8'h69;        memory[61132] <=  8'h77;        memory[61133] <=  8'h68;        memory[61134] <=  8'h61;        memory[61135] <=  8'h74;        memory[61136] <=  8'h61;        memory[61137] <=  8'h6e;        memory[61138] <=  8'h61;        memory[61139] <=  8'h62;        memory[61140] <=  8'h61;        memory[61141] <=  8'h63;        memory[61142] <=  8'h61;        memory[61143] <=  8'h74;        memory[61144] <=  8'h61;        memory[61145] <=  8'h62;        memory[61146] <=  8'h61;        memory[61147] <=  8'h72;        memory[61148] <=  8'h63;        memory[61149] <=  8'h61;        memory[61150] <=  8'h68;        memory[61151] <=  8'h64;        memory[61152] <=  8'h75;        memory[61153] <=  8'h63;        memory[61154] <=  8'h74;        memory[61155] <=  8'h61;        memory[61156] <=  8'h64;        memory[61157] <=  8'h61;        memory[61158] <=  8'h61;        memory[61159] <=  8'h63;        memory[61160] <=  8'h61;        memory[61161] <=  8'h72;        memory[61162] <=  8'h62;        memory[61163] <=  8'h61;        memory[61164] <=  8'h72;        memory[61165] <=  8'h74;        memory[61166] <=  8'h78;        memory[61167] <=  8'h61;        memory[61168] <=  8'h74;        memory[61169] <=  8'h6b;        memory[61170] <=  8'h73;        memory[61171] <=  8'h68;        memory[61172] <=  8'h63;        memory[61173] <=  8'h66;        memory[61174] <=  8'h69;        memory[61175] <=  8'h77;        memory[61176] <=  8'h68;        memory[61177] <=  8'h61;        memory[61178] <=  8'h74;        memory[61179] <=  8'h61;        memory[61180] <=  8'h6e;        memory[61181] <=  8'h61;        memory[61182] <=  8'h62;        memory[61183] <=  8'h61;        memory[61184] <=  8'h63;        memory[61185] <=  8'h61;        memory[61186] <=  8'h74;        memory[61187] <=  8'h61;        memory[61188] <=  8'h62;        memory[61189] <=  8'h61;        memory[61190] <=  8'h72;        memory[61191] <=  8'h63;        memory[61192] <=  8'h61;        memory[61193] <=  8'h68;        memory[61194] <=  8'h64;        memory[61195] <=  8'h75;        memory[61196] <=  8'h63;        memory[61197] <=  8'h74;        memory[61198] <=  8'h61;        memory[61199] <=  8'h64;        memory[61200] <=  8'h61;        memory[61201] <=  8'h61;        memory[61202] <=  8'h63;        memory[61203] <=  8'h61;        memory[61204] <=  8'h72;        memory[61205] <=  8'h62;        memory[61206] <=  8'h61;        memory[61207] <=  8'h72;        memory[61208] <=  8'h74;        memory[61209] <=  8'h74;        memory[61210] <=  8'h62;        memory[61211] <=  8'h61;        memory[61212] <=  8'h72;        memory[61213] <=  8'h74;        memory[61214] <=  8'h78;        memory[61215] <=  8'h61;        memory[61216] <=  8'h74;        memory[61217] <=  8'h6b;        memory[61218] <=  8'h73;        memory[61219] <=  8'h68;        memory[61220] <=  8'h63;        memory[61221] <=  8'h66;        memory[61222] <=  8'h69;        memory[61223] <=  8'h77;        memory[61224] <=  8'h68;        memory[61225] <=  8'h61;        memory[61226] <=  8'h74;        memory[61227] <=  8'h61;        memory[61228] <=  8'h6e;        memory[61229] <=  8'h61;        memory[61230] <=  8'h62;        memory[61231] <=  8'h61;        memory[61232] <=  8'h63;        memory[61233] <=  8'h61;        memory[61234] <=  8'h74;        memory[61235] <=  8'h61;        memory[61236] <=  8'h62;        memory[61237] <=  8'h61;        memory[61238] <=  8'h72;        memory[61239] <=  8'h63;        memory[61240] <=  8'h61;        memory[61241] <=  8'h68;        memory[61242] <=  8'h64;        memory[61243] <=  8'h75;        memory[61244] <=  8'h63;        memory[61245] <=  8'h74;        memory[61246] <=  8'h61;        memory[61247] <=  8'h64;        memory[61248] <=  8'h61;        memory[61249] <=  8'h61;        memory[61250] <=  8'h63;        memory[61251] <=  8'h61;        memory[61252] <=  8'h72;        memory[61253] <=  8'h63;        memory[61254] <=  8'h74;        memory[61255] <=  8'h72;        memory[61256] <=  8'h63;        memory[61257] <=  8'h61;        memory[61258] <=  8'h74;        memory[61259] <=  8'h72;        memory[61260] <=  8'h63;        memory[61261] <=  8'h61;        memory[61262] <=  8'h74;        memory[61263] <=  8'h63;        memory[61264] <=  8'h62;        memory[61265] <=  8'h61;        memory[61266] <=  8'h74;        memory[61267] <=  8'h62;        memory[61268] <=  8'h72;        memory[61269] <=  8'h63;        memory[61270] <=  8'h61;        memory[61271] <=  8'h72;        memory[61272] <=  8'h62;        memory[61273] <=  8'h78;        memory[61274] <=  8'h74;        memory[61275] <=  8'h61;        memory[61276] <=  8'h72;        memory[61277] <=  8'h64;        memory[61278] <=  8'h66;        memory[61279] <=  8'h73;        memory[61280] <=  8'h67;        memory[61281] <=  8'h76;        memory[61282] <=  8'h68;        memory[61283] <=  8'h62;        memory[61284] <=  8'h6b;        memory[61285] <=  8'h6a;        memory[61286] <=  8'h6e;        memory[61287] <=  8'h6d;        memory[61288] <=  8'h62;        memory[61289] <=  8'h76;        memory[61290] <=  8'h78;        memory[61291] <=  8'h63;        memory[61292] <=  8'h73;        memory[61293] <=  8'h66;        memory[61294] <=  8'h72;        memory[61295] <=  8'h74;        memory[61296] <=  8'h79;        memory[61297] <=  8'h75;        memory[61298] <=  8'h6a;        memory[61299] <=  8'h6e;        memory[61300] <=  8'h62;        memory[61301] <=  8'h76;        memory[61302] <=  8'h63;        memory[61303] <=  8'h64;        memory[61304] <=  8'h74;        memory[61305] <=  8'h79;        memory[61306] <=  8'h75;        memory[61307] <=  8'h69;        memory[61308] <=  8'h6b;        memory[61309] <=  8'h6d;        memory[61310] <=  8'h6e;        memory[61311] <=  8'h62;        memory[61312] <=  8'h76;        memory[61313] <=  8'h63;        memory[61314] <=  8'h78;        memory[61315] <=  8'h73;        memory[61316] <=  8'h64;        memory[61317] <=  8'h72;        memory[61318] <=  8'h74;        memory[61319] <=  8'h79;        memory[61320] <=  8'h75;        memory[61321] <=  8'h69;        memory[61322] <=  8'h6b;        memory[61323] <=  8'h6d;        memory[61324] <=  8'h6e;        memory[61325] <=  8'h62;        memory[61326] <=  8'h76;        memory[61327] <=  8'h63;        memory[61328] <=  8'h73;        memory[61329] <=  8'h77;        memory[61330] <=  8'h33;        memory[61331] <=  8'h34;        memory[61332] <=  8'h35;        memory[61333] <=  8'h36;        memory[61334] <=  8'h37;        memory[61335] <=  8'h38;        memory[61336] <=  8'h69;        memory[61337] <=  8'h6b;        memory[61338] <=  8'h6d;        memory[61339] <=  8'h6e;        memory[61340] <=  8'h62;        memory[61341] <=  8'h76;        memory[61342] <=  8'h63;        memory[61343] <=  8'h64;        memory[61344] <=  8'h65;        memory[61345] <=  8'h72;        memory[61346] <=  8'h36;        memory[61347] <=  8'h37;        memory[61348] <=  8'h38;        memory[61349] <=  8'h69;        memory[61350] <=  8'h6f;        memory[61351] <=  8'h6b;        memory[61352] <=  8'h6a;        memory[61353] <=  8'h6e;        memory[61354] <=  8'h62;        memory[61355] <=  8'h76;        memory[61356] <=  8'h63;        memory[61357] <=  8'h64;        memory[61358] <=  8'h72;        memory[61359] <=  8'h74;        memory[61360] <=  8'h79;        memory[61361] <=  8'h75;        memory[61362] <=  8'h73;        memory[61363] <=  8'h6a;        memory[61364] <=  8'h63;        memory[61365] <=  8'h6e;        memory[61366] <=  8'h62;        memory[61367] <=  8'h64;        memory[61368] <=  8'h66;        memory[61369] <=  8'h73;        memory[61370] <=  8'h74;        memory[61371] <=  8'h79;        memory[61372] <=  8'h75;        memory[61373] <=  8'h61;        memory[61374] <=  8'h69;        memory[61375] <=  8'h6b;        memory[61376] <=  8'h78;        memory[61377] <=  8'h6d;        memory[61378] <=  8'h6e;        memory[61379] <=  8'h73;        memory[61380] <=  8'h6a;        memory[61381] <=  8'h6f;        memory[61382] <=  8'h64;        memory[61383] <=  8'h6c;        memory[61384] <=  8'h63;        memory[61385] <=  8'h78;        memory[61386] <=  8'h2c;        memory[61387] <=  8'h6d;        memory[61388] <=  8'h73;        memory[61389] <=  8'h6b;        memory[61390] <=  8'h64;        memory[61391] <=  8'h6c;        memory[61392] <=  8'h70;        memory[61393] <=  8'h5b;        memory[61394] <=  8'h3b;        memory[61395] <=  8'h73;        memory[61396] <=  8'h6c;        memory[61397] <=  8'h64;        memory[61398] <=  8'h70;        memory[61399] <=  8'h76;        memory[61400] <=  8'h63;        memory[61401] <=  8'h5b;        memory[61402] <=  8'h78;        memory[61403] <=  8'h76;        memory[61404] <=  8'h63;        memory[61405] <=  8'h5b;        memory[61406] <=  8'h78;        memory[61407] <=  8'h70;        memory[61408] <=  8'h6f;        memory[61409] <=  8'h20;        memory[61410] <=  8'h62;        memory[61411] <=  8'h61;        memory[61412] <=  8'h72;        memory[61413] <=  8'h74;        memory[61414] <=  8'h74;        memory[61415] <=  8'h62;        memory[61416] <=  8'h61;        memory[61417] <=  8'h72;        memory[61418] <=  8'h74;        memory[61419] <=  8'h78;        memory[61420] <=  8'h61;        memory[61421] <=  8'h74;        memory[61422] <=  8'h6b;        memory[61423] <=  8'h73;        memory[61424] <=  8'h68;        memory[61425] <=  8'h63;        memory[61426] <=  8'h66;        memory[61427] <=  8'h69;        memory[61428] <=  8'h77;        memory[61429] <=  8'h68;        memory[61430] <=  8'h61;        memory[61431] <=  8'h69;        memory[61432] <=  8'h6a;        memory[61433] <=  8'h78;        memory[61434] <=  8'h5d;        memory[61435] <=  8'h65;        memory[61436] <=  8'h6b;        memory[61437] <=  8'h6f;        memory[61438] <=  8'h39;        memory[61439] <=  8'h64;        memory[61440] <=  8'h75;        memory[61441] <=  8'h38;        memory[61442] <=  8'h79;        memory[61443] <=  8'h20;        memory[61444] <=  8'h37;        memory[61445] <=  8'h63;        memory[61446] <=  8'h67;        memory[61447] <=  8'h78;        memory[61448] <=  8'h63;        memory[61449] <=  8'h75;        memory[61450] <=  8'h68;        memory[61451] <=  8'h69;        memory[61452] <=  8'h6a;        memory[61453] <=  8'h77;        memory[61454] <=  8'h69;        memory[61455] <=  8'h64;        memory[61456] <=  8'h66;        memory[61457] <=  8'h68;        memory[61458] <=  8'h75;        memory[61459] <=  8'h76;        memory[61460] <=  8'h64;        memory[61461] <=  8'h62;        memory[61462] <=  8'h66;        memory[61463] <=  8'h6a;        memory[61464] <=  8'h6e;        memory[61465] <=  8'h6b;        memory[61466] <=  8'h6a;        memory[61467] <=  8'h65;        memory[61468] <=  8'h38;        memory[61469] <=  8'h66;        memory[61470] <=  8'h37;        memory[61471] <=  8'h67;        memory[61472] <=  8'h79;        memory[61473] <=  8'h76;        memory[61474] <=  8'h63;        memory[61475] <=  8'h68;        memory[61476] <=  8'h69;        memory[61477] <=  8'h6a;        memory[61478] <=  8'h33;        memory[61479] <=  8'h65;        memory[61480] <=  8'h67;        memory[61481] <=  8'h79;        memory[61482] <=  8'h72;        memory[61483] <=  8'h64;        memory[61484] <=  8'h62;        memory[61485] <=  8'h6e;        memory[61486] <=  8'h63;        memory[61487] <=  8'h7a;        memory[61488] <=  8'h6a;        memory[61489] <=  8'h6f;        memory[61490] <=  8'h66;        memory[61491] <=  8'h78;        memory[61492] <=  8'h6a;        memory[61493] <=  8'h69;        memory[61494] <=  8'h63;        memory[61495] <=  8'h68;        memory[61496] <=  8'h62;        memory[61497] <=  8'h6e;        memory[61498] <=  8'h6d;        memory[61499] <=  8'h63;        memory[61500] <=  8'h73;        memory[61501] <=  8'h6c;        memory[61502] <=  8'h6b;        memory[61503] <=  8'h6a;        memory[61504] <=  8'h69;        memory[61505] <=  8'h68;        memory[61506] <=  8'h76;        memory[61507] <=  8'h75;        memory[61508] <=  8'h69;        memory[61509] <=  8'h64;        memory[61510] <=  8'h68;        memory[61511] <=  8'h75;        memory[61512] <=  8'h67;        memory[61513] <=  8'h79;        memory[61514] <=  8'h62;        memory[61515] <=  8'h68;        memory[61516] <=  8'h65;        memory[61517] <=  8'h6a;        memory[61518] <=  8'h72;        memory[61519] <=  8'h6b;        memory[61520] <=  8'h6a;        memory[61521] <=  8'h6f;        memory[61522] <=  8'h64;        memory[61523] <=  8'h67;        memory[61524] <=  8'h69;        memory[61525] <=  8'h75;        memory[61526] <=  8'h69;        memory[61527] <=  8'h67;        memory[61528] <=  8'h76;        memory[61529] <=  8'h79;        memory[61530] <=  8'h75;        memory[61531] <=  8'h67;        memory[61532] <=  8'h78;        memory[61533] <=  8'h68;        memory[61534] <=  8'h63;        memory[61535] <=  8'h20;        memory[61536] <=  8'h20;        memory[61537] <=  8'h20;        memory[61538] <=  8'h78;        memory[61539] <=  8'h76;        memory[61540] <=  8'h20;        memory[61541] <=  8'h63;        memory[61542] <=  8'h78;        memory[61543] <=  8'h67;        memory[61544] <=  8'h79;        memory[61545] <=  8'h63;        memory[61546] <=  8'h75;        memory[61547] <=  8'h68;        memory[61548] <=  8'h6a;        memory[61549] <=  8'h6b;        memory[61550] <=  8'h61;        memory[61551] <=  8'h6c;        memory[61552] <=  8'h78;        memory[61553] <=  8'h76;        memory[61554] <=  8'h70;        memory[61555] <=  8'h6f;        memory[61556] <=  8'h69;        memory[61557] <=  8'h6a;        memory[61558] <=  8'h69;        memory[61559] <=  8'h68;        memory[61560] <=  8'h6a;        memory[61561] <=  8'h62;        memory[61562] <=  8'h77;        memory[61563] <=  8'h65;        memory[61564] <=  8'h6e;        memory[61565] <=  8'h61;        memory[61566] <=  8'h66;        memory[61567] <=  8'h6d;        memory[61568] <=  8'h64;        memory[61569] <=  8'h6b;        memory[61570] <=  8'h6d;        memory[61571] <=  8'h76;        memory[61572] <=  8'h6c;        memory[61573] <=  8'h63;        memory[61574] <=  8'h6f;        memory[61575] <=  8'h64;        memory[61576] <=  8'h69;        memory[61577] <=  8'h75;        memory[61578] <=  8'h68;        memory[61579] <=  8'h73;        memory[61580] <=  8'h66;        memory[61581] <=  8'h65;        memory[61582] <=  8'h62;        memory[61583] <=  8'h6e;        memory[61584] <=  8'h64;        memory[61585] <=  8'h73;        memory[61586] <=  8'h63;        memory[61587] <=  8'h6b;        memory[61588] <=  8'h20;        memory[61589] <=  8'h78;        memory[61590] <=  8'h6a;        memory[61591] <=  8'h78;        memory[61592] <=  8'h63;        memory[61593] <=  8'h73;        memory[61594] <=  8'h64;        memory[61595] <=  8'h66;        memory[61596] <=  8'h6b;        memory[61597] <=  8'h64;        memory[61598] <=  8'h6e;        memory[61599] <=  8'h6d;        memory[61600] <=  8'h64;        memory[61601] <=  8'h73;        memory[61602] <=  8'h63;        memory[61603] <=  8'h6b;        memory[61604] <=  8'h78;        memory[61605] <=  8'h6c;        memory[61606] <=  8'h6f;        memory[61607] <=  8'h66;        memory[61608] <=  8'h6a;        memory[61609] <=  8'h69;        memory[61610] <=  8'h61;        memory[61611] <=  8'h62;        memory[61612] <=  8'h6e;        memory[61613] <=  8'h20;        memory[61614] <=  8'h78;        memory[61615] <=  8'h6b;        memory[61616] <=  8'h6d;        memory[61617] <=  8'h20;        memory[61618] <=  8'h6f;        memory[61619] <=  8'h63;        memory[61620] <=  8'h76;        memory[61621] <=  8'h73;        memory[61622] <=  8'h64;        memory[61623] <=  8'h69;        memory[61624] <=  8'h66;        memory[61625] <=  8'h68;        memory[61626] <=  8'h65;        memory[61627] <=  8'h71;        memory[61628] <=  8'h6a;        memory[61629] <=  8'h77;        memory[61630] <=  8'h62;        memory[61631] <=  8'h65;        memory[61632] <=  8'h6e;        memory[61633] <=  8'h20;        memory[61634] <=  8'h6d;        memory[61635] <=  8'h64;        memory[61636] <=  8'h73;        memory[61637] <=  8'h6c;        memory[61638] <=  8'h76;        memory[61639] <=  8'h6b;        memory[61640] <=  8'h63;        memory[61641] <=  8'h78;        memory[61642] <=  8'h20;        memory[61643] <=  8'h6f;        memory[61644] <=  8'h78;        memory[61645] <=  8'h69;        memory[61646] <=  8'h63;        memory[61647] <=  8'h6a;        memory[61648] <=  8'h76;        memory[61649] <=  8'h64;        memory[61650] <=  8'h66;        memory[61651] <=  8'h65;        memory[61652] <=  8'h71;        memory[61653] <=  8'h6e;        memory[61654] <=  8'h20;        memory[61655] <=  8'h64;        memory[61656] <=  8'h6d;        memory[61657] <=  8'h73;        memory[61658] <=  8'h6c;        memory[61659] <=  8'h63;        memory[61660] <=  8'h78;        memory[61661] <=  8'h6b;        memory[61662] <=  8'h20;        memory[61663] <=  8'h6f;        memory[61664] <=  8'h78;        memory[61665] <=  8'h63;        memory[61666] <=  8'h76;        memory[61667] <=  8'h6a;        memory[61668] <=  8'h64;        memory[61669] <=  8'h62;        memory[61670] <=  8'h71;        memory[61671] <=  8'h77;        memory[61672] <=  8'h65;        memory[61673] <=  8'h6e;        memory[61674] <=  8'h6d;        memory[61675] <=  8'h64;        memory[61676] <=  8'h6c;        memory[61677] <=  8'h73;        memory[61678] <=  8'h2c;        memory[61679] <=  8'h76;        memory[61680] <=  8'h63;        memory[61681] <=  8'h78;        memory[61682] <=  8'h20;        memory[61683] <=  8'h63;        memory[61684] <=  8'h6f;        memory[61685] <=  8'h69;        memory[61686] <=  8'h76;        memory[61687] <=  8'h68;        memory[61688] <=  8'h73;        memory[61689] <=  8'h64;        memory[61690] <=  8'h62;        memory[61691] <=  8'h71;        memory[61692] <=  8'h77;        memory[61693] <=  8'h65;        memory[61694] <=  8'h6e;        memory[61695] <=  8'h64;        memory[61696] <=  8'h6b;        memory[61697] <=  8'h73;        memory[61698] <=  8'h76;        memory[61699] <=  8'h6f;        memory[61700] <=  8'h63;        memory[61701] <=  8'h20;        memory[61702] <=  8'h76;        memory[61703] <=  8'h69;        memory[61704] <=  8'h75;        memory[61705] <=  8'h69;        memory[61706] <=  8'h68;        memory[61707] <=  8'h63;        memory[61708] <=  8'h78;        memory[61709] <=  8'h69;        memory[61710] <=  8'h6f;        memory[61711] <=  8'h76;        memory[61712] <=  8'h73;        memory[61713] <=  8'h64;        memory[61714] <=  8'h61;        memory[61715] <=  8'h64;        memory[61716] <=  8'h6e;        memory[61717] <=  8'h77;        memory[61718] <=  8'h71;        memory[61719] <=  8'h6b;        memory[61720] <=  8'h6c;        memory[61721] <=  8'h73;        memory[61722] <=  8'h76;        memory[61723] <=  8'h6e;        memory[61724] <=  8'h62;        memory[61725] <=  8'h20;        memory[61726] <=  8'h64;        memory[61727] <=  8'h66;        memory[61728] <=  8'h6a;        memory[61729] <=  8'h6b;        memory[61730] <=  8'h71;        memory[61731] <=  8'h64;        memory[61732] <=  8'h77;        memory[61733] <=  8'h65;        memory[61734] <=  8'h6e;        memory[61735] <=  8'h62;        memory[61736] <=  8'h20;        memory[61737] <=  8'h64;        memory[61738] <=  8'h73;        memory[61739] <=  8'h76;        memory[61740] <=  8'h68;        memory[61741] <=  8'h64;        memory[61742] <=  8'h61;        memory[61743] <=  8'h71;        memory[61744] <=  8'h77;        memory[61745] <=  8'h6a;        memory[61746] <=  8'h65;        memory[61747] <=  8'h6e;        memory[61748] <=  8'h64;        memory[61749] <=  8'h20;        memory[61750] <=  8'h61;        memory[61751] <=  8'h63;        memory[61752] <=  8'h62;        memory[61753] <=  8'h68;        memory[61754] <=  8'h64;        memory[61755] <=  8'h61;        memory[61756] <=  8'h77;        memory[61757] <=  8'h71;        memory[61758] <=  8'h6e;        memory[61759] <=  8'h20;        memory[61760] <=  8'h62;        memory[61761] <=  8'h73;        memory[61762] <=  8'h76;        memory[61763] <=  8'h61;        memory[61764] <=  8'h67;        memory[61765] <=  8'h76;        memory[61766] <=  8'h68;        memory[61767] <=  8'h67;        memory[61768] <=  8'h61;        memory[61769] <=  8'h73;        memory[61770] <=  8'h6a;        memory[61771] <=  8'h6b;        memory[61772] <=  8'h63;        memory[61773] <=  8'h78;        memory[61774] <=  8'h76;        memory[61775] <=  8'h6e;        memory[61776] <=  8'h73;        memory[61777] <=  8'h64;        memory[61778] <=  8'h20;        memory[61779] <=  8'h66;        memory[61780] <=  8'h62;        memory[61781] <=  8'h64;        memory[61782] <=  8'h61;        memory[61783] <=  8'h73;        memory[61784] <=  8'h76;        memory[61785] <=  8'h67;        memory[61786] <=  8'h63;        memory[61787] <=  8'h79;        memory[61788] <=  8'h7a;        memory[61789] <=  8'h78;        memory[61790] <=  8'h79;        memory[61791] <=  8'h75;        memory[61792] <=  8'h20;        memory[61793] <=  8'h69;        memory[61794] <=  8'h6a;        memory[61795] <=  8'h64;        memory[61796] <=  8'h66;        memory[61797] <=  8'h6b;        memory[61798] <=  8'h61;        memory[61799] <=  8'h64;        memory[61800] <=  8'h63;        memory[61801] <=  8'h78;        memory[61802] <=  8'h68;        memory[61803] <=  8'h20;        memory[61804] <=  8'h67;        memory[61805] <=  8'h61;        memory[61806] <=  8'h68;        memory[61807] <=  8'h75;        memory[61808] <=  8'h64;        memory[61809] <=  8'h73;        memory[61810] <=  8'h69;        memory[61811] <=  8'h6a;        memory[61812] <=  8'h61;        memory[61813] <=  8'h6b;        memory[61814] <=  8'h63;        memory[61815] <=  8'h62;        memory[61816] <=  8'h61;        memory[61817] <=  8'h72;        memory[61818] <=  8'h73;        memory[61819] <=  8'h68;        memory[61820] <=  8'h64;        memory[61821] <=  8'h66;        memory[61822] <=  8'h67;        memory[61823] <=  8'h73;        memory[61824] <=  8'h68;        memory[61825] <=  8'h64;        memory[61826] <=  8'h66;        memory[61827] <=  8'h68;        memory[61828] <=  8'h64;        memory[61829] <=  8'h6a;        memory[61830] <=  8'h68;        memory[61831] <=  8'h62;        memory[61832] <=  8'h67;        memory[61833] <=  8'h63;        memory[61834] <=  8'h61;        memory[61835] <=  8'h66;        memory[61836] <=  8'h73;        memory[61837] <=  8'h79;        memory[61838] <=  8'h67;        memory[61839] <=  8'h6b;        memory[61840] <=  8'h75;        memory[61841] <=  8'h64;        memory[61842] <=  8'h68;        memory[61843] <=  8'h62;        memory[61844] <=  8'h77;        memory[61845] <=  8'h76;        memory[61846] <=  8'h67;        memory[61847] <=  8'h61;        memory[61848] <=  8'h66;        memory[61849] <=  8'h64;        memory[61850] <=  8'h74;        memory[61851] <=  8'h75;        memory[61852] <=  8'h66;        memory[61853] <=  8'h79;        memory[61854] <=  8'h67;        memory[61855] <=  8'h69;        memory[61856] <=  8'h75;        memory[61857] <=  8'h68;        memory[61858] <=  8'h6c;        memory[61859] <=  8'h6a;        memory[61860] <=  8'h62;        memory[61861] <=  8'h6b;        memory[61862] <=  8'h68;        memory[61863] <=  8'h76;        memory[61864] <=  8'h67;        memory[61865] <=  8'h63;        memory[61866] <=  8'h66;        memory[61867] <=  8'h78;        memory[61868] <=  8'h64;        memory[61869] <=  8'h74;        memory[61870] <=  8'h75;        memory[61871] <=  8'h79;        memory[61872] <=  8'h69;        memory[61873] <=  8'h75;        memory[61874] <=  8'h68;        memory[61875] <=  8'h6c;        memory[61876] <=  8'h6a;        memory[61877] <=  8'h6b;        memory[61878] <=  8'h67;        memory[61879] <=  8'h6a;        memory[61880] <=  8'h63;        memory[61881] <=  8'h66;        memory[61882] <=  8'h68;        memory[61883] <=  8'h64;        memory[61884] <=  8'h67;        memory[61885] <=  8'h72;        memory[61886] <=  8'h79;        memory[61887] <=  8'h74;        memory[61888] <=  8'h66;        memory[61889] <=  8'h75;        memory[61890] <=  8'h79;        memory[61891] <=  8'h69;        memory[61892] <=  8'h68;        memory[61893] <=  8'h6c;        memory[61894] <=  8'h62;        memory[61895] <=  8'h6d;        memory[61896] <=  8'h76;        memory[61897] <=  8'h6e;        memory[61898] <=  8'h63;        memory[61899] <=  8'h66;        memory[61900] <=  8'h68;        memory[61901] <=  8'h64;        memory[61902] <=  8'h74;        memory[61903] <=  8'h75;        memory[61904] <=  8'h67;        memory[61905] <=  8'h79;        memory[61906] <=  8'h69;        memory[61907] <=  8'h68;        memory[61908] <=  8'h75;        memory[61909] <=  8'h6a;        memory[61910] <=  8'h6c;        memory[61911] <=  8'h62;        memory[61912] <=  8'h6d;        memory[61913] <=  8'h76;        memory[61914] <=  8'h6e;        memory[61915] <=  8'h63;        memory[61916] <=  8'h66;        memory[61917] <=  8'h68;        memory[61918] <=  8'h67;        memory[61919] <=  8'h79;        memory[61920] <=  8'h68;        memory[61921] <=  8'h75;        memory[61922] <=  8'h6a;        memory[61923] <=  8'h6e;        memory[61924] <=  8'h2c;        memory[61925] <=  8'h62;        memory[61926] <=  8'h6e;        memory[61927] <=  8'h6d;        memory[61928] <=  8'h76;        memory[61929] <=  8'h6e;        memory[61930] <=  8'h63;        memory[61931] <=  8'h66;        memory[61932] <=  8'h68;        memory[61933] <=  8'h74;        memory[61934] <=  8'h79;        memory[61935] <=  8'h69;        memory[61936] <=  8'h75;        memory[61937] <=  8'h6c;        memory[61938] <=  8'h6a;        memory[61939] <=  8'h62;        memory[61940] <=  8'h6d;        memory[61941] <=  8'h76;        memory[61942] <=  8'h6e;        memory[61943] <=  8'h63;        memory[61944] <=  8'h66;        memory[61945] <=  8'h74;        memory[61946] <=  8'h75;        memory[61947] <=  8'h79;        memory[61948] <=  8'h69;        memory[61949] <=  8'h68;        memory[61950] <=  8'h6b;        memory[61951] <=  8'h62;        memory[61952] <=  8'h76;        memory[61953] <=  8'h63;        memory[61954] <=  8'h66;        memory[61955] <=  8'h67;        memory[61956] <=  8'h74;        memory[61957] <=  8'h75;        memory[61958] <=  8'h79;        memory[61959] <=  8'h69;        memory[61960] <=  8'h75;        memory[61961] <=  8'h68;        memory[61962] <=  8'h6a;        memory[61963] <=  8'h6b;        memory[61964] <=  8'h62;        memory[61965] <=  8'h76;        memory[61966] <=  8'h63;        memory[61967] <=  8'h66;        memory[61968] <=  8'h74;        memory[61969] <=  8'h75;        memory[61970] <=  8'h79;        memory[61971] <=  8'h69;        memory[61972] <=  8'h75;        memory[61973] <=  8'h6a;        memory[61974] <=  8'h6b;        memory[61975] <=  8'h6e;        memory[61976] <=  8'h62;        memory[61977] <=  8'h76;        memory[61978] <=  8'h67;        memory[61979] <=  8'h66;        memory[61980] <=  8'h74;        memory[61981] <=  8'h79;        memory[61982] <=  8'h75;        memory[61983] <=  8'h75;        memory[61984] <=  8'h69;        memory[61985] <=  8'h6a;        memory[61986] <=  8'h6b;        memory[61987] <=  8'h68;        memory[61988] <=  8'h62;        memory[61989] <=  8'h6a;        memory[61990] <=  8'h67;        memory[61991] <=  8'h68;        memory[61992] <=  8'h66;        memory[61993] <=  8'h79;        memory[61994] <=  8'h74;        memory[61995] <=  8'h79;        memory[61996] <=  8'h69;        memory[61997] <=  8'h75;        memory[61998] <=  8'h64;        memory[61999] <=  8'h6a;        memory[62000] <=  8'h6b;        memory[62001] <=  8'h68;        memory[62002] <=  8'h63;        memory[62003] <=  8'h7a;        memory[62004] <=  8'h67;        memory[62005] <=  8'h68;        memory[62006] <=  8'h74;        memory[62007] <=  8'h75;        memory[62008] <=  8'h79;        memory[62009] <=  8'h69;        memory[62010] <=  8'h61;        memory[62011] <=  8'h73;        memory[62012] <=  8'h75;        memory[62013] <=  8'h6a;        memory[62014] <=  8'h6b;        memory[62015] <=  8'h62;        memory[62016] <=  8'h6e;        memory[62017] <=  8'h61;        memory[62018] <=  8'h76;        memory[62019] <=  8'h63;        memory[62020] <=  8'h66;        memory[62021] <=  8'h68;        memory[62022] <=  8'h75;        memory[62023] <=  8'h61;        memory[62024] <=  8'h73;        memory[62025] <=  8'h79;        memory[62026] <=  8'h64;        memory[62027] <=  8'h75;        memory[62028] <=  8'h69;        memory[62029] <=  8'h6a;        memory[62030] <=  8'h61;        memory[62031] <=  8'h6b;        memory[62032] <=  8'h62;        memory[62033] <=  8'h63;        memory[62034] <=  8'h78;        memory[62035] <=  8'h68;        memory[62036] <=  8'h67;        memory[62037] <=  8'h79;        memory[62038] <=  8'h75;        memory[62039] <=  8'h7a;        memory[62040] <=  8'h63;        memory[62041] <=  8'h61;        memory[62042] <=  8'h73;        memory[62043] <=  8'h69;        memory[62044] <=  8'h75;        memory[62045] <=  8'h6f;        memory[62046] <=  8'h69;        memory[62047] <=  8'h6a;        memory[62048] <=  8'h61;        memory[62049] <=  8'h6c;        memory[62050] <=  8'h63;        memory[62051] <=  8'h78;        memory[62052] <=  8'h62;        memory[62053] <=  8'h63;        memory[62054] <=  8'h20;        memory[62055] <=  8'h6e;        memory[62056] <=  8'h76;        memory[62057] <=  8'h63;        memory[62058] <=  8'h61;        memory[62059] <=  8'h64;        memory[62060] <=  8'h73;        memory[62061] <=  8'h67;        memory[62062] <=  8'h79;        memory[62063] <=  8'h68;        memory[62064] <=  8'h75;        memory[62065] <=  8'h61;        memory[62066] <=  8'h6a;        memory[62067] <=  8'h6b;        memory[62068] <=  8'h78;        memory[62069] <=  8'h62;        memory[62070] <=  8'h20;        memory[62071] <=  8'h6e;        memory[62072] <=  8'h76;        memory[62073] <=  8'h63;        memory[62074] <=  8'h61;        memory[62075] <=  8'h73;        memory[62076] <=  8'h67;        memory[62077] <=  8'h68;        memory[62078] <=  8'h75;        memory[62079] <=  8'h6a;        memory[62080] <=  8'h6c;        memory[62081] <=  8'h6b;        memory[62082] <=  8'h63;        memory[62083] <=  8'h78;        memory[62084] <=  8'h20;        memory[62085] <=  8'h6a;        memory[62086] <=  8'h6b;        memory[62087] <=  8'h68;        memory[62088] <=  8'h61;        memory[62089] <=  8'h73;        memory[62090] <=  8'h76;        memory[62091] <=  8'h64;        memory[62092] <=  8'h6e;        memory[62093] <=  8'h20;        memory[62094] <=  8'h62;        memory[62095] <=  8'h6e;        memory[62096] <=  8'h6d;        memory[62097] <=  8'h6b;        memory[62098] <=  8'h77;        memory[62099] <=  8'h64;        memory[62100] <=  8'h6f;        memory[62101] <=  8'h77;        memory[62102] <=  8'h69;        memory[62103] <=  8'h6f;        memory[62104] <=  8'h75;        memory[62105] <=  8'h69;        memory[62106] <=  8'h68;        memory[62107] <=  8'h62;        memory[62108] <=  8'h6e;        memory[62109] <=  8'h6b;        memory[62110] <=  8'h77;        memory[62111] <=  8'h69;        memory[62112] <=  8'h6f;        memory[62113] <=  8'h75;        memory[62114] <=  8'h71;        memory[62115] <=  8'h69;        memory[62116] <=  8'h79;        memory[62117] <=  8'h67;        memory[62118] <=  8'h6a;        memory[62119] <=  8'h64;        memory[62120] <=  8'h61;        memory[62121] <=  8'h76;        memory[62122] <=  8'h62;        memory[62123] <=  8'h6e;        memory[62124] <=  8'h6b;        memory[62125] <=  8'h6f;        memory[62126] <=  8'h70;        memory[62127] <=  8'h64;        memory[62128] <=  8'h76;        memory[62129] <=  8'h69;        memory[62130] <=  8'h6f;        memory[62131] <=  8'h75;        memory[62132] <=  8'h69;        memory[62133] <=  8'h48;        memory[62134] <=  8'h42;        memory[62135] <=  8'h6b;        memory[62136] <=  8'h64;        memory[62137] <=  8'h6e;        memory[62138] <=  8'h6c;        memory[62139] <=  8'h71;        memory[62140] <=  8'h6b;        memory[62141] <=  8'h6d;        memory[62142] <=  8'h6a;        memory[62143] <=  8'h70;        memory[62144] <=  8'h69;        memory[62145] <=  8'h6f;        memory[62146] <=  8'h68;        memory[62147] <=  8'h65;        memory[62148] <=  8'h66;        memory[62149] <=  8'h75;        memory[62150] <=  8'h67;        memory[62151] <=  8'h69;        memory[62152] <=  8'h73;        memory[62153] <=  8'h61;        memory[62154] <=  8'h62;        memory[62155] <=  8'h64;        memory[62156] <=  8'h6b;        memory[62157] <=  8'h6a;        memory[62158] <=  8'h6b;        memory[62159] <=  8'h6c;        memory[62160] <=  8'h6a;        memory[62161] <=  8'h69;        memory[62162] <=  8'h73;        memory[62163] <=  8'h6f;        memory[62164] <=  8'h71;        memory[62165] <=  8'h68;        memory[62166] <=  8'h77;        memory[62167] <=  8'h67;        memory[62168] <=  8'h69;        memory[62169] <=  8'h79;        memory[62170] <=  8'h6a;        memory[62171] <=  8'h64;        memory[62172] <=  8'h76;        memory[62173] <=  8'h62;        memory[62174] <=  8'h6e;        memory[62175] <=  8'h61;        memory[62176] <=  8'h73;        memory[62177] <=  8'h66;        memory[62178] <=  8'h6c;        memory[62179] <=  8'h6b;        memory[62180] <=  8'h64;        memory[62181] <=  8'h6a;        memory[62182] <=  8'h68;        memory[62183] <=  8'h63;        memory[62184] <=  8'h67;        memory[62185] <=  8'h6a;        memory[62186] <=  8'h76;        memory[62187] <=  8'h73;        memory[62188] <=  8'h64;        memory[62189] <=  8'h62;        memory[62190] <=  8'h62;        memory[62191] <=  8'h61;        memory[62192] <=  8'h72;        memory[62193] <=  8'h62;        memory[62194] <=  8'h62;        memory[62195] <=  8'h73;        memory[62196] <=  8'h62;        memory[62197] <=  8'h67;        memory[62198] <=  8'h73;        memory[62199] <=  8'h66;        memory[62200] <=  8'h67;        memory[62201] <=  8'h61;        memory[62202] <=  8'h68;        memory[62203] <=  8'h66;        memory[62204] <=  8'h73;        memory[62205] <=  8'h68;        memory[62206] <=  8'h61;        memory[62207] <=  8'h66;        memory[62208] <=  8'h73;        memory[62209] <=  8'h66;        memory[62210] <=  8'h68;        memory[62211] <=  8'h61;        memory[62212] <=  8'h69;        memory[62213] <=  8'h64;        memory[62214] <=  8'h75;        memory[62215] <=  8'h67;        memory[62216] <=  8'h64;        memory[62217] <=  8'h77;        memory[62218] <=  8'h62;        memory[62219] <=  8'h61;        memory[62220] <=  8'h62;        memory[62221] <=  8'h72;        memory[62222] <=  8'h62;        memory[62223] <=  8'h61;        memory[62224] <=  8'h62;        memory[62225] <=  8'h62;        memory[62226] <=  8'h74;        memory[62227] <=  8'h62;        memory[62228] <=  8'h62;        memory[62229] <=  8'h62;        memory[62230] <=  8'h62;        memory[62231] <=  8'h62;        memory[62232] <=  8'h62;        memory[62233] <=  8'h62;        memory[62234] <=  8'h62;        memory[62235] <=  8'h61;        memory[62236] <=  8'h62;        memory[62237] <=  8'h62;        memory[62238] <=  8'h72;        memory[62239] <=  8'h74;        memory[62240] <=  8'h62;        memory[62241] <=  8'h62;        memory[62242] <=  8'h61;        memory[62243] <=  8'h62;        memory[62244] <=  8'h72;        memory[62245] <=  8'h62;        memory[62246] <=  8'h74;        memory[62247] <=  8'h62;        memory[62248] <=  8'h62;        memory[62249] <=  8'h62;        memory[62250] <=  8'h63;        memory[62251] <=  8'h61;        memory[62252] <=  8'h72;        memory[62253] <=  8'h74;        memory[62254] <=  8'h73;        memory[62255] <=  8'h62;        memory[62256] <=  8'h61;        memory[62257] <=  8'h72;        memory[62258] <=  8'h74;        memory[62259] <=  8'h74;        memory[62260] <=  8'h62;        memory[62261] <=  8'h61;        memory[62262] <=  8'h72;        memory[62263] <=  8'h74;        memory[62264] <=  8'h78;        memory[62265] <=  8'h61;        memory[62266] <=  8'h74;        memory[62267] <=  8'h6b;        memory[62268] <=  8'h73;        memory[62269] <=  8'h68;        memory[62270] <=  8'h63;        memory[62271] <=  8'h66;        memory[62272] <=  8'h69;        memory[62273] <=  8'h77;        memory[62274] <=  8'h68;        memory[62275] <=  8'h61;        memory[62276] <=  8'h74;        memory[62277] <=  8'h61;        memory[62278] <=  8'h6e;        memory[62279] <=  8'h61;        memory[62280] <=  8'h62;        memory[62281] <=  8'h61;        memory[62282] <=  8'h63;        memory[62283] <=  8'h61;        memory[62284] <=  8'h74;        memory[62285] <=  8'h61;        memory[62286] <=  8'h62;        memory[62287] <=  8'h61;        memory[62288] <=  8'h72;        memory[62289] <=  8'h63;        memory[62290] <=  8'h61;        memory[62291] <=  8'h68;        memory[62292] <=  8'h64;        memory[62293] <=  8'h75;        memory[62294] <=  8'h63;        memory[62295] <=  8'h74;        memory[62296] <=  8'h61;        memory[62297] <=  8'h64;        memory[62298] <=  8'h61;        memory[62299] <=  8'h61;        memory[62300] <=  8'h63;        memory[62301] <=  8'h61;        memory[62302] <=  8'h72;        memory[62303] <=  8'h63;        memory[62304] <=  8'h74;        memory[62305] <=  8'h72;        memory[62306] <=  8'h63;        memory[62307] <=  8'h61;        memory[62308] <=  8'h74;        memory[62309] <=  8'h72;        memory[62310] <=  8'h63;        memory[62311] <=  8'h61;        memory[62312] <=  8'h74;        memory[62313] <=  8'h63;        memory[62314] <=  8'h62;        memory[62315] <=  8'h61;        memory[62316] <=  8'h74;        memory[62317] <=  8'h62;        memory[62318] <=  8'h72;        memory[62319] <=  8'h63;        memory[62320] <=  8'h61;        memory[62321] <=  8'h74;        memory[62322] <=  8'h72;        memory[62323] <=  8'h6e;        memory[62324] <=  8'h62;        memory[62325] <=  8'h61;        memory[62326] <=  8'h63;        memory[62327] <=  8'h61;        memory[62328] <=  8'h74;        memory[62329] <=  8'h79;        memory[62330] <=  8'h73;        memory[62331] <=  8'h6e;        memory[62332] <=  8'h63;        memory[62333] <=  8'h74;        memory[62334] <=  8'h61;        memory[62335] <=  8'h6e;        memory[62336] <=  8'h62;        memory[62337] <=  8'h61;        memory[62338] <=  8'h63;        memory[62339] <=  8'h72;        memory[62340] <=  8'h6e;        memory[62341] <=  8'h74;        memory[62342] <=  8'h61;        memory[62343] <=  8'h62;        memory[62344] <=  8'h74;        memory[62345] <=  8'h6e;        memory[62346] <=  8'h61;        memory[62347] <=  8'h72;        memory[62348] <=  8'h62;        memory[62349] <=  8'h78;        memory[62350] <=  8'h74;        memory[62351] <=  8'h61;        memory[62352] <=  8'h72;        memory[62353] <=  8'h62;        memory[62354] <=  8'h61;        memory[62355] <=  8'h72;        memory[62356] <=  8'h74;        memory[62357] <=  8'h74;        memory[62358] <=  8'h62;        memory[62359] <=  8'h61;        memory[62360] <=  8'h72;        memory[62361] <=  8'h74;        memory[62362] <=  8'h78;        memory[62363] <=  8'h61;        memory[62364] <=  8'h74;        memory[62365] <=  8'h6b;        memory[62366] <=  8'h73;        memory[62367] <=  8'h68;        memory[62368] <=  8'h63;        memory[62369] <=  8'h66;        memory[62370] <=  8'h69;        memory[62371] <=  8'h77;        memory[62372] <=  8'h68;        memory[62373] <=  8'h61;        memory[62374] <=  8'h74;        memory[62375] <=  8'h61;        memory[62376] <=  8'h6e;        memory[62377] <=  8'h61;        memory[62378] <=  8'h62;        memory[62379] <=  8'h61;        memory[62380] <=  8'h63;        memory[62381] <=  8'h61;        memory[62382] <=  8'h74;        memory[62383] <=  8'h61;        memory[62384] <=  8'h62;        memory[62385] <=  8'h61;        memory[62386] <=  8'h72;        memory[62387] <=  8'h63;        memory[62388] <=  8'h61;        memory[62389] <=  8'h68;        memory[62390] <=  8'h64;        memory[62391] <=  8'h75;        memory[62392] <=  8'h63;        memory[62393] <=  8'h74;        memory[62394] <=  8'h61;        memory[62395] <=  8'h64;        memory[62396] <=  8'h61;        memory[62397] <=  8'h61;        memory[62398] <=  8'h63;        memory[62399] <=  8'h61;        memory[62400] <=  8'h72;        memory[62401] <=  8'h63;        memory[62402] <=  8'h74;        memory[62403] <=  8'h72;        memory[62404] <=  8'h63;        memory[62405] <=  8'h61;        memory[62406] <=  8'h74;        memory[62407] <=  8'h72;        memory[62408] <=  8'h63;        memory[62409] <=  8'h61;        memory[62410] <=  8'h74;        memory[62411] <=  8'h63;        memory[62412] <=  8'h62;        memory[62413] <=  8'h61;        memory[62414] <=  8'h74;        memory[62415] <=  8'h62;        memory[62416] <=  8'h72;        memory[62417] <=  8'h63;        memory[62418] <=  8'h61;        memory[62419] <=  8'h74;        memory[62420] <=  8'h72;        memory[62421] <=  8'h6e;        memory[62422] <=  8'h62;        memory[62423] <=  8'h61;        memory[62424] <=  8'h63;        memory[62425] <=  8'h61;        memory[62426] <=  8'h74;        memory[62427] <=  8'h79;        memory[62428] <=  8'h73;        memory[62429] <=  8'h6e;        memory[62430] <=  8'h63;        memory[62431] <=  8'h74;        memory[62432] <=  8'h61;        memory[62433] <=  8'h6e;        memory[62434] <=  8'h62;        memory[62435] <=  8'h61;        memory[62436] <=  8'h63;        memory[62437] <=  8'h72;        memory[62438] <=  8'h6e;        memory[62439] <=  8'h74;        memory[62440] <=  8'h61;        memory[62441] <=  8'h62;        memory[62442] <=  8'h74;        memory[62443] <=  8'h6e;        memory[62444] <=  8'h61;        memory[62445] <=  8'h72;        memory[62446] <=  8'h62;        memory[62447] <=  8'h78;        memory[62448] <=  8'h74;        memory[62449] <=  8'h61;        memory[62450] <=  8'h72;        memory[62451] <=  8'h62;        memory[62452] <=  8'h61;        memory[62453] <=  8'h72;        memory[62454] <=  8'h74;        memory[62455] <=  8'h74;        memory[62456] <=  8'h62;        memory[62457] <=  8'h61;        memory[62458] <=  8'h72;        memory[62459] <=  8'h74;        memory[62460] <=  8'h78;        memory[62461] <=  8'h61;        memory[62462] <=  8'h74;        memory[62463] <=  8'h6b;        memory[62464] <=  8'h73;        memory[62465] <=  8'h68;        memory[62466] <=  8'h63;        memory[62467] <=  8'h66;        memory[62468] <=  8'h69;        memory[62469] <=  8'h77;        memory[62470] <=  8'h68;        memory[62471] <=  8'h61;        memory[62472] <=  8'h74;        memory[62473] <=  8'h61;        memory[62474] <=  8'h6e;        memory[62475] <=  8'h61;        memory[62476] <=  8'h62;        memory[62477] <=  8'h61;        memory[62478] <=  8'h63;        memory[62479] <=  8'h61;        memory[62480] <=  8'h74;        memory[62481] <=  8'h61;        memory[62482] <=  8'h62;        memory[62483] <=  8'h61;        memory[62484] <=  8'h72;        memory[62485] <=  8'h63;        memory[62486] <=  8'h61;        memory[62487] <=  8'h68;        memory[62488] <=  8'h64;        memory[62489] <=  8'h75;        memory[62490] <=  8'h63;        memory[62491] <=  8'h74;        memory[62492] <=  8'h61;        memory[62493] <=  8'h64;        memory[62494] <=  8'h61;        memory[62495] <=  8'h61;        memory[62496] <=  8'h63;        memory[62497] <=  8'h61;        memory[62498] <=  8'h72;        memory[62499] <=  8'h63;        memory[62500] <=  8'h74;        memory[62501] <=  8'h72;        memory[62502] <=  8'h63;        memory[62503] <=  8'h61;        memory[62504] <=  8'h74;        memory[62505] <=  8'h72;        memory[62506] <=  8'h63;        memory[62507] <=  8'h61;        memory[62508] <=  8'h74;        memory[62509] <=  8'h63;        memory[62510] <=  8'h62;        memory[62511] <=  8'h61;        memory[62512] <=  8'h74;        memory[62513] <=  8'h62;        memory[62514] <=  8'h72;        memory[62515] <=  8'h63;        memory[62516] <=  8'h61;        memory[62517] <=  8'h74;        memory[62518] <=  8'h72;        memory[62519] <=  8'h6e;        memory[62520] <=  8'h62;        memory[62521] <=  8'h61;        memory[62522] <=  8'h63;        memory[62523] <=  8'h61;        memory[62524] <=  8'h74;        memory[62525] <=  8'h79;        memory[62526] <=  8'h73;        memory[62527] <=  8'h6e;        memory[62528] <=  8'h63;        memory[62529] <=  8'h74;        memory[62530] <=  8'h61;        memory[62531] <=  8'h6e;        memory[62532] <=  8'h62;        memory[62533] <=  8'h61;        memory[62534] <=  8'h63;        memory[62535] <=  8'h72;        memory[62536] <=  8'h6e;        memory[62537] <=  8'h74;        memory[62538] <=  8'h61;        memory[62539] <=  8'h62;        memory[62540] <=  8'h74;        memory[62541] <=  8'h6e;        memory[62542] <=  8'h61;        memory[62543] <=  8'h72;        memory[62544] <=  8'h62;        memory[62545] <=  8'h78;        memory[62546] <=  8'h74;        memory[62547] <=  8'h61;        memory[62548] <=  8'h72;        memory[62549] <=  8'h5d;        memory[62550] <=  8'h5d;        memory[62551] <=  8'h65;        memory[62552] <=  8'h66;        memory[62553] <=  8'h77;        memory[62554] <=  8'h65;        memory[62555] <=  8'h5d;        memory[62556] <=  8'h65;        memory[62557] <=  8'h67;        memory[62558] <=  8'h73;        memory[62559] <=  8'h67;        memory[62560] <=  8'h66;        memory[62561] <=  8'h62;        memory[62562] <=  8'h61;        memory[62563] <=  8'h72;        memory[62564] <=  8'h74;        memory[62565] <=  8'h74;        memory[62566] <=  8'h62;        memory[62567] <=  8'h61;        memory[62568] <=  8'h72;        memory[62569] <=  8'h74;        memory[62570] <=  8'h78;        memory[62571] <=  8'h61;        memory[62572] <=  8'h74;        memory[62573] <=  8'h6b;        memory[62574] <=  8'h73;        memory[62575] <=  8'h68;        memory[62576] <=  8'h63;        memory[62577] <=  8'h66;        memory[62578] <=  8'h69;        memory[62579] <=  8'h77;        memory[62580] <=  8'h68;        memory[62581] <=  8'h61;        memory[62582] <=  8'h74;        memory[62583] <=  8'h61;        memory[62584] <=  8'h6e;        memory[62585] <=  8'h61;        memory[62586] <=  8'h62;        memory[62587] <=  8'h61;        memory[62588] <=  8'h63;        memory[62589] <=  8'h61;        memory[62590] <=  8'h74;        memory[62591] <=  8'h61;        memory[62592] <=  8'h62;        memory[62593] <=  8'h61;        memory[62594] <=  8'h72;        memory[62595] <=  8'h63;        memory[62596] <=  8'h61;        memory[62597] <=  8'h68;        memory[62598] <=  8'h64;        memory[62599] <=  8'h75;        memory[62600] <=  8'h63;        memory[62601] <=  8'h74;        memory[62602] <=  8'h61;        memory[62603] <=  8'h64;        memory[62604] <=  8'h61;        memory[62605] <=  8'h61;        memory[62606] <=  8'h63;        memory[62607] <=  8'h61;        memory[62608] <=  8'h72;        memory[62609] <=  8'h63;        memory[62610] <=  8'h74;        memory[62611] <=  8'h72;        memory[62612] <=  8'h63;        memory[62613] <=  8'h61;        memory[62614] <=  8'h74;        memory[62615] <=  8'h72;        memory[62616] <=  8'h63;        memory[62617] <=  8'h61;        memory[62618] <=  8'h74;        memory[62619] <=  8'h63;        memory[62620] <=  8'h62;        memory[62621] <=  8'h61;        memory[62622] <=  8'h74;        memory[62623] <=  8'h62;        memory[62624] <=  8'h72;        memory[62625] <=  8'h63;        memory[62626] <=  8'h61;        memory[62627] <=  8'h74;        memory[62628] <=  8'h72;        memory[62629] <=  8'h6e;        memory[62630] <=  8'h62;        memory[62631] <=  8'h61;        memory[62632] <=  8'h63;        memory[62633] <=  8'h61;        memory[62634] <=  8'h74;        memory[62635] <=  8'h79;        memory[62636] <=  8'h73;        memory[62637] <=  8'h6e;        memory[62638] <=  8'h63;        memory[62639] <=  8'h74;        memory[62640] <=  8'h61;        memory[62641] <=  8'h6e;        memory[62642] <=  8'h62;        memory[62643] <=  8'h61;        memory[62644] <=  8'h63;        memory[62645] <=  8'h72;        memory[62646] <=  8'h6e;        memory[62647] <=  8'h74;        memory[62648] <=  8'h61;        memory[62649] <=  8'h62;        memory[62650] <=  8'h74;        memory[62651] <=  8'h6e;        memory[62652] <=  8'h61;        memory[62653] <=  8'h72;        memory[62654] <=  8'h62;        memory[62655] <=  8'h78;        memory[62656] <=  8'h74;        memory[62657] <=  8'h61;        memory[62658] <=  8'h72;        memory[62659] <=  8'h62;        memory[62660] <=  8'h61;        memory[62661] <=  8'h72;        memory[62662] <=  8'h74;        memory[62663] <=  8'h74;        memory[62664] <=  8'h62;        memory[62665] <=  8'h61;        memory[62666] <=  8'h72;        memory[62667] <=  8'h74;        memory[62668] <=  8'h78;        memory[62669] <=  8'h61;        memory[62670] <=  8'h74;        memory[62671] <=  8'h6b;        memory[62672] <=  8'h73;        memory[62673] <=  8'h68;        memory[62674] <=  8'h63;        memory[62675] <=  8'h66;        memory[62676] <=  8'h69;        memory[62677] <=  8'h77;        memory[62678] <=  8'h68;        memory[62679] <=  8'h61;        memory[62680] <=  8'h74;        memory[62681] <=  8'h61;        memory[62682] <=  8'h6e;        memory[62683] <=  8'h61;        memory[62684] <=  8'h62;        memory[62685] <=  8'h61;        memory[62686] <=  8'h63;        memory[62687] <=  8'h61;        memory[62688] <=  8'h74;        memory[62689] <=  8'h61;        memory[62690] <=  8'h62;        memory[62691] <=  8'h61;        memory[62692] <=  8'h72;        memory[62693] <=  8'h63;        memory[62694] <=  8'h61;        memory[62695] <=  8'h68;        memory[62696] <=  8'h64;        memory[62697] <=  8'h75;        memory[62698] <=  8'h63;        memory[62699] <=  8'h74;        memory[62700] <=  8'h61;        memory[62701] <=  8'h64;        memory[62702] <=  8'h61;        memory[62703] <=  8'h61;        memory[62704] <=  8'h63;        memory[62705] <=  8'h61;        memory[62706] <=  8'h72;        memory[62707] <=  8'h63;        memory[62708] <=  8'h74;        memory[62709] <=  8'h72;        memory[62710] <=  8'h63;        memory[62711] <=  8'h61;        memory[62712] <=  8'h74;        memory[62713] <=  8'h72;        memory[62714] <=  8'h63;        memory[62715] <=  8'h61;        memory[62716] <=  8'h74;        memory[62717] <=  8'h63;        memory[62718] <=  8'h62;        memory[62719] <=  8'h61;        memory[62720] <=  8'h74;        memory[62721] <=  8'h62;        memory[62722] <=  8'h72;        memory[62723] <=  8'h63;        memory[62724] <=  8'h61;        memory[62725] <=  8'h74;        memory[62726] <=  8'h72;        memory[62727] <=  8'h6e;        memory[62728] <=  8'h62;        memory[62729] <=  8'h61;        memory[62730] <=  8'h63;        memory[62731] <=  8'h61;        memory[62732] <=  8'h74;        memory[62733] <=  8'h79;        memory[62734] <=  8'h73;        memory[62735] <=  8'h6e;        memory[62736] <=  8'h63;        memory[62737] <=  8'h74;        memory[62738] <=  8'h61;        memory[62739] <=  8'h6e;        memory[62740] <=  8'h62;        memory[62741] <=  8'h61;        memory[62742] <=  8'h63;        memory[62743] <=  8'h72;        memory[62744] <=  8'h6e;        memory[62745] <=  8'h74;        memory[62746] <=  8'h61;        memory[62747] <=  8'h62;        memory[62748] <=  8'h74;        memory[62749] <=  8'h6e;        memory[62750] <=  8'h61;        memory[62751] <=  8'h72;        memory[62752] <=  8'h62;        memory[62753] <=  8'h78;        memory[62754] <=  8'h74;        memory[62755] <=  8'h61;        memory[62756] <=  8'h72;        memory[62757] <=  8'h64;        memory[62758] <=  8'h66;        memory[62759] <=  8'h73;        memory[62760] <=  8'h67;        memory[62761] <=  8'h76;        memory[62762] <=  8'h68;        memory[62763] <=  8'h62;        memory[62764] <=  8'h6b;        memory[62765] <=  8'h6a;        memory[62766] <=  8'h6e;        memory[62767] <=  8'h6d;        memory[62768] <=  8'h62;        memory[62769] <=  8'h76;        memory[62770] <=  8'h78;        memory[62771] <=  8'h63;        memory[62772] <=  8'h73;        memory[62773] <=  8'h66;        memory[62774] <=  8'h72;        memory[62775] <=  8'h74;        memory[62776] <=  8'h79;        memory[62777] <=  8'h75;        memory[62778] <=  8'h6a;        memory[62779] <=  8'h6e;        memory[62780] <=  8'h62;        memory[62781] <=  8'h76;        memory[62782] <=  8'h63;        memory[62783] <=  8'h64;        memory[62784] <=  8'h74;        memory[62785] <=  8'h79;        memory[62786] <=  8'h75;        memory[62787] <=  8'h69;        memory[62788] <=  8'h6b;        memory[62789] <=  8'h6d;        memory[62790] <=  8'h6e;        memory[62791] <=  8'h62;        memory[62792] <=  8'h76;        memory[62793] <=  8'h63;        memory[62794] <=  8'h78;        memory[62795] <=  8'h73;        memory[62796] <=  8'h64;        memory[62797] <=  8'h72;        memory[62798] <=  8'h74;        memory[62799] <=  8'h79;        memory[62800] <=  8'h75;        memory[62801] <=  8'h69;        memory[62802] <=  8'h6b;        memory[62803] <=  8'h6d;        memory[62804] <=  8'h6e;        memory[62805] <=  8'h62;        memory[62806] <=  8'h76;        memory[62807] <=  8'h63;        memory[62808] <=  8'h73;        memory[62809] <=  8'h77;        memory[62810] <=  8'h33;        memory[62811] <=  8'h34;        memory[62812] <=  8'h35;        memory[62813] <=  8'h36;        memory[62814] <=  8'h37;        memory[62815] <=  8'h38;        memory[62816] <=  8'h69;        memory[62817] <=  8'h6b;        memory[62818] <=  8'h6d;        memory[62819] <=  8'h6e;        memory[62820] <=  8'h62;        memory[62821] <=  8'h76;        memory[62822] <=  8'h63;        memory[62823] <=  8'h64;        memory[62824] <=  8'h65;        memory[62825] <=  8'h72;        memory[62826] <=  8'h36;        memory[62827] <=  8'h37;        memory[62828] <=  8'h38;        memory[62829] <=  8'h69;        memory[62830] <=  8'h6f;        memory[62831] <=  8'h6b;        memory[62832] <=  8'h6a;        memory[62833] <=  8'h6e;        memory[62834] <=  8'h62;        memory[62835] <=  8'h76;        memory[62836] <=  8'h63;        memory[62837] <=  8'h64;        memory[62838] <=  8'h72;        memory[62839] <=  8'h74;        memory[62840] <=  8'h79;        memory[62841] <=  8'h75;        memory[62842] <=  8'h73;        memory[62843] <=  8'h6a;        memory[62844] <=  8'h63;        memory[62845] <=  8'h6e;        memory[62846] <=  8'h62;        memory[62847] <=  8'h64;        memory[62848] <=  8'h66;        memory[62849] <=  8'h73;        memory[62850] <=  8'h74;        memory[62851] <=  8'h79;        memory[62852] <=  8'h75;        memory[62853] <=  8'h61;        memory[62854] <=  8'h69;        memory[62855] <=  8'h6b;        memory[62856] <=  8'h78;        memory[62857] <=  8'h6d;        memory[62858] <=  8'h6e;        memory[62859] <=  8'h73;        memory[62860] <=  8'h6a;        memory[62861] <=  8'h6f;        memory[62862] <=  8'h64;        memory[62863] <=  8'h6c;        memory[62864] <=  8'h63;        memory[62865] <=  8'h78;        memory[62866] <=  8'h62;        memory[62867] <=  8'h61;        memory[62868] <=  8'h72;        memory[62869] <=  8'h74;        memory[62870] <=  8'h78;        memory[62871] <=  8'h61;        memory[62872] <=  8'h74;        memory[62873] <=  8'h6b;        memory[62874] <=  8'h73;        memory[62875] <=  8'h68;        memory[62876] <=  8'h63;        memory[62877] <=  8'h66;        memory[62878] <=  8'h69;        memory[62879] <=  8'h77;        memory[62880] <=  8'h68;        memory[62881] <=  8'h61;        memory[62882] <=  8'h74;        memory[62883] <=  8'h61;        memory[62884] <=  8'h6e;        memory[62885] <=  8'h61;        memory[62886] <=  8'h62;        memory[62887] <=  8'h61;        memory[62888] <=  8'h63;        memory[62889] <=  8'h61;        memory[62890] <=  8'h74;        memory[62891] <=  8'h61;        memory[62892] <=  8'h62;        memory[62893] <=  8'h61;        memory[62894] <=  8'h72;        memory[62895] <=  8'h63;        memory[62896] <=  8'h61;        memory[62897] <=  8'h68;        memory[62898] <=  8'h64;        memory[62899] <=  8'h75;        memory[62900] <=  8'h63;        memory[62901] <=  8'h74;        memory[62902] <=  8'h61;        memory[62903] <=  8'h64;        memory[62904] <=  8'h61;        memory[62905] <=  8'h61;        memory[62906] <=  8'h63;        memory[62907] <=  8'h61;        memory[62908] <=  8'h72;        memory[62909] <=  8'h62;        memory[62910] <=  8'h61;        memory[62911] <=  8'h72;        memory[62912] <=  8'h74;        memory[62913] <=  8'h78;        memory[62914] <=  8'h61;        memory[62915] <=  8'h74;        memory[62916] <=  8'h6b;        memory[62917] <=  8'h73;        memory[62918] <=  8'h68;        memory[62919] <=  8'h63;        memory[62920] <=  8'h66;        memory[62921] <=  8'h69;        memory[62922] <=  8'h77;        memory[62923] <=  8'h68;        memory[62924] <=  8'h61;        memory[62925] <=  8'h74;        memory[62926] <=  8'h61;        memory[62927] <=  8'h6e;        memory[62928] <=  8'h61;        memory[62929] <=  8'h62;        memory[62930] <=  8'h61;        memory[62931] <=  8'h63;        memory[62932] <=  8'h61;        memory[62933] <=  8'h74;        memory[62934] <=  8'h61;        memory[62935] <=  8'h62;        memory[62936] <=  8'h61;        memory[62937] <=  8'h72;        memory[62938] <=  8'h63;        memory[62939] <=  8'h61;        memory[62940] <=  8'h68;        memory[62941] <=  8'h64;        memory[62942] <=  8'h75;        memory[62943] <=  8'h63;        memory[62944] <=  8'h74;        memory[62945] <=  8'h61;        memory[62946] <=  8'h64;        memory[62947] <=  8'h61;        memory[62948] <=  8'h61;        memory[62949] <=  8'h63;        memory[62950] <=  8'h61;        memory[62951] <=  8'h72;        memory[62952] <=  8'h62;        memory[62953] <=  8'h61;        memory[62954] <=  8'h72;        memory[62955] <=  8'h74;        memory[62956] <=  8'h78;        memory[62957] <=  8'h61;        memory[62958] <=  8'h74;        memory[62959] <=  8'h6b;        memory[62960] <=  8'h73;        memory[62961] <=  8'h68;        memory[62962] <=  8'h63;        memory[62963] <=  8'h66;        memory[62964] <=  8'h69;        memory[62965] <=  8'h77;        memory[62966] <=  8'h68;        memory[62967] <=  8'h61;        memory[62968] <=  8'h74;        memory[62969] <=  8'h61;        memory[62970] <=  8'h6e;        memory[62971] <=  8'h61;        memory[62972] <=  8'h62;        memory[62973] <=  8'h61;        memory[62974] <=  8'h63;        memory[62975] <=  8'h61;        memory[62976] <=  8'h74;        memory[62977] <=  8'h61;        memory[62978] <=  8'h62;        memory[62979] <=  8'h61;        memory[62980] <=  8'h72;        memory[62981] <=  8'h63;        memory[62982] <=  8'h61;        memory[62983] <=  8'h68;        memory[62984] <=  8'h64;        memory[62985] <=  8'h75;        memory[62986] <=  8'h63;        memory[62987] <=  8'h74;        memory[62988] <=  8'h61;        memory[62989] <=  8'h64;        memory[62990] <=  8'h61;        memory[62991] <=  8'h61;        memory[62992] <=  8'h63;        memory[62993] <=  8'h61;        memory[62994] <=  8'h72;        memory[62995] <=  8'h62;        memory[62996] <=  8'h61;        memory[62997] <=  8'h72;        memory[62998] <=  8'h74;        memory[62999] <=  8'h78;        memory[63000] <=  8'h61;        memory[63001] <=  8'h74;        memory[63002] <=  8'h6b;        memory[63003] <=  8'h73;        memory[63004] <=  8'h68;        memory[63005] <=  8'h63;        memory[63006] <=  8'h66;        memory[63007] <=  8'h69;        memory[63008] <=  8'h77;        memory[63009] <=  8'h68;        memory[63010] <=  8'h61;        memory[63011] <=  8'h74;        memory[63012] <=  8'h61;        memory[63013] <=  8'h6e;        memory[63014] <=  8'h61;        memory[63015] <=  8'h62;        memory[63016] <=  8'h61;        memory[63017] <=  8'h63;        memory[63018] <=  8'h61;        memory[63019] <=  8'h74;        memory[63020] <=  8'h61;        memory[63021] <=  8'h62;        memory[63022] <=  8'h61;        memory[63023] <=  8'h72;        memory[63024] <=  8'h63;        memory[63025] <=  8'h61;        memory[63026] <=  8'h68;        memory[63027] <=  8'h64;        memory[63028] <=  8'h75;        memory[63029] <=  8'h63;        memory[63030] <=  8'h74;        memory[63031] <=  8'h61;        memory[63032] <=  8'h64;        memory[63033] <=  8'h61;        memory[63034] <=  8'h61;        memory[63035] <=  8'h63;        memory[63036] <=  8'h61;        memory[63037] <=  8'h72;        memory[63038] <=  8'h62;        memory[63039] <=  8'h61;        memory[63040] <=  8'h72;        memory[63041] <=  8'h74;        memory[63042] <=  8'h78;        memory[63043] <=  8'h61;        memory[63044] <=  8'h74;        memory[63045] <=  8'h6b;        memory[63046] <=  8'h73;        memory[63047] <=  8'h68;        memory[63048] <=  8'h63;        memory[63049] <=  8'h66;        memory[63050] <=  8'h69;        memory[63051] <=  8'h77;        memory[63052] <=  8'h68;        memory[63053] <=  8'h61;        memory[63054] <=  8'h74;        memory[63055] <=  8'h61;        memory[63056] <=  8'h6e;        memory[63057] <=  8'h61;        memory[63058] <=  8'h62;        memory[63059] <=  8'h61;        memory[63060] <=  8'h63;        memory[63061] <=  8'h61;        memory[63062] <=  8'h74;        memory[63063] <=  8'h61;        memory[63064] <=  8'h62;        memory[63065] <=  8'h61;        memory[63066] <=  8'h72;        memory[63067] <=  8'h63;        memory[63068] <=  8'h61;        memory[63069] <=  8'h68;        memory[63070] <=  8'h64;        memory[63071] <=  8'h75;        memory[63072] <=  8'h63;        memory[63073] <=  8'h74;        memory[63074] <=  8'h61;        memory[63075] <=  8'h64;        memory[63076] <=  8'h61;        memory[63077] <=  8'h61;        memory[63078] <=  8'h63;        memory[63079] <=  8'h61;        memory[63080] <=  8'h72;        memory[63081] <=  8'h62;        memory[63082] <=  8'h61;        memory[63083] <=  8'h72;        memory[63084] <=  8'h74;        memory[63085] <=  8'h78;        memory[63086] <=  8'h61;        memory[63087] <=  8'h74;        memory[63088] <=  8'h6b;        memory[63089] <=  8'h73;        memory[63090] <=  8'h68;        memory[63091] <=  8'h63;        memory[63092] <=  8'h66;        memory[63093] <=  8'h69;        memory[63094] <=  8'h77;        memory[63095] <=  8'h68;        memory[63096] <=  8'h61;        memory[63097] <=  8'h74;        memory[63098] <=  8'h61;        memory[63099] <=  8'h6e;        memory[63100] <=  8'h61;        memory[63101] <=  8'h62;        memory[63102] <=  8'h61;        memory[63103] <=  8'h63;        memory[63104] <=  8'h61;        memory[63105] <=  8'h74;        memory[63106] <=  8'h61;        memory[63107] <=  8'h62;        memory[63108] <=  8'h61;        memory[63109] <=  8'h72;        memory[63110] <=  8'h63;        memory[63111] <=  8'h61;        memory[63112] <=  8'h68;        memory[63113] <=  8'h64;        memory[63114] <=  8'h75;        memory[63115] <=  8'h63;        memory[63116] <=  8'h74;        memory[63117] <=  8'h61;        memory[63118] <=  8'h64;        memory[63119] <=  8'h61;        memory[63120] <=  8'h61;        memory[63121] <=  8'h63;        memory[63122] <=  8'h61;        memory[63123] <=  8'h72;        memory[63124] <=  8'h62;        memory[63125] <=  8'h61;        memory[63126] <=  8'h72;        memory[63127] <=  8'h74;        memory[63128] <=  8'h78;        memory[63129] <=  8'h61;        memory[63130] <=  8'h74;        memory[63131] <=  8'h6b;        memory[63132] <=  8'h73;        memory[63133] <=  8'h68;        memory[63134] <=  8'h63;        memory[63135] <=  8'h66;        memory[63136] <=  8'h69;        memory[63137] <=  8'h77;        memory[63138] <=  8'h68;        memory[63139] <=  8'h61;        memory[63140] <=  8'h74;        memory[63141] <=  8'h61;        memory[63142] <=  8'h6e;        memory[63143] <=  8'h61;        memory[63144] <=  8'h62;        memory[63145] <=  8'h61;        memory[63146] <=  8'h63;        memory[63147] <=  8'h61;        memory[63148] <=  8'h74;        memory[63149] <=  8'h61;        memory[63150] <=  8'h62;        memory[63151] <=  8'h61;        memory[63152] <=  8'h72;        memory[63153] <=  8'h63;        memory[63154] <=  8'h61;        memory[63155] <=  8'h68;        memory[63156] <=  8'h64;        memory[63157] <=  8'h75;        memory[63158] <=  8'h63;        memory[63159] <=  8'h74;        memory[63160] <=  8'h61;        memory[63161] <=  8'h64;        memory[63162] <=  8'h61;        memory[63163] <=  8'h61;        memory[63164] <=  8'h63;        memory[63165] <=  8'h61;        memory[63166] <=  8'h72;        memory[63167] <=  8'h62;        memory[63168] <=  8'h61;        memory[63169] <=  8'h72;        memory[63170] <=  8'h74;        memory[63171] <=  8'h78;        memory[63172] <=  8'h61;        memory[63173] <=  8'h74;        memory[63174] <=  8'h6b;        memory[63175] <=  8'h73;        memory[63176] <=  8'h68;        memory[63177] <=  8'h63;        memory[63178] <=  8'h66;        memory[63179] <=  8'h69;        memory[63180] <=  8'h77;        memory[63181] <=  8'h68;        memory[63182] <=  8'h61;        memory[63183] <=  8'h74;        memory[63184] <=  8'h61;        memory[63185] <=  8'h6e;        memory[63186] <=  8'h61;        memory[63187] <=  8'h62;        memory[63188] <=  8'h61;        memory[63189] <=  8'h63;        memory[63190] <=  8'h61;        memory[63191] <=  8'h74;        memory[63192] <=  8'h61;        memory[63193] <=  8'h62;        memory[63194] <=  8'h61;        memory[63195] <=  8'h72;        memory[63196] <=  8'h63;        memory[63197] <=  8'h61;        memory[63198] <=  8'h68;        memory[63199] <=  8'h64;        memory[63200] <=  8'h75;        memory[63201] <=  8'h63;        memory[63202] <=  8'h74;        memory[63203] <=  8'h61;        memory[63204] <=  8'h64;        memory[63205] <=  8'h61;        memory[63206] <=  8'h61;        memory[63207] <=  8'h63;        memory[63208] <=  8'h61;        memory[63209] <=  8'h72;        memory[63210] <=  8'h62;        memory[63211] <=  8'h61;        memory[63212] <=  8'h72;        memory[63213] <=  8'h74;        memory[63214] <=  8'h78;        memory[63215] <=  8'h61;        memory[63216] <=  8'h74;        memory[63217] <=  8'h6b;        memory[63218] <=  8'h73;        memory[63219] <=  8'h68;        memory[63220] <=  8'h63;        memory[63221] <=  8'h66;        memory[63222] <=  8'h69;        memory[63223] <=  8'h77;        memory[63224] <=  8'h68;        memory[63225] <=  8'h61;        memory[63226] <=  8'h74;        memory[63227] <=  8'h61;        memory[63228] <=  8'h6e;        memory[63229] <=  8'h61;        memory[63230] <=  8'h62;        memory[63231] <=  8'h61;        memory[63232] <=  8'h63;        memory[63233] <=  8'h61;        memory[63234] <=  8'h74;        memory[63235] <=  8'h61;        memory[63236] <=  8'h62;        memory[63237] <=  8'h61;        memory[63238] <=  8'h72;        memory[63239] <=  8'h63;        memory[63240] <=  8'h61;        memory[63241] <=  8'h68;        memory[63242] <=  8'h64;        memory[63243] <=  8'h75;        memory[63244] <=  8'h63;        memory[63245] <=  8'h74;        memory[63246] <=  8'h61;        memory[63247] <=  8'h64;        memory[63248] <=  8'h61;        memory[63249] <=  8'h61;        memory[63250] <=  8'h63;        memory[63251] <=  8'h61;        memory[63252] <=  8'h72;        memory[63253] <=  8'h62;        memory[63254] <=  8'h61;        memory[63255] <=  8'h72;        memory[63256] <=  8'h74;        memory[63257] <=  8'h74;        memory[63258] <=  8'h62;        memory[63259] <=  8'h61;        memory[63260] <=  8'h72;        memory[63261] <=  8'h74;        memory[63262] <=  8'h78;        memory[63263] <=  8'h61;        memory[63264] <=  8'h74;        memory[63265] <=  8'h6b;        memory[63266] <=  8'h73;        memory[63267] <=  8'h68;        memory[63268] <=  8'h63;        memory[63269] <=  8'h66;        memory[63270] <=  8'h69;        memory[63271] <=  8'h77;        memory[63272] <=  8'h68;        memory[63273] <=  8'h61;        memory[63274] <=  8'h74;        memory[63275] <=  8'h61;        memory[63276] <=  8'h6e;        memory[63277] <=  8'h61;        memory[63278] <=  8'h62;        memory[63279] <=  8'h61;        memory[63280] <=  8'h63;        memory[63281] <=  8'h61;        memory[63282] <=  8'h74;        memory[63283] <=  8'h61;        memory[63284] <=  8'h62;        memory[63285] <=  8'h61;        memory[63286] <=  8'h72;        memory[63287] <=  8'h63;        memory[63288] <=  8'h61;        memory[63289] <=  8'h68;        memory[63290] <=  8'h64;        memory[63291] <=  8'h75;        memory[63292] <=  8'h63;        memory[63293] <=  8'h74;        memory[63294] <=  8'h61;        memory[63295] <=  8'h64;        memory[63296] <=  8'h61;        memory[63297] <=  8'h61;        memory[63298] <=  8'h63;        memory[63299] <=  8'h61;        memory[63300] <=  8'h72;        memory[63301] <=  8'h63;        memory[63302] <=  8'h74;        memory[63303] <=  8'h72;        memory[63304] <=  8'h63;        memory[63305] <=  8'h61;        memory[63306] <=  8'h74;        memory[63307] <=  8'h72;        memory[63308] <=  8'h63;        memory[63309] <=  8'h61;        memory[63310] <=  8'h74;        memory[63311] <=  8'h63;        memory[63312] <=  8'h62;        memory[63313] <=  8'h61;        memory[63314] <=  8'h74;        memory[63315] <=  8'h62;        memory[63316] <=  8'h72;        memory[63317] <=  8'h63;        memory[63318] <=  8'h61;        memory[63319] <=  8'h72;        memory[63320] <=  8'h62;        memory[63321] <=  8'h78;        memory[63322] <=  8'h74;        memory[63323] <=  8'h61;        memory[63324] <=  8'h72;        memory[63325] <=  8'h64;        memory[63326] <=  8'h66;        memory[63327] <=  8'h73;        memory[63328] <=  8'h67;        memory[63329] <=  8'h76;        memory[63330] <=  8'h68;        memory[63331] <=  8'h62;        memory[63332] <=  8'h6b;        memory[63333] <=  8'h6a;        memory[63334] <=  8'h6e;        memory[63335] <=  8'h6d;        memory[63336] <=  8'h62;        memory[63337] <=  8'h76;        memory[63338] <=  8'h78;        memory[63339] <=  8'h63;        memory[63340] <=  8'h73;        memory[63341] <=  8'h66;        memory[63342] <=  8'h72;        memory[63343] <=  8'h74;        memory[63344] <=  8'h79;        memory[63345] <=  8'h75;        memory[63346] <=  8'h6a;        memory[63347] <=  8'h6e;        memory[63348] <=  8'h62;        memory[63349] <=  8'h76;        memory[63350] <=  8'h63;        memory[63351] <=  8'h64;        memory[63352] <=  8'h74;        memory[63353] <=  8'h79;        memory[63354] <=  8'h75;        memory[63355] <=  8'h69;        memory[63356] <=  8'h6b;        memory[63357] <=  8'h6d;        memory[63358] <=  8'h6e;        memory[63359] <=  8'h62;        memory[63360] <=  8'h76;        memory[63361] <=  8'h63;        memory[63362] <=  8'h78;        memory[63363] <=  8'h73;        memory[63364] <=  8'h64;        memory[63365] <=  8'h72;        memory[63366] <=  8'h74;        memory[63367] <=  8'h79;        memory[63368] <=  8'h75;        memory[63369] <=  8'h69;        memory[63370] <=  8'h6b;        memory[63371] <=  8'h6d;        memory[63372] <=  8'h6e;        memory[63373] <=  8'h62;        memory[63374] <=  8'h76;        memory[63375] <=  8'h63;        memory[63376] <=  8'h73;        memory[63377] <=  8'h77;        memory[63378] <=  8'h33;        memory[63379] <=  8'h34;        memory[63380] <=  8'h35;        memory[63381] <=  8'h36;        memory[63382] <=  8'h37;        memory[63383] <=  8'h38;        memory[63384] <=  8'h69;        memory[63385] <=  8'h6b;        memory[63386] <=  8'h6d;        memory[63387] <=  8'h6e;        memory[63388] <=  8'h62;        memory[63389] <=  8'h76;        memory[63390] <=  8'h63;        memory[63391] <=  8'h64;        memory[63392] <=  8'h65;        memory[63393] <=  8'h72;        memory[63394] <=  8'h36;        memory[63395] <=  8'h37;        memory[63396] <=  8'h38;        memory[63397] <=  8'h69;        memory[63398] <=  8'h6f;        memory[63399] <=  8'h6b;        memory[63400] <=  8'h6a;        memory[63401] <=  8'h6e;        memory[63402] <=  8'h62;        memory[63403] <=  8'h76;        memory[63404] <=  8'h63;        memory[63405] <=  8'h64;        memory[63406] <=  8'h72;        memory[63407] <=  8'h74;        memory[63408] <=  8'h79;        memory[63409] <=  8'h75;        memory[63410] <=  8'h73;        memory[63411] <=  8'h6a;        memory[63412] <=  8'h63;        memory[63413] <=  8'h6e;        memory[63414] <=  8'h62;        memory[63415] <=  8'h64;        memory[63416] <=  8'h66;        memory[63417] <=  8'h73;        memory[63418] <=  8'h74;        memory[63419] <=  8'h79;        memory[63420] <=  8'h75;        memory[63421] <=  8'h61;        memory[63422] <=  8'h69;        memory[63423] <=  8'h6b;        memory[63424] <=  8'h78;        memory[63425] <=  8'h6d;        memory[63426] <=  8'h6e;        memory[63427] <=  8'h73;        memory[63428] <=  8'h6a;        memory[63429] <=  8'h6f;        memory[63430] <=  8'h64;        memory[63431] <=  8'h6c;        memory[63432] <=  8'h63;        memory[63433] <=  8'h78;        memory[63434] <=  8'h2c;        memory[63435] <=  8'h6d;        memory[63436] <=  8'h73;        memory[63437] <=  8'h6b;        memory[63438] <=  8'h64;        memory[63439] <=  8'h6c;        memory[63440] <=  8'h70;        memory[63441] <=  8'h5b;        memory[63442] <=  8'h3b;        memory[63443] <=  8'h73;        memory[63444] <=  8'h6c;        memory[63445] <=  8'h64;        memory[63446] <=  8'h70;        memory[63447] <=  8'h76;        memory[63448] <=  8'h63;        memory[63449] <=  8'h5b;        memory[63450] <=  8'h78;        memory[63451] <=  8'h76;        memory[63452] <=  8'h63;        memory[63453] <=  8'h5b;        memory[63454] <=  8'h78;        memory[63455] <=  8'h70;        memory[63456] <=  8'h6f;        memory[63457] <=  8'h20;        memory[63458] <=  8'h62;        memory[63459] <=  8'h61;        memory[63460] <=  8'h72;        memory[63461] <=  8'h74;        memory[63462] <=  8'h74;        memory[63463] <=  8'h62;        memory[63464] <=  8'h61;        memory[63465] <=  8'h72;        memory[63466] <=  8'h74;        memory[63467] <=  8'h78;        memory[63468] <=  8'h61;        memory[63469] <=  8'h74;        memory[63470] <=  8'h6b;        memory[63471] <=  8'h73;        memory[63472] <=  8'h68;        memory[63473] <=  8'h63;        memory[63474] <=  8'h66;        memory[63475] <=  8'h69;        memory[63476] <=  8'h77;        memory[63477] <=  8'h68;        memory[63478] <=  8'h61;        memory[63479] <=  8'h69;        memory[63480] <=  8'h6a;        memory[63481] <=  8'h78;        memory[63482] <=  8'h5d;        memory[63483] <=  8'h65;        memory[63484] <=  8'h6b;        memory[63485] <=  8'h6f;        memory[63486] <=  8'h39;        memory[63487] <=  8'h64;        memory[63488] <=  8'h75;        memory[63489] <=  8'h38;        memory[63490] <=  8'h79;        memory[63491] <=  8'h20;        memory[63492] <=  8'h37;        memory[63493] <=  8'h63;        memory[63494] <=  8'h67;        memory[63495] <=  8'h78;        memory[63496] <=  8'h63;        memory[63497] <=  8'h75;        memory[63498] <=  8'h68;        memory[63499] <=  8'h69;        memory[63500] <=  8'h6a;        memory[63501] <=  8'h77;        memory[63502] <=  8'h69;        memory[63503] <=  8'h64;        memory[63504] <=  8'h66;        memory[63505] <=  8'h68;        memory[63506] <=  8'h75;        memory[63507] <=  8'h76;        memory[63508] <=  8'h64;        memory[63509] <=  8'h62;        memory[63510] <=  8'h66;        memory[63511] <=  8'h6a;        memory[63512] <=  8'h6e;        memory[63513] <=  8'h6b;        memory[63514] <=  8'h6a;        memory[63515] <=  8'h65;        memory[63516] <=  8'h38;        memory[63517] <=  8'h66;        memory[63518] <=  8'h37;        memory[63519] <=  8'h67;        memory[63520] <=  8'h79;        memory[63521] <=  8'h76;        memory[63522] <=  8'h63;        memory[63523] <=  8'h68;        memory[63524] <=  8'h69;        memory[63525] <=  8'h6a;        memory[63526] <=  8'h33;        memory[63527] <=  8'h65;        memory[63528] <=  8'h67;        memory[63529] <=  8'h79;        memory[63530] <=  8'h72;        memory[63531] <=  8'h64;        memory[63532] <=  8'h62;        memory[63533] <=  8'h6e;        memory[63534] <=  8'h63;        memory[63535] <=  8'h7a;        memory[63536] <=  8'h6a;        memory[63537] <=  8'h6f;        memory[63538] <=  8'h66;        memory[63539] <=  8'h78;        memory[63540] <=  8'h6a;        memory[63541] <=  8'h69;        memory[63542] <=  8'h63;        memory[63543] <=  8'h68;        memory[63544] <=  8'h62;        memory[63545] <=  8'h6e;        memory[63546] <=  8'h6d;        memory[63547] <=  8'h63;        memory[63548] <=  8'h73;        memory[63549] <=  8'h6c;        memory[63550] <=  8'h6b;        memory[63551] <=  8'h6a;        memory[63552] <=  8'h69;        memory[63553] <=  8'h68;        memory[63554] <=  8'h76;        memory[63555] <=  8'h75;        memory[63556] <=  8'h69;        memory[63557] <=  8'h64;        memory[63558] <=  8'h68;        memory[63559] <=  8'h75;        memory[63560] <=  8'h67;        memory[63561] <=  8'h79;        memory[63562] <=  8'h62;        memory[63563] <=  8'h68;        memory[63564] <=  8'h65;        memory[63565] <=  8'h6a;        memory[63566] <=  8'h72;        memory[63567] <=  8'h6b;        memory[63568] <=  8'h6a;        memory[63569] <=  8'h6f;        memory[63570] <=  8'h64;        memory[63571] <=  8'h67;        memory[63572] <=  8'h69;        memory[63573] <=  8'h75;        memory[63574] <=  8'h69;        memory[63575] <=  8'h67;        memory[63576] <=  8'h76;        memory[63577] <=  8'h79;        memory[63578] <=  8'h75;        memory[63579] <=  8'h67;        memory[63580] <=  8'h78;        memory[63581] <=  8'h68;        memory[63582] <=  8'h63;        memory[63583] <=  8'h20;        memory[63584] <=  8'h20;        memory[63585] <=  8'h20;        memory[63586] <=  8'h78;        memory[63587] <=  8'h76;        memory[63588] <=  8'h20;        memory[63589] <=  8'h63;        memory[63590] <=  8'h78;        memory[63591] <=  8'h67;        memory[63592] <=  8'h79;        memory[63593] <=  8'h63;        memory[63594] <=  8'h75;        memory[63595] <=  8'h68;        memory[63596] <=  8'h6a;        memory[63597] <=  8'h6b;        memory[63598] <=  8'h61;        memory[63599] <=  8'h6c;        memory[63600] <=  8'h78;        memory[63601] <=  8'h76;        memory[63602] <=  8'h70;        memory[63603] <=  8'h6f;        memory[63604] <=  8'h69;        memory[63605] <=  8'h6a;        memory[63606] <=  8'h69;        memory[63607] <=  8'h68;        memory[63608] <=  8'h6a;        memory[63609] <=  8'h62;        memory[63610] <=  8'h77;        memory[63611] <=  8'h65;        memory[63612] <=  8'h6e;        memory[63613] <=  8'h61;        memory[63614] <=  8'h66;        memory[63615] <=  8'h6d;        memory[63616] <=  8'h64;        memory[63617] <=  8'h6b;        memory[63618] <=  8'h6d;        memory[63619] <=  8'h76;        memory[63620] <=  8'h6c;        memory[63621] <=  8'h63;        memory[63622] <=  8'h6f;        memory[63623] <=  8'h64;        memory[63624] <=  8'h69;        memory[63625] <=  8'h75;        memory[63626] <=  8'h68;        memory[63627] <=  8'h73;        memory[63628] <=  8'h66;        memory[63629] <=  8'h65;        memory[63630] <=  8'h62;        memory[63631] <=  8'h6e;        memory[63632] <=  8'h64;        memory[63633] <=  8'h73;        memory[63634] <=  8'h63;        memory[63635] <=  8'h6b;        memory[63636] <=  8'h20;        memory[63637] <=  8'h78;        memory[63638] <=  8'h6a;        memory[63639] <=  8'h78;        memory[63640] <=  8'h63;        memory[63641] <=  8'h73;        memory[63642] <=  8'h64;        memory[63643] <=  8'h66;        memory[63644] <=  8'h6b;        memory[63645] <=  8'h64;        memory[63646] <=  8'h6e;        memory[63647] <=  8'h6d;        memory[63648] <=  8'h64;        memory[63649] <=  8'h73;        memory[63650] <=  8'h63;        memory[63651] <=  8'h6b;        memory[63652] <=  8'h78;        memory[63653] <=  8'h6c;        memory[63654] <=  8'h6f;        memory[63655] <=  8'h66;        memory[63656] <=  8'h6a;        memory[63657] <=  8'h69;        memory[63658] <=  8'h61;        memory[63659] <=  8'h62;        memory[63660] <=  8'h6e;        memory[63661] <=  8'h20;        memory[63662] <=  8'h78;        memory[63663] <=  8'h6b;        memory[63664] <=  8'h6d;        memory[63665] <=  8'h20;        memory[63666] <=  8'h6f;        memory[63667] <=  8'h63;        memory[63668] <=  8'h76;        memory[63669] <=  8'h73;        memory[63670] <=  8'h64;        memory[63671] <=  8'h69;        memory[63672] <=  8'h66;        memory[63673] <=  8'h68;        memory[63674] <=  8'h65;        memory[63675] <=  8'h71;        memory[63676] <=  8'h6a;        memory[63677] <=  8'h77;        memory[63678] <=  8'h62;        memory[63679] <=  8'h65;        memory[63680] <=  8'h6e;        memory[63681] <=  8'h20;        memory[63682] <=  8'h6d;        memory[63683] <=  8'h64;        memory[63684] <=  8'h73;        memory[63685] <=  8'h6c;        memory[63686] <=  8'h76;        memory[63687] <=  8'h6b;        memory[63688] <=  8'h63;        memory[63689] <=  8'h78;        memory[63690] <=  8'h20;        memory[63691] <=  8'h6f;        memory[63692] <=  8'h78;        memory[63693] <=  8'h69;        memory[63694] <=  8'h63;        memory[63695] <=  8'h6a;        memory[63696] <=  8'h76;        memory[63697] <=  8'h64;        memory[63698] <=  8'h66;        memory[63699] <=  8'h65;        memory[63700] <=  8'h71;        memory[63701] <=  8'h6e;        memory[63702] <=  8'h20;        memory[63703] <=  8'h64;        memory[63704] <=  8'h6d;        memory[63705] <=  8'h73;        memory[63706] <=  8'h6c;        memory[63707] <=  8'h63;        memory[63708] <=  8'h78;        memory[63709] <=  8'h6b;        memory[63710] <=  8'h20;        memory[63711] <=  8'h6f;        memory[63712] <=  8'h78;        memory[63713] <=  8'h63;        memory[63714] <=  8'h76;        memory[63715] <=  8'h6a;        memory[63716] <=  8'h64;        memory[63717] <=  8'h62;        memory[63718] <=  8'h71;        memory[63719] <=  8'h77;        memory[63720] <=  8'h65;        memory[63721] <=  8'h6e;        memory[63722] <=  8'h6d;        memory[63723] <=  8'h64;        memory[63724] <=  8'h6c;        memory[63725] <=  8'h73;        memory[63726] <=  8'h2c;        memory[63727] <=  8'h76;        memory[63728] <=  8'h63;        memory[63729] <=  8'h78;        memory[63730] <=  8'h20;        memory[63731] <=  8'h63;        memory[63732] <=  8'h6f;        memory[63733] <=  8'h69;        memory[63734] <=  8'h76;        memory[63735] <=  8'h68;        memory[63736] <=  8'h73;        memory[63737] <=  8'h64;        memory[63738] <=  8'h62;        memory[63739] <=  8'h71;        memory[63740] <=  8'h77;        memory[63741] <=  8'h65;        memory[63742] <=  8'h6e;        memory[63743] <=  8'h64;        memory[63744] <=  8'h6b;        memory[63745] <=  8'h73;        memory[63746] <=  8'h76;        memory[63747] <=  8'h6f;        memory[63748] <=  8'h63;        memory[63749] <=  8'h20;        memory[63750] <=  8'h76;        memory[63751] <=  8'h69;        memory[63752] <=  8'h75;        memory[63753] <=  8'h69;        memory[63754] <=  8'h68;        memory[63755] <=  8'h63;        memory[63756] <=  8'h78;        memory[63757] <=  8'h69;        memory[63758] <=  8'h6f;        memory[63759] <=  8'h76;        memory[63760] <=  8'h73;        memory[63761] <=  8'h64;        memory[63762] <=  8'h61;        memory[63763] <=  8'h64;        memory[63764] <=  8'h6e;        memory[63765] <=  8'h77;        memory[63766] <=  8'h71;        memory[63767] <=  8'h6b;        memory[63768] <=  8'h6c;        memory[63769] <=  8'h73;        memory[63770] <=  8'h76;        memory[63771] <=  8'h6e;        memory[63772] <=  8'h62;        memory[63773] <=  8'h20;        memory[63774] <=  8'h64;        memory[63775] <=  8'h66;        memory[63776] <=  8'h6a;        memory[63777] <=  8'h6b;        memory[63778] <=  8'h71;        memory[63779] <=  8'h64;        memory[63780] <=  8'h77;        memory[63781] <=  8'h65;        memory[63782] <=  8'h6e;        memory[63783] <=  8'h62;        memory[63784] <=  8'h20;        memory[63785] <=  8'h64;        memory[63786] <=  8'h73;        memory[63787] <=  8'h76;        memory[63788] <=  8'h68;        memory[63789] <=  8'h64;        memory[63790] <=  8'h61;        memory[63791] <=  8'h71;        memory[63792] <=  8'h77;        memory[63793] <=  8'h6a;        memory[63794] <=  8'h65;        memory[63795] <=  8'h6e;        memory[63796] <=  8'h64;        memory[63797] <=  8'h20;        memory[63798] <=  8'h61;        memory[63799] <=  8'h63;        memory[63800] <=  8'h62;        memory[63801] <=  8'h68;        memory[63802] <=  8'h64;        memory[63803] <=  8'h61;        memory[63804] <=  8'h77;        memory[63805] <=  8'h71;        memory[63806] <=  8'h6e;        memory[63807] <=  8'h20;        memory[63808] <=  8'h62;        memory[63809] <=  8'h73;        memory[63810] <=  8'h76;        memory[63811] <=  8'h61;        memory[63812] <=  8'h67;        memory[63813] <=  8'h76;        memory[63814] <=  8'h68;        memory[63815] <=  8'h67;        memory[63816] <=  8'h61;        memory[63817] <=  8'h73;        memory[63818] <=  8'h6a;        memory[63819] <=  8'h6b;        memory[63820] <=  8'h63;        memory[63821] <=  8'h78;        memory[63822] <=  8'h76;        memory[63823] <=  8'h6e;        memory[63824] <=  8'h73;        memory[63825] <=  8'h64;        memory[63826] <=  8'h20;        memory[63827] <=  8'h66;        memory[63828] <=  8'h62;        memory[63829] <=  8'h64;        memory[63830] <=  8'h61;        memory[63831] <=  8'h73;        memory[63832] <=  8'h76;        memory[63833] <=  8'h67;        memory[63834] <=  8'h63;        memory[63835] <=  8'h79;        memory[63836] <=  8'h7a;        memory[63837] <=  8'h78;        memory[63838] <=  8'h79;        memory[63839] <=  8'h75;        memory[63840] <=  8'h20;        memory[63841] <=  8'h69;        memory[63842] <=  8'h6a;        memory[63843] <=  8'h64;        memory[63844] <=  8'h66;        memory[63845] <=  8'h6b;        memory[63846] <=  8'h61;        memory[63847] <=  8'h64;        memory[63848] <=  8'h63;        memory[63849] <=  8'h78;        memory[63850] <=  8'h68;        memory[63851] <=  8'h20;        memory[63852] <=  8'h67;        memory[63853] <=  8'h61;        memory[63854] <=  8'h68;        memory[63855] <=  8'h75;        memory[63856] <=  8'h64;        memory[63857] <=  8'h73;        memory[63858] <=  8'h69;        memory[63859] <=  8'h6a;        memory[63860] <=  8'h61;        memory[63861] <=  8'h6b;        memory[63862] <=  8'h63;        memory[63863] <=  8'h62;        memory[63864] <=  8'h61;        memory[63865] <=  8'h72;        memory[63866] <=  8'h73;        memory[63867] <=  8'h68;        memory[63868] <=  8'h64;        memory[63869] <=  8'h66;        memory[63870] <=  8'h67;        memory[63871] <=  8'h73;        memory[63872] <=  8'h68;        memory[63873] <=  8'h64;        memory[63874] <=  8'h66;        memory[63875] <=  8'h68;        memory[63876] <=  8'h64;        memory[63877] <=  8'h6a;        memory[63878] <=  8'h68;        memory[63879] <=  8'h62;        memory[63880] <=  8'h67;        memory[63881] <=  8'h63;        memory[63882] <=  8'h61;        memory[63883] <=  8'h66;        memory[63884] <=  8'h73;        memory[63885] <=  8'h79;        memory[63886] <=  8'h67;        memory[63887] <=  8'h6b;        memory[63888] <=  8'h75;        memory[63889] <=  8'h64;        memory[63890] <=  8'h68;        memory[63891] <=  8'h62;        memory[63892] <=  8'h77;        memory[63893] <=  8'h76;        memory[63894] <=  8'h67;        memory[63895] <=  8'h61;        memory[63896] <=  8'h66;        memory[63897] <=  8'h64;        memory[63898] <=  8'h74;        memory[63899] <=  8'h75;        memory[63900] <=  8'h66;        memory[63901] <=  8'h79;        memory[63902] <=  8'h67;        memory[63903] <=  8'h69;        memory[63904] <=  8'h75;        memory[63905] <=  8'h68;        memory[63906] <=  8'h6c;        memory[63907] <=  8'h6a;        memory[63908] <=  8'h62;        memory[63909] <=  8'h6b;        memory[63910] <=  8'h68;        memory[63911] <=  8'h76;        memory[63912] <=  8'h67;        memory[63913] <=  8'h63;        memory[63914] <=  8'h66;        memory[63915] <=  8'h78;        memory[63916] <=  8'h64;        memory[63917] <=  8'h74;        memory[63918] <=  8'h75;        memory[63919] <=  8'h79;        memory[63920] <=  8'h69;        memory[63921] <=  8'h75;        memory[63922] <=  8'h68;        memory[63923] <=  8'h6c;        memory[63924] <=  8'h6a;        memory[63925] <=  8'h6b;        memory[63926] <=  8'h67;        memory[63927] <=  8'h6a;        memory[63928] <=  8'h63;        memory[63929] <=  8'h66;        memory[63930] <=  8'h68;        memory[63931] <=  8'h64;        memory[63932] <=  8'h67;        memory[63933] <=  8'h72;        memory[63934] <=  8'h79;        memory[63935] <=  8'h74;        memory[63936] <=  8'h66;        memory[63937] <=  8'h75;        memory[63938] <=  8'h79;        memory[63939] <=  8'h69;        memory[63940] <=  8'h68;        memory[63941] <=  8'h6c;        memory[63942] <=  8'h62;        memory[63943] <=  8'h6d;        memory[63944] <=  8'h76;        memory[63945] <=  8'h6e;        memory[63946] <=  8'h63;        memory[63947] <=  8'h66;        memory[63948] <=  8'h68;        memory[63949] <=  8'h64;        memory[63950] <=  8'h74;        memory[63951] <=  8'h75;        memory[63952] <=  8'h67;        memory[63953] <=  8'h79;        memory[63954] <=  8'h69;        memory[63955] <=  8'h68;        memory[63956] <=  8'h75;        memory[63957] <=  8'h6a;        memory[63958] <=  8'h6c;        memory[63959] <=  8'h62;        memory[63960] <=  8'h6d;        memory[63961] <=  8'h76;        memory[63962] <=  8'h6e;        memory[63963] <=  8'h63;        memory[63964] <=  8'h66;        memory[63965] <=  8'h68;        memory[63966] <=  8'h67;        memory[63967] <=  8'h79;        memory[63968] <=  8'h68;        memory[63969] <=  8'h75;        memory[63970] <=  8'h6a;        memory[63971] <=  8'h6e;        memory[63972] <=  8'h2c;        memory[63973] <=  8'h62;        memory[63974] <=  8'h6e;        memory[63975] <=  8'h6d;        memory[63976] <=  8'h76;        memory[63977] <=  8'h6e;        memory[63978] <=  8'h63;        memory[63979] <=  8'h66;        memory[63980] <=  8'h68;        memory[63981] <=  8'h74;        memory[63982] <=  8'h79;        memory[63983] <=  8'h69;        memory[63984] <=  8'h75;        memory[63985] <=  8'h6c;        memory[63986] <=  8'h6a;        memory[63987] <=  8'h62;        memory[63988] <=  8'h6d;        memory[63989] <=  8'h76;        memory[63990] <=  8'h6e;        memory[63991] <=  8'h63;        memory[63992] <=  8'h66;        memory[63993] <=  8'h74;        memory[63994] <=  8'h75;        memory[63995] <=  8'h79;        memory[63996] <=  8'h69;        memory[63997] <=  8'h68;        memory[63998] <=  8'h6b;        memory[63999] <=  8'h62;        memory[64000] <=  8'h76;        memory[64001] <=  8'h63;        memory[64002] <=  8'h66;        memory[64003] <=  8'h67;        memory[64004] <=  8'h74;        memory[64005] <=  8'h75;        memory[64006] <=  8'h79;        memory[64007] <=  8'h69;        memory[64008] <=  8'h75;        memory[64009] <=  8'h68;        memory[64010] <=  8'h6a;        memory[64011] <=  8'h6b;        memory[64012] <=  8'h62;        memory[64013] <=  8'h76;        memory[64014] <=  8'h63;        memory[64015] <=  8'h66;        memory[64016] <=  8'h74;        memory[64017] <=  8'h75;        memory[64018] <=  8'h79;        memory[64019] <=  8'h69;        memory[64020] <=  8'h75;        memory[64021] <=  8'h6a;        memory[64022] <=  8'h6b;        memory[64023] <=  8'h6e;        memory[64024] <=  8'h62;        memory[64025] <=  8'h76;        memory[64026] <=  8'h67;        memory[64027] <=  8'h66;        memory[64028] <=  8'h74;        memory[64029] <=  8'h79;        memory[64030] <=  8'h75;        memory[64031] <=  8'h75;        memory[64032] <=  8'h69;        memory[64033] <=  8'h6a;        memory[64034] <=  8'h6b;        memory[64035] <=  8'h68;        memory[64036] <=  8'h62;        memory[64037] <=  8'h6a;        memory[64038] <=  8'h67;        memory[64039] <=  8'h68;        memory[64040] <=  8'h66;        memory[64041] <=  8'h79;        memory[64042] <=  8'h74;        memory[64043] <=  8'h79;        memory[64044] <=  8'h69;        memory[64045] <=  8'h75;        memory[64046] <=  8'h64;        memory[64047] <=  8'h6a;        memory[64048] <=  8'h6b;        memory[64049] <=  8'h68;        memory[64050] <=  8'h63;        memory[64051] <=  8'h7a;        memory[64052] <=  8'h67;        memory[64053] <=  8'h68;        memory[64054] <=  8'h74;        memory[64055] <=  8'h75;        memory[64056] <=  8'h79;        memory[64057] <=  8'h69;        memory[64058] <=  8'h61;        memory[64059] <=  8'h73;        memory[64060] <=  8'h75;        memory[64061] <=  8'h6a;        memory[64062] <=  8'h6b;        memory[64063] <=  8'h62;        memory[64064] <=  8'h6e;        memory[64065] <=  8'h61;        memory[64066] <=  8'h76;        memory[64067] <=  8'h63;        memory[64068] <=  8'h66;        memory[64069] <=  8'h68;        memory[64070] <=  8'h75;        memory[64071] <=  8'h61;        memory[64072] <=  8'h73;        memory[64073] <=  8'h79;        memory[64074] <=  8'h64;        memory[64075] <=  8'h75;        memory[64076] <=  8'h69;        memory[64077] <=  8'h6a;        memory[64078] <=  8'h61;        memory[64079] <=  8'h6b;        memory[64080] <=  8'h62;        memory[64081] <=  8'h63;        memory[64082] <=  8'h78;        memory[64083] <=  8'h68;        memory[64084] <=  8'h67;        memory[64085] <=  8'h79;        memory[64086] <=  8'h75;        memory[64087] <=  8'h7a;        memory[64088] <=  8'h63;        memory[64089] <=  8'h61;        memory[64090] <=  8'h73;        memory[64091] <=  8'h69;        memory[64092] <=  8'h75;        memory[64093] <=  8'h6f;        memory[64094] <=  8'h69;        memory[64095] <=  8'h6a;        memory[64096] <=  8'h61;        memory[64097] <=  8'h6c;        memory[64098] <=  8'h63;        memory[64099] <=  8'h78;        memory[64100] <=  8'h62;        memory[64101] <=  8'h63;        memory[64102] <=  8'h20;        memory[64103] <=  8'h6e;        memory[64104] <=  8'h76;        memory[64105] <=  8'h63;        memory[64106] <=  8'h61;        memory[64107] <=  8'h64;        memory[64108] <=  8'h73;        memory[64109] <=  8'h67;        memory[64110] <=  8'h79;        memory[64111] <=  8'h68;        memory[64112] <=  8'h75;        memory[64113] <=  8'h61;        memory[64114] <=  8'h6a;        memory[64115] <=  8'h6b;        memory[64116] <=  8'h78;        memory[64117] <=  8'h62;        memory[64118] <=  8'h20;        memory[64119] <=  8'h6e;        memory[64120] <=  8'h76;        memory[64121] <=  8'h63;        memory[64122] <=  8'h61;        memory[64123] <=  8'h73;        memory[64124] <=  8'h67;        memory[64125] <=  8'h68;        memory[64126] <=  8'h75;        memory[64127] <=  8'h6a;        memory[64128] <=  8'h6c;        memory[64129] <=  8'h6b;        memory[64130] <=  8'h63;        memory[64131] <=  8'h78;        memory[64132] <=  8'h20;        memory[64133] <=  8'h6a;        memory[64134] <=  8'h6b;        memory[64135] <=  8'h68;        memory[64136] <=  8'h61;        memory[64137] <=  8'h73;        memory[64138] <=  8'h76;        memory[64139] <=  8'h64;        memory[64140] <=  8'h6e;        memory[64141] <=  8'h20;        memory[64142] <=  8'h62;        memory[64143] <=  8'h6e;        memory[64144] <=  8'h6d;        memory[64145] <=  8'h6b;        memory[64146] <=  8'h77;        memory[64147] <=  8'h64;        memory[64148] <=  8'h6f;        memory[64149] <=  8'h77;        memory[64150] <=  8'h69;        memory[64151] <=  8'h6f;        memory[64152] <=  8'h75;        memory[64153] <=  8'h69;        memory[64154] <=  8'h68;        memory[64155] <=  8'h62;        memory[64156] <=  8'h6e;        memory[64157] <=  8'h6b;        memory[64158] <=  8'h77;        memory[64159] <=  8'h69;        memory[64160] <=  8'h6f;        memory[64161] <=  8'h75;        memory[64162] <=  8'h71;        memory[64163] <=  8'h69;        memory[64164] <=  8'h79;        memory[64165] <=  8'h67;        memory[64166] <=  8'h6a;        memory[64167] <=  8'h64;        memory[64168] <=  8'h61;        memory[64169] <=  8'h76;        memory[64170] <=  8'h62;        memory[64171] <=  8'h6e;        memory[64172] <=  8'h6b;        memory[64173] <=  8'h6f;        memory[64174] <=  8'h70;        memory[64175] <=  8'h64;        memory[64176] <=  8'h76;        memory[64177] <=  8'h69;        memory[64178] <=  8'h6f;        memory[64179] <=  8'h75;        memory[64180] <=  8'h69;        memory[64181] <=  8'h48;        memory[64182] <=  8'h42;        memory[64183] <=  8'h6b;        memory[64184] <=  8'h64;        memory[64185] <=  8'h6e;        memory[64186] <=  8'h6c;        memory[64187] <=  8'h71;        memory[64188] <=  8'h6b;        memory[64189] <=  8'h6d;        memory[64190] <=  8'h6a;        memory[64191] <=  8'h70;        memory[64192] <=  8'h69;        memory[64193] <=  8'h6f;        memory[64194] <=  8'h68;        memory[64195] <=  8'h65;        memory[64196] <=  8'h66;        memory[64197] <=  8'h75;        memory[64198] <=  8'h67;        memory[64199] <=  8'h69;        memory[64200] <=  8'h73;        memory[64201] <=  8'h61;        memory[64202] <=  8'h62;        memory[64203] <=  8'h64;        memory[64204] <=  8'h6b;        memory[64205] <=  8'h6a;        memory[64206] <=  8'h6b;        memory[64207] <=  8'h6c;        memory[64208] <=  8'h6a;        memory[64209] <=  8'h69;        memory[64210] <=  8'h73;        memory[64211] <=  8'h6f;        memory[64212] <=  8'h71;        memory[64213] <=  8'h68;        memory[64214] <=  8'h77;        memory[64215] <=  8'h67;        memory[64216] <=  8'h69;        memory[64217] <=  8'h79;        memory[64218] <=  8'h6a;        memory[64219] <=  8'h64;        memory[64220] <=  8'h76;        memory[64221] <=  8'h62;        memory[64222] <=  8'h6e;        memory[64223] <=  8'h61;        memory[64224] <=  8'h73;        memory[64225] <=  8'h66;        memory[64226] <=  8'h6c;        memory[64227] <=  8'h6b;        memory[64228] <=  8'h64;        memory[64229] <=  8'h6a;        memory[64230] <=  8'h68;        memory[64231] <=  8'h63;        memory[64232] <=  8'h67;        memory[64233] <=  8'h6a;        memory[64234] <=  8'h76;        memory[64235] <=  8'h73;        memory[64236] <=  8'h64;        memory[64237] <=  8'h62;        memory[64238] <=  8'h62;        memory[64239] <=  8'h61;        memory[64240] <=  8'h72;        memory[64241] <=  8'h62;        memory[64242] <=  8'h62;        memory[64243] <=  8'h73;        memory[64244] <=  8'h62;        memory[64245] <=  8'h67;        memory[64246] <=  8'h73;        memory[64247] <=  8'h66;        memory[64248] <=  8'h67;        memory[64249] <=  8'h61;        memory[64250] <=  8'h68;        memory[64251] <=  8'h66;        memory[64252] <=  8'h73;        memory[64253] <=  8'h68;        memory[64254] <=  8'h61;        memory[64255] <=  8'h66;        memory[64256] <=  8'h73;        memory[64257] <=  8'h66;        memory[64258] <=  8'h68;        memory[64259] <=  8'h61;        memory[64260] <=  8'h69;        memory[64261] <=  8'h64;        memory[64262] <=  8'h75;        memory[64263] <=  8'h67;        memory[64264] <=  8'h64;        memory[64265] <=  8'h77;        memory[64266] <=  8'h62;        memory[64267] <=  8'h61;        memory[64268] <=  8'h62;        memory[64269] <=  8'h72;        memory[64270] <=  8'h62;        memory[64271] <=  8'h61;        memory[64272] <=  8'h62;        memory[64273] <=  8'h62;        memory[64274] <=  8'h74;        memory[64275] <=  8'h62;        memory[64276] <=  8'h62;        memory[64277] <=  8'h62;        memory[64278] <=  8'h62;        memory[64279] <=  8'h62;        memory[64280] <=  8'h62;        memory[64281] <=  8'h62;        memory[64282] <=  8'h62;        memory[64283] <=  8'h61;        memory[64284] <=  8'h62;        memory[64285] <=  8'h62;        memory[64286] <=  8'h72;        memory[64287] <=  8'h74;        memory[64288] <=  8'h62;        memory[64289] <=  8'h62;        memory[64290] <=  8'h61;        memory[64291] <=  8'h62;        memory[64292] <=  8'h72;        memory[64293] <=  8'h62;        memory[64294] <=  8'h74;        memory[64295] <=  8'h62;        memory[64296] <=  8'h62;        memory[64297] <=  8'h62;        memory[64298] <=  8'h63;        memory[64299] <=  8'h61;        memory[64300] <=  8'h72;        memory[64301] <=  8'h74;        memory[64302] <=  8'h73;        memory[64303] <=  8'h62;        memory[64304] <=  8'h61;        memory[64305] <=  8'h72;        memory[64306] <=  8'h74;        memory[64307] <=  8'h74;        memory[64308] <=  8'h62;        memory[64309] <=  8'h61;        memory[64310] <=  8'h72;        memory[64311] <=  8'h74;        memory[64312] <=  8'h78;        memory[64313] <=  8'h61;        memory[64314] <=  8'h74;        memory[64315] <=  8'h6b;        memory[64316] <=  8'h73;        memory[64317] <=  8'h68;        memory[64318] <=  8'h63;        memory[64319] <=  8'h66;        memory[64320] <=  8'h69;        memory[64321] <=  8'h77;        memory[64322] <=  8'h68;        memory[64323] <=  8'h61;        memory[64324] <=  8'h74;        memory[64325] <=  8'h61;        memory[64326] <=  8'h6e;        memory[64327] <=  8'h61;        memory[64328] <=  8'h62;        memory[64329] <=  8'h61;        memory[64330] <=  8'h63;        memory[64331] <=  8'h61;        memory[64332] <=  8'h74;        memory[64333] <=  8'h61;        memory[64334] <=  8'h62;        memory[64335] <=  8'h61;        memory[64336] <=  8'h72;        memory[64337] <=  8'h63;        memory[64338] <=  8'h61;        memory[64339] <=  8'h68;        memory[64340] <=  8'h64;        memory[64341] <=  8'h75;        memory[64342] <=  8'h63;        memory[64343] <=  8'h74;        memory[64344] <=  8'h61;        memory[64345] <=  8'h64;        memory[64346] <=  8'h61;        memory[64347] <=  8'h61;        memory[64348] <=  8'h63;        memory[64349] <=  8'h61;        memory[64350] <=  8'h72;        memory[64351] <=  8'h63;        memory[64352] <=  8'h74;        memory[64353] <=  8'h72;        memory[64354] <=  8'h63;        memory[64355] <=  8'h61;        memory[64356] <=  8'h74;        memory[64357] <=  8'h72;        memory[64358] <=  8'h63;        memory[64359] <=  8'h61;        memory[64360] <=  8'h74;        memory[64361] <=  8'h63;        memory[64362] <=  8'h62;        memory[64363] <=  8'h61;        memory[64364] <=  8'h74;        memory[64365] <=  8'h62;        memory[64366] <=  8'h72;        memory[64367] <=  8'h63;        memory[64368] <=  8'h61;        memory[64369] <=  8'h74;        memory[64370] <=  8'h72;        memory[64371] <=  8'h6e;        memory[64372] <=  8'h62;        memory[64373] <=  8'h61;        memory[64374] <=  8'h63;        memory[64375] <=  8'h61;        memory[64376] <=  8'h74;        memory[64377] <=  8'h79;        memory[64378] <=  8'h73;        memory[64379] <=  8'h6e;        memory[64380] <=  8'h63;        memory[64381] <=  8'h74;        memory[64382] <=  8'h61;        memory[64383] <=  8'h6e;        memory[64384] <=  8'h62;        memory[64385] <=  8'h61;        memory[64386] <=  8'h63;        memory[64387] <=  8'h72;        memory[64388] <=  8'h6e;        memory[64389] <=  8'h74;        memory[64390] <=  8'h61;        memory[64391] <=  8'h62;        memory[64392] <=  8'h74;        memory[64393] <=  8'h6e;        memory[64394] <=  8'h61;        memory[64395] <=  8'h72;        memory[64396] <=  8'h62;        memory[64397] <=  8'h78;        memory[64398] <=  8'h74;        memory[64399] <=  8'h61;        memory[64400] <=  8'h72;        memory[64401] <=  8'h62;        memory[64402] <=  8'h61;        memory[64403] <=  8'h72;        memory[64404] <=  8'h74;        memory[64405] <=  8'h74;        memory[64406] <=  8'h62;        memory[64407] <=  8'h61;        memory[64408] <=  8'h72;        memory[64409] <=  8'h74;        memory[64410] <=  8'h78;        memory[64411] <=  8'h61;        memory[64412] <=  8'h74;        memory[64413] <=  8'h6b;        memory[64414] <=  8'h73;        memory[64415] <=  8'h68;        memory[64416] <=  8'h63;        memory[64417] <=  8'h66;        memory[64418] <=  8'h69;        memory[64419] <=  8'h77;        memory[64420] <=  8'h68;        memory[64421] <=  8'h61;        memory[64422] <=  8'h74;        memory[64423] <=  8'h61;        memory[64424] <=  8'h6e;        memory[64425] <=  8'h61;        memory[64426] <=  8'h62;        memory[64427] <=  8'h61;        memory[64428] <=  8'h63;        memory[64429] <=  8'h61;        memory[64430] <=  8'h74;        memory[64431] <=  8'h61;        memory[64432] <=  8'h62;        memory[64433] <=  8'h61;        memory[64434] <=  8'h72;        memory[64435] <=  8'h63;        memory[64436] <=  8'h61;        memory[64437] <=  8'h68;        memory[64438] <=  8'h64;        memory[64439] <=  8'h75;        memory[64440] <=  8'h63;        memory[64441] <=  8'h74;        memory[64442] <=  8'h61;        memory[64443] <=  8'h64;        memory[64444] <=  8'h61;        memory[64445] <=  8'h61;        memory[64446] <=  8'h63;        memory[64447] <=  8'h61;        memory[64448] <=  8'h72;        memory[64449] <=  8'h63;        memory[64450] <=  8'h74;        memory[64451] <=  8'h72;        memory[64452] <=  8'h63;        memory[64453] <=  8'h61;        memory[64454] <=  8'h74;        memory[64455] <=  8'h72;        memory[64456] <=  8'h63;        memory[64457] <=  8'h61;        memory[64458] <=  8'h74;        memory[64459] <=  8'h63;        memory[64460] <=  8'h62;        memory[64461] <=  8'h61;        memory[64462] <=  8'h74;        memory[64463] <=  8'h62;        memory[64464] <=  8'h72;        memory[64465] <=  8'h63;        memory[64466] <=  8'h61;        memory[64467] <=  8'h74;        memory[64468] <=  8'h72;        memory[64469] <=  8'h6e;        memory[64470] <=  8'h62;        memory[64471] <=  8'h61;        memory[64472] <=  8'h63;        memory[64473] <=  8'h61;        memory[64474] <=  8'h74;        memory[64475] <=  8'h79;        memory[64476] <=  8'h73;        memory[64477] <=  8'h6e;        memory[64478] <=  8'h63;        memory[64479] <=  8'h74;        memory[64480] <=  8'h61;        memory[64481] <=  8'h6e;        memory[64482] <=  8'h62;        memory[64483] <=  8'h61;        memory[64484] <=  8'h63;        memory[64485] <=  8'h72;        memory[64486] <=  8'h6e;        memory[64487] <=  8'h74;        memory[64488] <=  8'h61;        memory[64489] <=  8'h62;        memory[64490] <=  8'h74;        memory[64491] <=  8'h6e;        memory[64492] <=  8'h61;        memory[64493] <=  8'h72;        memory[64494] <=  8'h62;        memory[64495] <=  8'h78;        memory[64496] <=  8'h74;        memory[64497] <=  8'h61;        memory[64498] <=  8'h72;        memory[64499] <=  8'h62;        memory[64500] <=  8'h61;        memory[64501] <=  8'h72;        memory[64502] <=  8'h74;        memory[64503] <=  8'h74;        memory[64504] <=  8'h62;        memory[64505] <=  8'h61;        memory[64506] <=  8'h72;        memory[64507] <=  8'h74;        memory[64508] <=  8'h78;        memory[64509] <=  8'h61;        memory[64510] <=  8'h74;        memory[64511] <=  8'h6b;        memory[64512] <=  8'h73;        memory[64513] <=  8'h68;        memory[64514] <=  8'h63;        memory[64515] <=  8'h66;        memory[64516] <=  8'h69;        memory[64517] <=  8'h77;        memory[64518] <=  8'h68;        memory[64519] <=  8'h61;        memory[64520] <=  8'h74;        memory[64521] <=  8'h61;        memory[64522] <=  8'h6e;        memory[64523] <=  8'h61;        memory[64524] <=  8'h62;        memory[64525] <=  8'h61;        memory[64526] <=  8'h63;        memory[64527] <=  8'h61;        memory[64528] <=  8'h74;        memory[64529] <=  8'h61;        memory[64530] <=  8'h62;        memory[64531] <=  8'h61;        memory[64532] <=  8'h72;        memory[64533] <=  8'h63;        memory[64534] <=  8'h61;        memory[64535] <=  8'h68;        memory[64536] <=  8'h64;        memory[64537] <=  8'h75;        memory[64538] <=  8'h63;        memory[64539] <=  8'h74;        memory[64540] <=  8'h61;        memory[64541] <=  8'h64;        memory[64542] <=  8'h61;        memory[64543] <=  8'h61;        memory[64544] <=  8'h63;        memory[64545] <=  8'h61;        memory[64546] <=  8'h72;        memory[64547] <=  8'h63;        memory[64548] <=  8'h74;        memory[64549] <=  8'h72;        memory[64550] <=  8'h63;        memory[64551] <=  8'h61;        memory[64552] <=  8'h74;        memory[64553] <=  8'h72;        memory[64554] <=  8'h63;        memory[64555] <=  8'h61;        memory[64556] <=  8'h74;        memory[64557] <=  8'h63;        memory[64558] <=  8'h62;        memory[64559] <=  8'h61;        memory[64560] <=  8'h74;        memory[64561] <=  8'h62;        memory[64562] <=  8'h72;        memory[64563] <=  8'h63;        memory[64564] <=  8'h61;        memory[64565] <=  8'h74;        memory[64566] <=  8'h72;        memory[64567] <=  8'h6e;        memory[64568] <=  8'h62;        memory[64569] <=  8'h61;        memory[64570] <=  8'h63;        memory[64571] <=  8'h61;        memory[64572] <=  8'h74;        memory[64573] <=  8'h79;        memory[64574] <=  8'h73;        memory[64575] <=  8'h6e;        memory[64576] <=  8'h63;        memory[64577] <=  8'h74;        memory[64578] <=  8'h61;        memory[64579] <=  8'h6e;        memory[64580] <=  8'h62;        memory[64581] <=  8'h61;        memory[64582] <=  8'h63;        memory[64583] <=  8'h72;        memory[64584] <=  8'h6e;        memory[64585] <=  8'h74;        memory[64586] <=  8'h61;        memory[64587] <=  8'h62;        memory[64588] <=  8'h74;        memory[64589] <=  8'h6e;        memory[64590] <=  8'h61;        memory[64591] <=  8'h72;        memory[64592] <=  8'h62;        memory[64593] <=  8'h78;        memory[64594] <=  8'h74;        memory[64595] <=  8'h61;        memory[64596] <=  8'h72;        memory[64597] <=  8'h5d;        memory[64598] <=  8'h5d;        memory[64599] <=  8'h65;        memory[64600] <=  8'h66;        memory[64601] <=  8'h77;        memory[64602] <=  8'h65;        memory[64603] <=  8'h5d;        memory[64604] <=  8'h65;        memory[64605] <=  8'h67;        memory[64606] <=  8'h73;        memory[64607] <=  8'h67;        memory[64608] <=  8'h66;        memory[64609] <=  8'h62;        memory[64610] <=  8'h61;        memory[64611] <=  8'h72;        memory[64612] <=  8'h74;        memory[64613] <=  8'h74;        memory[64614] <=  8'h62;        memory[64615] <=  8'h61;        memory[64616] <=  8'h72;        memory[64617] <=  8'h74;        memory[64618] <=  8'h78;        memory[64619] <=  8'h61;        memory[64620] <=  8'h74;        memory[64621] <=  8'h6b;        memory[64622] <=  8'h73;        memory[64623] <=  8'h68;        memory[64624] <=  8'h63;        memory[64625] <=  8'h66;        memory[64626] <=  8'h69;        memory[64627] <=  8'h77;        memory[64628] <=  8'h68;        memory[64629] <=  8'h61;        memory[64630] <=  8'h74;        memory[64631] <=  8'h61;        memory[64632] <=  8'h6e;        memory[64633] <=  8'h61;        memory[64634] <=  8'h62;        memory[64635] <=  8'h61;        memory[64636] <=  8'h63;        memory[64637] <=  8'h61;        memory[64638] <=  8'h74;        memory[64639] <=  8'h61;        memory[64640] <=  8'h62;        memory[64641] <=  8'h61;        memory[64642] <=  8'h72;        memory[64643] <=  8'h63;        memory[64644] <=  8'h61;        memory[64645] <=  8'h68;        memory[64646] <=  8'h64;        memory[64647] <=  8'h75;        memory[64648] <=  8'h63;        memory[64649] <=  8'h74;        memory[64650] <=  8'h61;        memory[64651] <=  8'h64;        memory[64652] <=  8'h61;        memory[64653] <=  8'h61;        memory[64654] <=  8'h63;        memory[64655] <=  8'h61;        memory[64656] <=  8'h72;        memory[64657] <=  8'h63;        memory[64658] <=  8'h74;        memory[64659] <=  8'h72;        memory[64660] <=  8'h63;        memory[64661] <=  8'h61;        memory[64662] <=  8'h74;        memory[64663] <=  8'h72;        memory[64664] <=  8'h63;        memory[64665] <=  8'h61;        memory[64666] <=  8'h74;        memory[64667] <=  8'h63;        memory[64668] <=  8'h62;        memory[64669] <=  8'h61;        memory[64670] <=  8'h74;        memory[64671] <=  8'h62;        memory[64672] <=  8'h72;        memory[64673] <=  8'h63;        memory[64674] <=  8'h61;        memory[64675] <=  8'h74;        memory[64676] <=  8'h72;        memory[64677] <=  8'h6e;        memory[64678] <=  8'h62;        memory[64679] <=  8'h61;        memory[64680] <=  8'h63;        memory[64681] <=  8'h61;        memory[64682] <=  8'h74;        memory[64683] <=  8'h79;        memory[64684] <=  8'h73;        memory[64685] <=  8'h6e;        memory[64686] <=  8'h63;        memory[64687] <=  8'h74;        memory[64688] <=  8'h61;        memory[64689] <=  8'h6e;        memory[64690] <=  8'h62;        memory[64691] <=  8'h61;        memory[64692] <=  8'h63;        memory[64693] <=  8'h72;        memory[64694] <=  8'h6e;        memory[64695] <=  8'h74;        memory[64696] <=  8'h61;        memory[64697] <=  8'h62;        memory[64698] <=  8'h74;        memory[64699] <=  8'h6e;        memory[64700] <=  8'h61;        memory[64701] <=  8'h72;        memory[64702] <=  8'h62;        memory[64703] <=  8'h78;        memory[64704] <=  8'h74;        memory[64705] <=  8'h61;        memory[64706] <=  8'h72;        memory[64707] <=  8'h62;        memory[64708] <=  8'h61;        memory[64709] <=  8'h72;        memory[64710] <=  8'h74;        memory[64711] <=  8'h74;        memory[64712] <=  8'h62;        memory[64713] <=  8'h61;        memory[64714] <=  8'h72;        memory[64715] <=  8'h74;        memory[64716] <=  8'h78;        memory[64717] <=  8'h61;        memory[64718] <=  8'h74;        memory[64719] <=  8'h6b;        memory[64720] <=  8'h73;        memory[64721] <=  8'h68;        memory[64722] <=  8'h63;        memory[64723] <=  8'h66;        memory[64724] <=  8'h69;        memory[64725] <=  8'h77;        memory[64726] <=  8'h68;        memory[64727] <=  8'h61;        memory[64728] <=  8'h74;        memory[64729] <=  8'h61;        memory[64730] <=  8'h6e;        memory[64731] <=  8'h61;        memory[64732] <=  8'h62;        memory[64733] <=  8'h61;        memory[64734] <=  8'h63;        memory[64735] <=  8'h61;        memory[64736] <=  8'h74;        memory[64737] <=  8'h61;        memory[64738] <=  8'h62;        memory[64739] <=  8'h61;        memory[64740] <=  8'h72;        memory[64741] <=  8'h63;        memory[64742] <=  8'h61;        memory[64743] <=  8'h68;        memory[64744] <=  8'h64;        memory[64745] <=  8'h75;        memory[64746] <=  8'h63;        memory[64747] <=  8'h74;        memory[64748] <=  8'h61;        memory[64749] <=  8'h64;        memory[64750] <=  8'h61;        memory[64751] <=  8'h61;        memory[64752] <=  8'h63;        memory[64753] <=  8'h61;        memory[64754] <=  8'h72;        memory[64755] <=  8'h63;        memory[64756] <=  8'h74;        memory[64757] <=  8'h72;        memory[64758] <=  8'h63;        memory[64759] <=  8'h61;        memory[64760] <=  8'h74;        memory[64761] <=  8'h72;        memory[64762] <=  8'h63;        memory[64763] <=  8'h61;        memory[64764] <=  8'h74;        memory[64765] <=  8'h63;        memory[64766] <=  8'h62;        memory[64767] <=  8'h61;        memory[64768] <=  8'h74;        memory[64769] <=  8'h62;        memory[64770] <=  8'h72;        memory[64771] <=  8'h63;        memory[64772] <=  8'h61;        memory[64773] <=  8'h74;        memory[64774] <=  8'h72;        memory[64775] <=  8'h6e;        memory[64776] <=  8'h62;        memory[64777] <=  8'h61;        memory[64778] <=  8'h63;        memory[64779] <=  8'h61;        memory[64780] <=  8'h74;        memory[64781] <=  8'h79;        memory[64782] <=  8'h73;        memory[64783] <=  8'h6e;        memory[64784] <=  8'h63;        memory[64785] <=  8'h74;        memory[64786] <=  8'h61;        memory[64787] <=  8'h6e;        memory[64788] <=  8'h62;        memory[64789] <=  8'h61;        memory[64790] <=  8'h63;        memory[64791] <=  8'h72;        memory[64792] <=  8'h6e;        memory[64793] <=  8'h74;        memory[64794] <=  8'h61;        memory[64795] <=  8'h62;        memory[64796] <=  8'h74;        memory[64797] <=  8'h6e;        memory[64798] <=  8'h61;        memory[64799] <=  8'h72;        memory[64800] <=  8'h62;        memory[64801] <=  8'h78;        memory[64802] <=  8'h74;        memory[64803] <=  8'h61;        memory[64804] <=  8'h72;        memory[64805] <=  8'h64;        memory[64806] <=  8'h66;        memory[64807] <=  8'h73;        memory[64808] <=  8'h67;        memory[64809] <=  8'h76;        memory[64810] <=  8'h68;        memory[64811] <=  8'h62;        memory[64812] <=  8'h6b;        memory[64813] <=  8'h6a;        memory[64814] <=  8'h6e;        memory[64815] <=  8'h6d;        memory[64816] <=  8'h62;        memory[64817] <=  8'h76;        memory[64818] <=  8'h78;        memory[64819] <=  8'h63;        memory[64820] <=  8'h73;        memory[64821] <=  8'h66;        memory[64822] <=  8'h72;        memory[64823] <=  8'h74;        memory[64824] <=  8'h79;        memory[64825] <=  8'h75;        memory[64826] <=  8'h6a;        memory[64827] <=  8'h6e;        memory[64828] <=  8'h62;        memory[64829] <=  8'h76;        memory[64830] <=  8'h63;        memory[64831] <=  8'h64;        memory[64832] <=  8'h74;        memory[64833] <=  8'h79;        memory[64834] <=  8'h75;        memory[64835] <=  8'h69;        memory[64836] <=  8'h6b;        memory[64837] <=  8'h6d;        memory[64838] <=  8'h6e;        memory[64839] <=  8'h62;        memory[64840] <=  8'h76;        memory[64841] <=  8'h63;        memory[64842] <=  8'h78;        memory[64843] <=  8'h73;        memory[64844] <=  8'h64;        memory[64845] <=  8'h72;        memory[64846] <=  8'h74;        memory[64847] <=  8'h79;        memory[64848] <=  8'h75;        memory[64849] <=  8'h69;        memory[64850] <=  8'h6b;        memory[64851] <=  8'h6d;        memory[64852] <=  8'h6e;        memory[64853] <=  8'h62;        memory[64854] <=  8'h76;        memory[64855] <=  8'h63;        memory[64856] <=  8'h73;        memory[64857] <=  8'h77;        memory[64858] <=  8'h33;        memory[64859] <=  8'h34;        memory[64860] <=  8'h35;        memory[64861] <=  8'h36;        memory[64862] <=  8'h37;        memory[64863] <=  8'h38;        memory[64864] <=  8'h69;        memory[64865] <=  8'h6b;        memory[64866] <=  8'h6d;        memory[64867] <=  8'h6e;        memory[64868] <=  8'h62;        memory[64869] <=  8'h76;        memory[64870] <=  8'h63;        memory[64871] <=  8'h64;        memory[64872] <=  8'h65;        memory[64873] <=  8'h72;        memory[64874] <=  8'h36;        memory[64875] <=  8'h37;        memory[64876] <=  8'h38;        memory[64877] <=  8'h69;        memory[64878] <=  8'h6f;        memory[64879] <=  8'h6b;        memory[64880] <=  8'h6a;        memory[64881] <=  8'h6e;        memory[64882] <=  8'h62;        memory[64883] <=  8'h76;        memory[64884] <=  8'h63;        memory[64885] <=  8'h64;        memory[64886] <=  8'h72;        memory[64887] <=  8'h74;        memory[64888] <=  8'h79;        memory[64889] <=  8'h75;        memory[64890] <=  8'h73;        memory[64891] <=  8'h6a;        memory[64892] <=  8'h63;        memory[64893] <=  8'h6e;        memory[64894] <=  8'h62;        memory[64895] <=  8'h64;        memory[64896] <=  8'h66;        memory[64897] <=  8'h73;        memory[64898] <=  8'h74;        memory[64899] <=  8'h79;        memory[64900] <=  8'h75;        memory[64901] <=  8'h61;        memory[64902] <=  8'h69;        memory[64903] <=  8'h6b;        memory[64904] <=  8'h78;        memory[64905] <=  8'h6d;        memory[64906] <=  8'h6e;        memory[64907] <=  8'h73;        memory[64908] <=  8'h6a;        memory[64909] <=  8'h6f;        memory[64910] <=  8'h64;        memory[64911] <=  8'h6c;        memory[64912] <=  8'h63;        memory[64913] <=  8'h78;        memory[64914] <=  8'h62;        memory[64915] <=  8'h61;        memory[64916] <=  8'h72;        memory[64917] <=  8'h74;        memory[64918] <=  8'h78;        memory[64919] <=  8'h61;        memory[64920] <=  8'h74;        memory[64921] <=  8'h6b;        memory[64922] <=  8'h73;        memory[64923] <=  8'h68;        memory[64924] <=  8'h63;        memory[64925] <=  8'h66;        memory[64926] <=  8'h69;        memory[64927] <=  8'h77;        memory[64928] <=  8'h68;        memory[64929] <=  8'h61;        memory[64930] <=  8'h74;        memory[64931] <=  8'h61;        memory[64932] <=  8'h6e;        memory[64933] <=  8'h61;        memory[64934] <=  8'h62;        memory[64935] <=  8'h61;        memory[64936] <=  8'h63;        memory[64937] <=  8'h61;        memory[64938] <=  8'h74;        memory[64939] <=  8'h61;        memory[64940] <=  8'h62;        memory[64941] <=  8'h61;        memory[64942] <=  8'h72;        memory[64943] <=  8'h63;        memory[64944] <=  8'h61;        memory[64945] <=  8'h68;        memory[64946] <=  8'h64;        memory[64947] <=  8'h75;        memory[64948] <=  8'h63;        memory[64949] <=  8'h74;        memory[64950] <=  8'h61;        memory[64951] <=  8'h64;        memory[64952] <=  8'h61;        memory[64953] <=  8'h61;        memory[64954] <=  8'h63;        memory[64955] <=  8'h61;        memory[64956] <=  8'h72;        memory[64957] <=  8'h62;        memory[64958] <=  8'h61;        memory[64959] <=  8'h72;        memory[64960] <=  8'h74;        memory[64961] <=  8'h78;        memory[64962] <=  8'h61;        memory[64963] <=  8'h74;        memory[64964] <=  8'h6b;        memory[64965] <=  8'h73;        memory[64966] <=  8'h68;        memory[64967] <=  8'h63;        memory[64968] <=  8'h66;        memory[64969] <=  8'h69;        memory[64970] <=  8'h77;        memory[64971] <=  8'h68;        memory[64972] <=  8'h61;        memory[64973] <=  8'h74;        memory[64974] <=  8'h61;        memory[64975] <=  8'h6e;        memory[64976] <=  8'h61;        memory[64977] <=  8'h62;        memory[64978] <=  8'h61;        memory[64979] <=  8'h63;        memory[64980] <=  8'h61;        memory[64981] <=  8'h74;        memory[64982] <=  8'h61;        memory[64983] <=  8'h62;        memory[64984] <=  8'h61;        memory[64985] <=  8'h72;        memory[64986] <=  8'h63;        memory[64987] <=  8'h61;        memory[64988] <=  8'h68;        memory[64989] <=  8'h64;        memory[64990] <=  8'h75;        memory[64991] <=  8'h63;        memory[64992] <=  8'h74;        memory[64993] <=  8'h61;        memory[64994] <=  8'h64;        memory[64995] <=  8'h61;        memory[64996] <=  8'h61;        memory[64997] <=  8'h63;        memory[64998] <=  8'h61;        memory[64999] <=  8'h72;        memory[65000] <=  8'h62;        memory[65001] <=  8'h61;        memory[65002] <=  8'h72;        memory[65003] <=  8'h74;        memory[65004] <=  8'h78;        memory[65005] <=  8'h61;        memory[65006] <=  8'h74;        memory[65007] <=  8'h6b;        memory[65008] <=  8'h73;        memory[65009] <=  8'h68;        memory[65010] <=  8'h63;        memory[65011] <=  8'h66;        memory[65012] <=  8'h69;        memory[65013] <=  8'h77;        memory[65014] <=  8'h68;        memory[65015] <=  8'h61;        memory[65016] <=  8'h74;        memory[65017] <=  8'h61;        memory[65018] <=  8'h6e;        memory[65019] <=  8'h61;        memory[65020] <=  8'h62;        memory[65021] <=  8'h61;        memory[65022] <=  8'h63;        memory[65023] <=  8'h61;        memory[65024] <=  8'h74;        memory[65025] <=  8'h61;        memory[65026] <=  8'h62;        memory[65027] <=  8'h61;        memory[65028] <=  8'h72;        memory[65029] <=  8'h63;        memory[65030] <=  8'h61;        memory[65031] <=  8'h68;        memory[65032] <=  8'h64;        memory[65033] <=  8'h75;        memory[65034] <=  8'h63;        memory[65035] <=  8'h74;        memory[65036] <=  8'h61;        memory[65037] <=  8'h64;        memory[65038] <=  8'h61;        memory[65039] <=  8'h61;        memory[65040] <=  8'h63;        memory[65041] <=  8'h61;        memory[65042] <=  8'h72;        memory[65043] <=  8'h62;        memory[65044] <=  8'h61;        memory[65045] <=  8'h72;        memory[65046] <=  8'h74;        memory[65047] <=  8'h78;        memory[65048] <=  8'h61;        memory[65049] <=  8'h74;        memory[65050] <=  8'h6b;        memory[65051] <=  8'h73;        memory[65052] <=  8'h68;        memory[65053] <=  8'h63;        memory[65054] <=  8'h66;        memory[65055] <=  8'h69;        memory[65056] <=  8'h77;        memory[65057] <=  8'h68;        memory[65058] <=  8'h61;        memory[65059] <=  8'h74;        memory[65060] <=  8'h61;        memory[65061] <=  8'h6e;        memory[65062] <=  8'h61;        memory[65063] <=  8'h62;        memory[65064] <=  8'h61;        memory[65065] <=  8'h63;        memory[65066] <=  8'h61;        memory[65067] <=  8'h74;        memory[65068] <=  8'h61;        memory[65069] <=  8'h62;        memory[65070] <=  8'h61;        memory[65071] <=  8'h72;        memory[65072] <=  8'h63;        memory[65073] <=  8'h61;        memory[65074] <=  8'h68;        memory[65075] <=  8'h64;        memory[65076] <=  8'h75;        memory[65077] <=  8'h63;        memory[65078] <=  8'h74;        memory[65079] <=  8'h61;        memory[65080] <=  8'h64;        memory[65081] <=  8'h61;        memory[65082] <=  8'h61;        memory[65083] <=  8'h63;        memory[65084] <=  8'h61;        memory[65085] <=  8'h72;        memory[65086] <=  8'h62;        memory[65087] <=  8'h61;        memory[65088] <=  8'h72;        memory[65089] <=  8'h74;        memory[65090] <=  8'h78;        memory[65091] <=  8'h61;        memory[65092] <=  8'h74;        memory[65093] <=  8'h6b;        memory[65094] <=  8'h73;        memory[65095] <=  8'h68;        memory[65096] <=  8'h63;        memory[65097] <=  8'h66;        memory[65098] <=  8'h69;        memory[65099] <=  8'h77;        memory[65100] <=  8'h68;        memory[65101] <=  8'h61;        memory[65102] <=  8'h74;        memory[65103] <=  8'h61;        memory[65104] <=  8'h6e;        memory[65105] <=  8'h61;        memory[65106] <=  8'h62;        memory[65107] <=  8'h61;        memory[65108] <=  8'h63;        memory[65109] <=  8'h61;        memory[65110] <=  8'h74;        memory[65111] <=  8'h61;        memory[65112] <=  8'h62;        memory[65113] <=  8'h61;        memory[65114] <=  8'h72;        memory[65115] <=  8'h63;        memory[65116] <=  8'h61;        memory[65117] <=  8'h68;        memory[65118] <=  8'h64;        memory[65119] <=  8'h75;        memory[65120] <=  8'h63;        memory[65121] <=  8'h74;        memory[65122] <=  8'h61;        memory[65123] <=  8'h64;        memory[65124] <=  8'h61;        memory[65125] <=  8'h61;        memory[65126] <=  8'h63;        memory[65127] <=  8'h61;        memory[65128] <=  8'h72;        memory[65129] <=  8'h62;        memory[65130] <=  8'h61;        memory[65131] <=  8'h72;        memory[65132] <=  8'h74;        memory[65133] <=  8'h78;        memory[65134] <=  8'h61;        memory[65135] <=  8'h74;        memory[65136] <=  8'h6b;        memory[65137] <=  8'h73;        memory[65138] <=  8'h68;        memory[65139] <=  8'h63;        memory[65140] <=  8'h66;        memory[65141] <=  8'h69;        memory[65142] <=  8'h77;        memory[65143] <=  8'h68;        memory[65144] <=  8'h61;        memory[65145] <=  8'h74;        memory[65146] <=  8'h61;        memory[65147] <=  8'h6e;        memory[65148] <=  8'h61;        memory[65149] <=  8'h62;        memory[65150] <=  8'h61;        memory[65151] <=  8'h63;        memory[65152] <=  8'h61;        memory[65153] <=  8'h74;        memory[65154] <=  8'h61;        memory[65155] <=  8'h62;        memory[65156] <=  8'h61;        memory[65157] <=  8'h72;        memory[65158] <=  8'h63;        memory[65159] <=  8'h61;        memory[65160] <=  8'h68;        memory[65161] <=  8'h64;        memory[65162] <=  8'h75;        memory[65163] <=  8'h63;        memory[65164] <=  8'h74;        memory[65165] <=  8'h61;        memory[65166] <=  8'h64;        memory[65167] <=  8'h61;        memory[65168] <=  8'h61;        memory[65169] <=  8'h63;        memory[65170] <=  8'h61;        memory[65171] <=  8'h72;        memory[65172] <=  8'h62;        memory[65173] <=  8'h61;        memory[65174] <=  8'h72;        memory[65175] <=  8'h74;        memory[65176] <=  8'h78;        memory[65177] <=  8'h61;        memory[65178] <=  8'h74;        memory[65179] <=  8'h6b;        memory[65180] <=  8'h73;        memory[65181] <=  8'h68;        memory[65182] <=  8'h63;        memory[65183] <=  8'h66;        memory[65184] <=  8'h69;        memory[65185] <=  8'h77;        memory[65186] <=  8'h68;        memory[65187] <=  8'h61;        memory[65188] <=  8'h74;        memory[65189] <=  8'h61;        memory[65190] <=  8'h6e;        memory[65191] <=  8'h61;        memory[65192] <=  8'h62;        memory[65193] <=  8'h61;        memory[65194] <=  8'h63;        memory[65195] <=  8'h61;        memory[65196] <=  8'h74;        memory[65197] <=  8'h61;        memory[65198] <=  8'h62;        memory[65199] <=  8'h61;        memory[65200] <=  8'h72;        memory[65201] <=  8'h63;        memory[65202] <=  8'h61;        memory[65203] <=  8'h68;        memory[65204] <=  8'h64;        memory[65205] <=  8'h75;        memory[65206] <=  8'h63;        memory[65207] <=  8'h74;        memory[65208] <=  8'h61;        memory[65209] <=  8'h64;        memory[65210] <=  8'h61;        memory[65211] <=  8'h61;        memory[65212] <=  8'h63;        memory[65213] <=  8'h61;        memory[65214] <=  8'h72;        memory[65215] <=  8'h62;        memory[65216] <=  8'h61;        memory[65217] <=  8'h72;        memory[65218] <=  8'h74;        memory[65219] <=  8'h78;        memory[65220] <=  8'h61;        memory[65221] <=  8'h74;        memory[65222] <=  8'h6b;        memory[65223] <=  8'h73;        memory[65224] <=  8'h68;        memory[65225] <=  8'h63;        memory[65226] <=  8'h66;        memory[65227] <=  8'h69;        memory[65228] <=  8'h77;        memory[65229] <=  8'h68;        memory[65230] <=  8'h61;        memory[65231] <=  8'h74;        memory[65232] <=  8'h61;        memory[65233] <=  8'h6e;        memory[65234] <=  8'h61;        memory[65235] <=  8'h62;        memory[65236] <=  8'h61;        memory[65237] <=  8'h63;        memory[65238] <=  8'h61;        memory[65239] <=  8'h74;        memory[65240] <=  8'h61;        memory[65241] <=  8'h62;        memory[65242] <=  8'h61;        memory[65243] <=  8'h72;        memory[65244] <=  8'h63;        memory[65245] <=  8'h61;        memory[65246] <=  8'h68;        memory[65247] <=  8'h64;        memory[65248] <=  8'h75;        memory[65249] <=  8'h63;        memory[65250] <=  8'h74;        memory[65251] <=  8'h61;        memory[65252] <=  8'h64;        memory[65253] <=  8'h61;        memory[65254] <=  8'h61;        memory[65255] <=  8'h63;        memory[65256] <=  8'h61;        memory[65257] <=  8'h72;        memory[65258] <=  8'h62;        memory[65259] <=  8'h61;        memory[65260] <=  8'h72;        memory[65261] <=  8'h74;        memory[65262] <=  8'h78;        memory[65263] <=  8'h61;        memory[65264] <=  8'h74;        memory[65265] <=  8'h6b;        memory[65266] <=  8'h73;        memory[65267] <=  8'h68;        memory[65268] <=  8'h63;        memory[65269] <=  8'h66;        memory[65270] <=  8'h69;        memory[65271] <=  8'h77;        memory[65272] <=  8'h68;        memory[65273] <=  8'h61;        memory[65274] <=  8'h74;        memory[65275] <=  8'h61;        memory[65276] <=  8'h6e;        memory[65277] <=  8'h61;        memory[65278] <=  8'h62;        memory[65279] <=  8'h61;        memory[65280] <=  8'h63;        memory[65281] <=  8'h61;        memory[65282] <=  8'h74;        memory[65283] <=  8'h61;        memory[65284] <=  8'h62;        memory[65285] <=  8'h61;        memory[65286] <=  8'h72;        memory[65287] <=  8'h63;        memory[65288] <=  8'h61;        memory[65289] <=  8'h68;        memory[65290] <=  8'h64;        memory[65291] <=  8'h75;        memory[65292] <=  8'h63;        memory[65293] <=  8'h74;        memory[65294] <=  8'h61;        memory[65295] <=  8'h64;        memory[65296] <=  8'h61;        memory[65297] <=  8'h61;        memory[65298] <=  8'h63;        memory[65299] <=  8'h61;        memory[65300] <=  8'h72;        memory[65301] <=  8'h00;        memory[65302] <=  8'h00;        memory[65303] <=  8'h00;        memory[65304] <=  8'h00;        memory[65305] <=  8'h00;        memory[65306] <=  8'h00;        memory[65307] <=  8'h00;        memory[65308] <=  8'h00;        memory[65309] <=  8'h00;        memory[65310] <=  8'h00;        memory[65311] <=  8'h00;        memory[65312] <=  8'h00;        memory[65313] <=  8'h00;        memory[65314] <=  8'h00;        memory[65315] <=  8'h00;        memory[65316] <=  8'h00;        memory[65317] <=  8'h00;        memory[65318] <=  8'h00;        memory[65319] <=  8'h00;        memory[65320] <=  8'h00;        memory[65321] <=  8'h00;        memory[65322] <=  8'h00;        memory[65323] <=  8'h00;        memory[65324] <=  8'h00;        memory[65325] <=  8'h00;        memory[65326] <=  8'h00;        memory[65327] <=  8'h00;        memory[65328] <=  8'h00;        memory[65329] <=  8'h00;        memory[65330] <=  8'h00;        memory[65331] <=  8'h00;        memory[65332] <=  8'h00;        memory[65333] <=  8'h00;        memory[65334] <=  8'h00;        memory[65335] <=  8'h00;        memory[65336] <=  8'h00;        memory[65337] <=  8'h00;        memory[65338] <=  8'h00;        memory[65339] <=  8'h00;        memory[65340] <=  8'h00;        memory[65341] <=  8'h00;        memory[65342] <=  8'h00;        memory[65343] <=  8'h00;        memory[65344] <=  8'h00;        memory[65345] <=  8'h00;        memory[65346] <=  8'h00;        memory[65347] <=  8'h00;        memory[65348] <=  8'h00;        memory[65349] <=  8'h00;        memory[65350] <=  8'h00;        memory[65351] <=  8'h00;        memory[65352] <=  8'h00;        memory[65353] <=  8'h00;        memory[65354] <=  8'h00;        memory[65355] <=  8'h00;        memory[65356] <=  8'h00;        memory[65357] <=  8'h00;        memory[65358] <=  8'h00;        memory[65359] <=  8'h00;        memory[65360] <=  8'h00;        memory[65361] <=  8'h00;        memory[65362] <=  8'h00;        memory[65363] <=  8'h00;        memory[65364] <=  8'h00;        memory[65365] <=  8'h00;        memory[65366] <=  8'h00;        memory[65367] <=  8'h00;        memory[65368] <=  8'h00;        memory[65369] <=  8'h00;        memory[65370] <=  8'h00;        memory[65371] <=  8'h00;        memory[65372] <=  8'h00;        memory[65373] <=  8'h00;        memory[65374] <=  8'h00;        memory[65375] <=  8'h00;        memory[65376] <=  8'h00;        memory[65377] <=  8'h00;        memory[65378] <=  8'h00;        memory[65379] <=  8'h00;        memory[65380] <=  8'h00;        memory[65381] <=  8'h00;        memory[65382] <=  8'h00;        memory[65383] <=  8'h00;        memory[65384] <=  8'h00;        memory[65385] <=  8'h00;        memory[65386] <=  8'h00;        memory[65387] <=  8'h00;        memory[65388] <=  8'h00;        memory[65389] <=  8'h00;        memory[65390] <=  8'h00;        memory[65391] <=  8'h00;        memory[65392] <=  8'h00;        memory[65393] <=  8'h00;        memory[65394] <=  8'h00;        memory[65395] <=  8'h00;        memory[65396] <=  8'h00;        memory[65397] <=  8'h00;        memory[65398] <=  8'h00;        memory[65399] <=  8'h00;        memory[65400] <=  8'h00;        memory[65401] <=  8'h00;        memory[65402] <=  8'h00;        memory[65403] <=  8'h00;        memory[65404] <=  8'h00;        memory[65405] <=  8'h00;        memory[65406] <=  8'h00;        memory[65407] <=  8'h00;        memory[65408] <=  8'h00;        memory[65409] <=  8'h00;        memory[65410] <=  8'h00;        memory[65411] <=  8'h00;        memory[65412] <=  8'h00;        memory[65413] <=  8'h00;        memory[65414] <=  8'h00;        memory[65415] <=  8'h00;        memory[65416] <=  8'h00;        memory[65417] <=  8'h00;        memory[65418] <=  8'h00;        memory[65419] <=  8'h00;        memory[65420] <=  8'h00;        memory[65421] <=  8'h00;        memory[65422] <=  8'h00;        memory[65423] <=  8'h00;        memory[65424] <=  8'h00;        memory[65425] <=  8'h00;        memory[65426] <=  8'h00;        memory[65427] <=  8'h00;        memory[65428] <=  8'h00;        memory[65429] <=  8'h00;        memory[65430] <=  8'h00;        memory[65431] <=  8'h00;        memory[65432] <=  8'h00;        memory[65433] <=  8'h00;        memory[65434] <=  8'h00;        memory[65435] <=  8'h00;        memory[65436] <=  8'h00;        memory[65437] <=  8'h00;        memory[65438] <=  8'h00;        memory[65439] <=  8'h00;        memory[65440] <=  8'h00;        memory[65441] <=  8'h00;        memory[65442] <=  8'h00;        memory[65443] <=  8'h00;        memory[65444] <=  8'h00;        memory[65445] <=  8'h00;        memory[65446] <=  8'h00;        memory[65447] <=  8'h00;        memory[65448] <=  8'h00;        memory[65449] <=  8'h00;        memory[65450] <=  8'h00;        memory[65451] <=  8'h00;        memory[65452] <=  8'h00;        memory[65453] <=  8'h00;        memory[65454] <=  8'h00;        memory[65455] <=  8'h00;        memory[65456] <=  8'h00;        memory[65457] <=  8'h00;        memory[65458] <=  8'h00;        memory[65459] <=  8'h00;        memory[65460] <=  8'h00;        memory[65461] <=  8'h00;        memory[65462] <=  8'h00;        memory[65463] <=  8'h00;        memory[65464] <=  8'h00;        memory[65465] <=  8'h00;        memory[65466] <=  8'h00;        memory[65467] <=  8'h00;        memory[65468] <=  8'h00;        memory[65469] <=  8'h00;        memory[65470] <=  8'h00;        memory[65471] <=  8'h00;        memory[65472] <=  8'h00;        memory[65473] <=  8'h00;        memory[65474] <=  8'h00;        memory[65475] <=  8'h00;        memory[65476] <=  8'h00;        memory[65477] <=  8'h00;        memory[65478] <=  8'h00;        memory[65479] <=  8'h00;        memory[65480] <=  8'h00;        memory[65481] <=  8'h00;        memory[65482] <=  8'h00;        memory[65483] <=  8'h00;        memory[65484] <=  8'h00;        memory[65485] <=  8'h00;        memory[65486] <=  8'h00;        memory[65487] <=  8'h00;        memory[65488] <=  8'h00;        memory[65489] <=  8'h00;        memory[65490] <=  8'h00;        memory[65491] <=  8'h00;        memory[65492] <=  8'h00;        memory[65493] <=  8'h00;        memory[65494] <=  8'h00;        memory[65495] <=  8'h00;        memory[65496] <=  8'h00;        memory[65497] <=  8'h00;        memory[65498] <=  8'h00;        memory[65499] <=  8'h00;        memory[65500] <=  8'h00;        memory[65501] <=  8'h00;        memory[65502] <=  8'h00;        memory[65503] <=  8'h00;        memory[65504] <=  8'h00;        memory[65505] <=  8'h00;        memory[65506] <=  8'h00;        memory[65507] <=  8'h00;        memory[65508] <=  8'h00;        memory[65509] <=  8'h00;        memory[65510] <=  8'h00;        memory[65511] <=  8'h00;        memory[65512] <=  8'h00;        memory[65513] <=  8'h00;        memory[65514] <=  8'h00;        memory[65515] <=  8'h00;        memory[65516] <=  8'h00;        memory[65517] <=  8'h00;        memory[65518] <=  8'h00;        memory[65519] <=  8'h00;        memory[65520] <=  8'h00;        memory[65521] <=  8'h00;        memory[65522] <=  8'h00;        memory[65523] <=  8'h00;        memory[65524] <=  8'h00;        memory[65525] <=  8'h00;        memory[65526] <=  8'h00;        memory[65527] <=  8'h00;        memory[65528] <=  8'h00;        memory[65529] <=  8'h00;        memory[65530] <=  8'h00;        memory[65531] <=  8'h00;        memory[65532] <=  8'h00;        memory[65533] <=  8'h00;        memory[65534] <=  8'h00;        memory[65535] <=  8'h00;    
    end

    always @(posedge clk) begin
        if (enable) begin
            if (we) begin
                memory[addr] <= write_data; // Write operation when we and enable are high
                reg_last_written_data <= write_data;
                reg_last_written_addr <= addr;
            end
        read_data_buff2  <= memory[addr]; // Read operation when enable is high
            read_data_buff1  <= read_data_buff2; // Read operation when enable is high
            read_data <= read_data_buff1; // Read operation when enable is high

        end
    end
 
endmodule





module BRAM_empty_AUTO (
    input wire clk,           // Clock signal 
    input wire [15:0] addr,    // Address input (8 bits)
    input wire we,            // Write enable signal
    input wire [7:0] write_data, // Data input (8 bits)
    input wire enable,        // Enable signal for read and write operations
    output reg [7:0] read_data // Data output (9 bits)
);
  reg [7:0] memory [0:65535]; // 65536x8-bit Block RAM

    reg [7:0] read_data_buff1, read_data_buff2, reg_last_written_data, reg_last_written_addr;
    initial begin
reg_last_written_data <= 8'b0;
reg_last_written_addr <= 8'b0;
read_data_buff1 <= 8'h00;
read_data_buff2 <= 8'h00;
read_data <=   8'h00;


    memory[0] <=  8'h00;      memory[1] <=  8'h00;      memory[2] <=  8'h00;      memory[3] <=  8'h00;      memory[4] <=  8'h00;      memory[5] <=  8'h00;      memory[6] <=  8'h00;      memory[7] <=  8'h00;      memory[8] <=  8'h00;      memory[9] <=  8'h00;      memory[10] <=  8'h00;      memory[11] <=  8'h00;      memory[12] <=  8'h00;      memory[13] <=  8'h00;      memory[14] <=  8'h00;      memory[15] <=  8'h00;      memory[16] <=  8'h00;      memory[17] <=  8'h00;      memory[18] <=  8'h00;      memory[19] <=  8'h00;      memory[20] <=  8'h00;      memory[21] <=  8'h00;      memory[22] <=  8'h00;      memory[23] <=  8'h00;      memory[24] <=  8'h00;      memory[25] <=  8'h00;      memory[26] <=  8'h00;      memory[27] <=  8'h00;      memory[28] <=  8'h00;      memory[29] <=  8'h00;      memory[30] <=  8'h00;      memory[31] <=  8'h00;      memory[32] <=  8'h00;      memory[33] <=  8'h00;      memory[34] <=  8'h00;      memory[35] <=  8'h00;      memory[36] <=  8'h00;      memory[37] <=  8'h00;      memory[38] <=  8'h00;      memory[39] <=  8'h00;      memory[40] <=  8'h00;      memory[41] <=  8'h00;      memory[42] <=  8'h00;      memory[43] <=  8'h00;      memory[44] <=  8'h00;      memory[45] <=  8'h00;      memory[46] <=  8'h00;      memory[47] <=  8'h00;      memory[48] <=  8'h00;      memory[49] <=  8'h00;      memory[50] <=  8'h00;      memory[51] <=  8'h00;      memory[52] <=  8'h00;      memory[53] <=  8'h00;      memory[54] <=  8'h00;      memory[55] <=  8'h00;      memory[56] <=  8'h00;      memory[57] <=  8'h00;      memory[58] <=  8'h00;      memory[59] <=  8'h00;      memory[60] <=  8'h00;      memory[61] <=  8'h00;      memory[62] <=  8'h00;      memory[63] <=  8'h00;      memory[64] <=  8'h00;      memory[65] <=  8'h00;      memory[66] <=  8'h00;      memory[67] <=  8'h00;      memory[68] <=  8'h00;      memory[69] <=  8'h00;      memory[70] <=  8'h00;      memory[71] <=  8'h00;      memory[72] <=  8'h00;      memory[73] <=  8'h00;      memory[74] <=  8'h00;      memory[75] <=  8'h00;      memory[76] <=  8'h00;      memory[77] <=  8'h00;      memory[78] <=  8'h00;      memory[79] <=  8'h00;      memory[80] <=  8'h00;      memory[81] <=  8'h00;      memory[82] <=  8'h00;      memory[83] <=  8'h00;      memory[84] <=  8'h00;      memory[85] <=  8'h00;      memory[86] <=  8'h00;      memory[87] <=  8'h00;      memory[88] <=  8'h00;      memory[89] <=  8'h00;      memory[90] <=  8'h00;      memory[91] <=  8'h00;      memory[92] <=  8'h00;      memory[93] <=  8'h00;      memory[94] <=  8'h00;      memory[95] <=  8'h00;      memory[96] <=  8'h00;      memory[97] <=  8'h00;      memory[98] <=  8'h00;      memory[99] <=  8'h00;      memory[100] <=  8'h00;      memory[101] <=  8'h00;      memory[102] <=  8'h00;      memory[103] <=  8'h00;      memory[104] <=  8'h00;      memory[105] <=  8'h00;      memory[106] <=  8'h00;      memory[107] <=  8'h00;      memory[108] <=  8'h00;      memory[109] <=  8'h00;      memory[110] <=  8'h00;      memory[111] <=  8'h00;      memory[112] <=  8'h00;      memory[113] <=  8'h00;      memory[114] <=  8'h00;      memory[115] <=  8'h00;      memory[116] <=  8'h00;      memory[117] <=  8'h00;      memory[118] <=  8'h00;      memory[119] <=  8'h00;      memory[120] <=  8'h00;      memory[121] <=  8'h00;      memory[122] <=  8'h00;      memory[123] <=  8'h00;      memory[124] <=  8'h00;      memory[125] <=  8'h00;      memory[126] <=  8'h00;      memory[127] <=  8'h00;      memory[128] <=  8'h00;      memory[129] <=  8'h00;      memory[130] <=  8'h00;      memory[131] <=  8'h00;      memory[132] <=  8'h00;      memory[133] <=  8'h00;      memory[134] <=  8'h00;      memory[135] <=  8'h00;      memory[136] <=  8'h00;      memory[137] <=  8'h00;      memory[138] <=  8'h00;      memory[139] <=  8'h00;      memory[140] <=  8'h00;      memory[141] <=  8'h00;      memory[142] <=  8'h00;      memory[143] <=  8'h00;      memory[144] <=  8'h00;      memory[145] <=  8'h00;      memory[146] <=  8'h00;      memory[147] <=  8'h00;      memory[148] <=  8'h00;      memory[149] <=  8'h00;      memory[150] <=  8'h00;      memory[151] <=  8'h00;      memory[152] <=  8'h00;      memory[153] <=  8'h00;      memory[154] <=  8'h00;      memory[155] <=  8'h00;      memory[156] <=  8'h00;      memory[157] <=  8'h00;      memory[158] <=  8'h00;      memory[159] <=  8'h00;      memory[160] <=  8'h00;      memory[161] <=  8'h00;      memory[162] <=  8'h00;      memory[163] <=  8'h00;      memory[164] <=  8'h00;      memory[165] <=  8'h00;      memory[166] <=  8'h00;      memory[167] <=  8'h00;      memory[168] <=  8'h00;      memory[169] <=  8'h00;      memory[170] <=  8'h00;      memory[171] <=  8'h00;      memory[172] <=  8'h00;      memory[173] <=  8'h00;      memory[174] <=  8'h00;      memory[175] <=  8'h00;      memory[176] <=  8'h00;      memory[177] <=  8'h00;      memory[178] <=  8'h00;      memory[179] <=  8'h00;      memory[180] <=  8'h00;      memory[181] <=  8'h00;      memory[182] <=  8'h00;      memory[183] <=  8'h00;      memory[184] <=  8'h00;      memory[185] <=  8'h00;      memory[186] <=  8'h00;      memory[187] <=  8'h00;      memory[188] <=  8'h00;      memory[189] <=  8'h00;      memory[190] <=  8'h00;      memory[191] <=  8'h00;      memory[192] <=  8'h00;      memory[193] <=  8'h00;      memory[194] <=  8'h00;      memory[195] <=  8'h00;      memory[196] <=  8'h00;      memory[197] <=  8'h00;      memory[198] <=  8'h00;      memory[199] <=  8'h00;      memory[200] <=  8'h00;      memory[201] <=  8'h00;      memory[202] <=  8'h00;      memory[203] <=  8'h00;      memory[204] <=  8'h00;      memory[205] <=  8'h00;      memory[206] <=  8'h00;      memory[207] <=  8'h00;      memory[208] <=  8'h00;      memory[209] <=  8'h00;      memory[210] <=  8'h00;      memory[211] <=  8'h00;      memory[212] <=  8'h00;      memory[213] <=  8'h00;      memory[214] <=  8'h00;      memory[215] <=  8'h00;      memory[216] <=  8'h00;      memory[217] <=  8'h00;      memory[218] <=  8'h00;      memory[219] <=  8'h00;      memory[220] <=  8'h00;      memory[221] <=  8'h00;      memory[222] <=  8'h00;      memory[223] <=  8'h00;      memory[224] <=  8'h00;      memory[225] <=  8'h00;      memory[226] <=  8'h00;      memory[227] <=  8'h00;      memory[228] <=  8'h00;      memory[229] <=  8'h00;      memory[230] <=  8'h00;      memory[231] <=  8'h00;      memory[232] <=  8'h00;      memory[233] <=  8'h00;      memory[234] <=  8'h00;      memory[235] <=  8'h00;      memory[236] <=  8'h00;      memory[237] <=  8'h00;      memory[238] <=  8'h00;      memory[239] <=  8'h00;      memory[240] <=  8'h00;      memory[241] <=  8'h00;      memory[242] <=  8'h00;      memory[243] <=  8'h00;      memory[244] <=  8'h00;      memory[245] <=  8'h00;      memory[246] <=  8'h00;      memory[247] <=  8'h00;      memory[248] <=  8'h00;      memory[249] <=  8'h00;      memory[250] <=  8'h00;      memory[251] <=  8'h00;      memory[252] <=  8'h00;      memory[253] <=  8'h00;      memory[254] <=  8'h00;      memory[255] <=  8'h00;      memory[256] <=  8'h00;      memory[257] <=  8'h00;      memory[258] <=  8'h00;      memory[259] <=  8'h00;      memory[260] <=  8'h00;      memory[261] <=  8'h00;      memory[262] <=  8'h00;      memory[263] <=  8'h00;      memory[264] <=  8'h00;      memory[265] <=  8'h00;      memory[266] <=  8'h00;      memory[267] <=  8'h00;      memory[268] <=  8'h00;      memory[269] <=  8'h00;      memory[270] <=  8'h00;      memory[271] <=  8'h00;      memory[272] <=  8'h00;      memory[273] <=  8'h00;      memory[274] <=  8'h00;      memory[275] <=  8'h00;      memory[276] <=  8'h00;      memory[277] <=  8'h00;      memory[278] <=  8'h00;      memory[279] <=  8'h00;      memory[280] <=  8'h00;      memory[281] <=  8'h00;      memory[282] <=  8'h00;      memory[283] <=  8'h00;      memory[284] <=  8'h00;      memory[285] <=  8'h00;      memory[286] <=  8'h00;      memory[287] <=  8'h00;      memory[288] <=  8'h00;      memory[289] <=  8'h00;      memory[290] <=  8'h00;      memory[291] <=  8'h00;      memory[292] <=  8'h00;      memory[293] <=  8'h00;      memory[294] <=  8'h00;      memory[295] <=  8'h00;      memory[296] <=  8'h00;      memory[297] <=  8'h00;      memory[298] <=  8'h00;      memory[299] <=  8'h00;      memory[300] <=  8'h00;      memory[301] <=  8'h00;      memory[302] <=  8'h00;      memory[303] <=  8'h00;      memory[304] <=  8'h00;      memory[305] <=  8'h00;      memory[306] <=  8'h00;      memory[307] <=  8'h00;      memory[308] <=  8'h00;      memory[309] <=  8'h00;      memory[310] <=  8'h00;      memory[311] <=  8'h00;      memory[312] <=  8'h00;      memory[313] <=  8'h00;      memory[314] <=  8'h00;      memory[315] <=  8'h00;      memory[316] <=  8'h00;      memory[317] <=  8'h00;      memory[318] <=  8'h00;      memory[319] <=  8'h00;      memory[320] <=  8'h00;      memory[321] <=  8'h00;      memory[322] <=  8'h00;      memory[323] <=  8'h00;      memory[324] <=  8'h00;      memory[325] <=  8'h00;      memory[326] <=  8'h00;      memory[327] <=  8'h00;      memory[328] <=  8'h00;      memory[329] <=  8'h00;      memory[330] <=  8'h00;      memory[331] <=  8'h00;      memory[332] <=  8'h00;      memory[333] <=  8'h00;      memory[334] <=  8'h00;      memory[335] <=  8'h00;      memory[336] <=  8'h00;      memory[337] <=  8'h00;      memory[338] <=  8'h00;      memory[339] <=  8'h00;      memory[340] <=  8'h00;      memory[341] <=  8'h00;      memory[342] <=  8'h00;      memory[343] <=  8'h00;      memory[344] <=  8'h00;      memory[345] <=  8'h00;      memory[346] <=  8'h00;      memory[347] <=  8'h00;      memory[348] <=  8'h00;      memory[349] <=  8'h00;      memory[350] <=  8'h00;      memory[351] <=  8'h00;      memory[352] <=  8'h00;      memory[353] <=  8'h00;      memory[354] <=  8'h00;      memory[355] <=  8'h00;      memory[356] <=  8'h00;      memory[357] <=  8'h00;      memory[358] <=  8'h00;      memory[359] <=  8'h00;      memory[360] <=  8'h00;      memory[361] <=  8'h00;      memory[362] <=  8'h00;      memory[363] <=  8'h00;      memory[364] <=  8'h00;      memory[365] <=  8'h00;      memory[366] <=  8'h00;      memory[367] <=  8'h00;      memory[368] <=  8'h00;      memory[369] <=  8'h00;      memory[370] <=  8'h00;      memory[371] <=  8'h00;      memory[372] <=  8'h00;      memory[373] <=  8'h00;      memory[374] <=  8'h00;      memory[375] <=  8'h00;      memory[376] <=  8'h00;      memory[377] <=  8'h00;      memory[378] <=  8'h00;      memory[379] <=  8'h00;      memory[380] <=  8'h00;      memory[381] <=  8'h00;      memory[382] <=  8'h00;      memory[383] <=  8'h00;      memory[384] <=  8'h00;      memory[385] <=  8'h00;      memory[386] <=  8'h00;      memory[387] <=  8'h00;      memory[388] <=  8'h00;      memory[389] <=  8'h00;      memory[390] <=  8'h00;      memory[391] <=  8'h00;      memory[392] <=  8'h00;      memory[393] <=  8'h00;      memory[394] <=  8'h00;      memory[395] <=  8'h00;      memory[396] <=  8'h00;      memory[397] <=  8'h00;      memory[398] <=  8'h00;      memory[399] <=  8'h00;      memory[400] <=  8'h00;      memory[401] <=  8'h00;      memory[402] <=  8'h00;      memory[403] <=  8'h00;      memory[404] <=  8'h00;      memory[405] <=  8'h00;      memory[406] <=  8'h00;      memory[407] <=  8'h00;      memory[408] <=  8'h00;      memory[409] <=  8'h00;      memory[410] <=  8'h00;      memory[411] <=  8'h00;      memory[412] <=  8'h00;      memory[413] <=  8'h00;      memory[414] <=  8'h00;      memory[415] <=  8'h00;      memory[416] <=  8'h00;      memory[417] <=  8'h00;      memory[418] <=  8'h00;      memory[419] <=  8'h00;      memory[420] <=  8'h00;      memory[421] <=  8'h00;      memory[422] <=  8'h00;      memory[423] <=  8'h00;      memory[424] <=  8'h00;      memory[425] <=  8'h00;      memory[426] <=  8'h00;      memory[427] <=  8'h00;      memory[428] <=  8'h00;      memory[429] <=  8'h00;      memory[430] <=  8'h00;      memory[431] <=  8'h00;      memory[432] <=  8'h00;      memory[433] <=  8'h00;      memory[434] <=  8'h00;      memory[435] <=  8'h00;      memory[436] <=  8'h00;      memory[437] <=  8'h00;      memory[438] <=  8'h00;      memory[439] <=  8'h00;      memory[440] <=  8'h00;      memory[441] <=  8'h00;      memory[442] <=  8'h00;      memory[443] <=  8'h00;      memory[444] <=  8'h00;      memory[445] <=  8'h00;      memory[446] <=  8'h00;      memory[447] <=  8'h00;      memory[448] <=  8'h00;      memory[449] <=  8'h00;      memory[450] <=  8'h00;      memory[451] <=  8'h00;      memory[452] <=  8'h00;      memory[453] <=  8'h00;      memory[454] <=  8'h00;      memory[455] <=  8'h00;      memory[456] <=  8'h00;      memory[457] <=  8'h00;      memory[458] <=  8'h00;      memory[459] <=  8'h00;      memory[460] <=  8'h00;      memory[461] <=  8'h00;      memory[462] <=  8'h00;      memory[463] <=  8'h00;      memory[464] <=  8'h00;      memory[465] <=  8'h00;      memory[466] <=  8'h00;      memory[467] <=  8'h00;      memory[468] <=  8'h00;      memory[469] <=  8'h00;      memory[470] <=  8'h00;      memory[471] <=  8'h00;      memory[472] <=  8'h00;      memory[473] <=  8'h00;      memory[474] <=  8'h00;      memory[475] <=  8'h00;      memory[476] <=  8'h00;      memory[477] <=  8'h00;      memory[478] <=  8'h00;      memory[479] <=  8'h00;      memory[480] <=  8'h00;      memory[481] <=  8'h00;      memory[482] <=  8'h00;      memory[483] <=  8'h00;      memory[484] <=  8'h00;      memory[485] <=  8'h00;      memory[486] <=  8'h00;      memory[487] <=  8'h00;      memory[488] <=  8'h00;      memory[489] <=  8'h00;      memory[490] <=  8'h00;      memory[491] <=  8'h00;      memory[492] <=  8'h00;      memory[493] <=  8'h00;      memory[494] <=  8'h00;      memory[495] <=  8'h00;      memory[496] <=  8'h00;      memory[497] <=  8'h00;      memory[498] <=  8'h00;      memory[499] <=  8'h00;      memory[500] <=  8'h00;      memory[501] <=  8'h00;      memory[502] <=  8'h00;      memory[503] <=  8'h00;      memory[504] <=  8'h00;      memory[505] <=  8'h00;      memory[506] <=  8'h00;      memory[507] <=  8'h00;      memory[508] <=  8'h00;      memory[509] <=  8'h00;      memory[510] <=  8'h00;      memory[511] <=  8'h00;      memory[512] <=  8'h00;      memory[513] <=  8'h00;      memory[514] <=  8'h00;      memory[515] <=  8'h00;      memory[516] <=  8'h00;      memory[517] <=  8'h00;      memory[518] <=  8'h00;      memory[519] <=  8'h00;      memory[520] <=  8'h00;      memory[521] <=  8'h00;      memory[522] <=  8'h00;      memory[523] <=  8'h00;      memory[524] <=  8'h00;      memory[525] <=  8'h00;      memory[526] <=  8'h00;      memory[527] <=  8'h00;      memory[528] <=  8'h00;      memory[529] <=  8'h00;      memory[530] <=  8'h00;      memory[531] <=  8'h00;      memory[532] <=  8'h00;      memory[533] <=  8'h00;      memory[534] <=  8'h00;      memory[535] <=  8'h00;      memory[536] <=  8'h00;      memory[537] <=  8'h00;      memory[538] <=  8'h00;      memory[539] <=  8'h00;      memory[540] <=  8'h00;      memory[541] <=  8'h00;      memory[542] <=  8'h00;      memory[543] <=  8'h00;      memory[544] <=  8'h00;      memory[545] <=  8'h00;      memory[546] <=  8'h00;      memory[547] <=  8'h00;      memory[548] <=  8'h00;      memory[549] <=  8'h00;      memory[550] <=  8'h00;      memory[551] <=  8'h00;      memory[552] <=  8'h00;      memory[553] <=  8'h00;      memory[554] <=  8'h00;      memory[555] <=  8'h00;      memory[556] <=  8'h00;      memory[557] <=  8'h00;      memory[558] <=  8'h00;      memory[559] <=  8'h00;      memory[560] <=  8'h00;      memory[561] <=  8'h00;      memory[562] <=  8'h00;      memory[563] <=  8'h00;      memory[564] <=  8'h00;      memory[565] <=  8'h00;      memory[566] <=  8'h00;      memory[567] <=  8'h00;      memory[568] <=  8'h00;      memory[569] <=  8'h00;      memory[570] <=  8'h00;      memory[571] <=  8'h00;      memory[572] <=  8'h00;      memory[573] <=  8'h00;      memory[574] <=  8'h00;      memory[575] <=  8'h00;      memory[576] <=  8'h00;      memory[577] <=  8'h00;      memory[578] <=  8'h00;      memory[579] <=  8'h00;      memory[580] <=  8'h00;      memory[581] <=  8'h00;      memory[582] <=  8'h00;      memory[583] <=  8'h00;      memory[584] <=  8'h00;      memory[585] <=  8'h00;      memory[586] <=  8'h00;      memory[587] <=  8'h00;      memory[588] <=  8'h00;      memory[589] <=  8'h00;      memory[590] <=  8'h00;      memory[591] <=  8'h00;      memory[592] <=  8'h00;      memory[593] <=  8'h00;      memory[594] <=  8'h00;      memory[595] <=  8'h00;      memory[596] <=  8'h00;      memory[597] <=  8'h00;      memory[598] <=  8'h00;      memory[599] <=  8'h00;      memory[600] <=  8'h00;      memory[601] <=  8'h00;      memory[602] <=  8'h00;      memory[603] <=  8'h00;      memory[604] <=  8'h00;      memory[605] <=  8'h00;      memory[606] <=  8'h00;      memory[607] <=  8'h00;      memory[608] <=  8'h00;      memory[609] <=  8'h00;      memory[610] <=  8'h00;      memory[611] <=  8'h00;      memory[612] <=  8'h00;      memory[613] <=  8'h00;      memory[614] <=  8'h00;      memory[615] <=  8'h00;      memory[616] <=  8'h00;      memory[617] <=  8'h00;      memory[618] <=  8'h00;      memory[619] <=  8'h00;      memory[620] <=  8'h00;      memory[621] <=  8'h00;      memory[622] <=  8'h00;      memory[623] <=  8'h00;      memory[624] <=  8'h00;      memory[625] <=  8'h00;      memory[626] <=  8'h00;      memory[627] <=  8'h00;      memory[628] <=  8'h00;      memory[629] <=  8'h00;      memory[630] <=  8'h00;      memory[631] <=  8'h00;      memory[632] <=  8'h00;      memory[633] <=  8'h00;      memory[634] <=  8'h00;      memory[635] <=  8'h00;      memory[636] <=  8'h00;      memory[637] <=  8'h00;      memory[638] <=  8'h00;      memory[639] <=  8'h00;      memory[640] <=  8'h00;      memory[641] <=  8'h00;      memory[642] <=  8'h00;      memory[643] <=  8'h00;      memory[644] <=  8'h00;      memory[645] <=  8'h00;      memory[646] <=  8'h00;      memory[647] <=  8'h00;      memory[648] <=  8'h00;      memory[649] <=  8'h00;      memory[650] <=  8'h00;      memory[651] <=  8'h00;      memory[652] <=  8'h00;      memory[653] <=  8'h00;      memory[654] <=  8'h00;      memory[655] <=  8'h00;      memory[656] <=  8'h00;      memory[657] <=  8'h00;      memory[658] <=  8'h00;      memory[659] <=  8'h00;      memory[660] <=  8'h00;      memory[661] <=  8'h00;      memory[662] <=  8'h00;      memory[663] <=  8'h00;      memory[664] <=  8'h00;      memory[665] <=  8'h00;      memory[666] <=  8'h00;      memory[667] <=  8'h00;      memory[668] <=  8'h00;      memory[669] <=  8'h00;      memory[670] <=  8'h00;      memory[671] <=  8'h00;      memory[672] <=  8'h00;      memory[673] <=  8'h00;      memory[674] <=  8'h00;      memory[675] <=  8'h00;      memory[676] <=  8'h00;      memory[677] <=  8'h00;      memory[678] <=  8'h00;      memory[679] <=  8'h00;      memory[680] <=  8'h00;      memory[681] <=  8'h00;      memory[682] <=  8'h00;      memory[683] <=  8'h00;      memory[684] <=  8'h00;      memory[685] <=  8'h00;      memory[686] <=  8'h00;      memory[687] <=  8'h00;      memory[688] <=  8'h00;      memory[689] <=  8'h00;      memory[690] <=  8'h00;      memory[691] <=  8'h00;      memory[692] <=  8'h00;      memory[693] <=  8'h00;      memory[694] <=  8'h00;      memory[695] <=  8'h00;      memory[696] <=  8'h00;      memory[697] <=  8'h00;      memory[698] <=  8'h00;      memory[699] <=  8'h00;      memory[700] <=  8'h00;      memory[701] <=  8'h00;      memory[702] <=  8'h00;      memory[703] <=  8'h00;      memory[704] <=  8'h00;      memory[705] <=  8'h00;      memory[706] <=  8'h00;      memory[707] <=  8'h00;      memory[708] <=  8'h00;      memory[709] <=  8'h00;      memory[710] <=  8'h00;      memory[711] <=  8'h00;      memory[712] <=  8'h00;      memory[713] <=  8'h00;      memory[714] <=  8'h00;      memory[715] <=  8'h00;      memory[716] <=  8'h00;      memory[717] <=  8'h00;      memory[718] <=  8'h00;      memory[719] <=  8'h00;      memory[720] <=  8'h00;      memory[721] <=  8'h00;      memory[722] <=  8'h00;      memory[723] <=  8'h00;      memory[724] <=  8'h00;      memory[725] <=  8'h00;      memory[726] <=  8'h00;      memory[727] <=  8'h00;      memory[728] <=  8'h00;      memory[729] <=  8'h00;      memory[730] <=  8'h00;      memory[731] <=  8'h00;      memory[732] <=  8'h00;      memory[733] <=  8'h00;      memory[734] <=  8'h00;      memory[735] <=  8'h00;      memory[736] <=  8'h00;      memory[737] <=  8'h00;      memory[738] <=  8'h00;      memory[739] <=  8'h00;      memory[740] <=  8'h00;      memory[741] <=  8'h00;      memory[742] <=  8'h00;      memory[743] <=  8'h00;      memory[744] <=  8'h00;      memory[745] <=  8'h00;      memory[746] <=  8'h00;      memory[747] <=  8'h00;      memory[748] <=  8'h00;      memory[749] <=  8'h00;      memory[750] <=  8'h00;      memory[751] <=  8'h00;      memory[752] <=  8'h00;      memory[753] <=  8'h00;      memory[754] <=  8'h00;      memory[755] <=  8'h00;      memory[756] <=  8'h00;      memory[757] <=  8'h00;      memory[758] <=  8'h00;      memory[759] <=  8'h00;      memory[760] <=  8'h00;      memory[761] <=  8'h00;      memory[762] <=  8'h00;      memory[763] <=  8'h00;      memory[764] <=  8'h00;      memory[765] <=  8'h00;      memory[766] <=  8'h00;      memory[767] <=  8'h00;      memory[768] <=  8'h00;      memory[769] <=  8'h00;      memory[770] <=  8'h00;      memory[771] <=  8'h00;      memory[772] <=  8'h00;      memory[773] <=  8'h00;      memory[774] <=  8'h00;      memory[775] <=  8'h00;      memory[776] <=  8'h00;      memory[777] <=  8'h00;      memory[778] <=  8'h00;      memory[779] <=  8'h00;      memory[780] <=  8'h00;      memory[781] <=  8'h00;      memory[782] <=  8'h00;      memory[783] <=  8'h00;      memory[784] <=  8'h00;      memory[785] <=  8'h00;      memory[786] <=  8'h00;      memory[787] <=  8'h00;      memory[788] <=  8'h00;      memory[789] <=  8'h00;      memory[790] <=  8'h00;      memory[791] <=  8'h00;      memory[792] <=  8'h00;      memory[793] <=  8'h00;      memory[794] <=  8'h00;      memory[795] <=  8'h00;      memory[796] <=  8'h00;      memory[797] <=  8'h00;      memory[798] <=  8'h00;      memory[799] <=  8'h00;      memory[800] <=  8'h00;      memory[801] <=  8'h00;      memory[802] <=  8'h00;      memory[803] <=  8'h00;      memory[804] <=  8'h00;      memory[805] <=  8'h00;      memory[806] <=  8'h00;      memory[807] <=  8'h00;      memory[808] <=  8'h00;      memory[809] <=  8'h00;      memory[810] <=  8'h00;      memory[811] <=  8'h00;      memory[812] <=  8'h00;      memory[813] <=  8'h00;      memory[814] <=  8'h00;      memory[815] <=  8'h00;      memory[816] <=  8'h00;      memory[817] <=  8'h00;      memory[818] <=  8'h00;      memory[819] <=  8'h00;      memory[820] <=  8'h00;      memory[821] <=  8'h00;      memory[822] <=  8'h00;      memory[823] <=  8'h00;      memory[824] <=  8'h00;      memory[825] <=  8'h00;      memory[826] <=  8'h00;      memory[827] <=  8'h00;      memory[828] <=  8'h00;      memory[829] <=  8'h00;      memory[830] <=  8'h00;      memory[831] <=  8'h00;      memory[832] <=  8'h00;      memory[833] <=  8'h00;      memory[834] <=  8'h00;      memory[835] <=  8'h00;      memory[836] <=  8'h00;      memory[837] <=  8'h00;      memory[838] <=  8'h00;      memory[839] <=  8'h00;      memory[840] <=  8'h00;      memory[841] <=  8'h00;      memory[842] <=  8'h00;      memory[843] <=  8'h00;      memory[844] <=  8'h00;      memory[845] <=  8'h00;      memory[846] <=  8'h00;      memory[847] <=  8'h00;      memory[848] <=  8'h00;      memory[849] <=  8'h00;      memory[850] <=  8'h00;      memory[851] <=  8'h00;      memory[852] <=  8'h00;      memory[853] <=  8'h00;      memory[854] <=  8'h00;      memory[855] <=  8'h00;      memory[856] <=  8'h00;      memory[857] <=  8'h00;      memory[858] <=  8'h00;      memory[859] <=  8'h00;      memory[860] <=  8'h00;      memory[861] <=  8'h00;      memory[862] <=  8'h00;      memory[863] <=  8'h00;      memory[864] <=  8'h00;      memory[865] <=  8'h00;      memory[866] <=  8'h00;      memory[867] <=  8'h00;      memory[868] <=  8'h00;      memory[869] <=  8'h00;      memory[870] <=  8'h00;      memory[871] <=  8'h00;      memory[872] <=  8'h00;      memory[873] <=  8'h00;      memory[874] <=  8'h00;      memory[875] <=  8'h00;      memory[876] <=  8'h00;      memory[877] <=  8'h00;      memory[878] <=  8'h00;      memory[879] <=  8'h00;      memory[880] <=  8'h00;      memory[881] <=  8'h00;      memory[882] <=  8'h00;      memory[883] <=  8'h00;      memory[884] <=  8'h00;      memory[885] <=  8'h00;      memory[886] <=  8'h00;      memory[887] <=  8'h00;      memory[888] <=  8'h00;      memory[889] <=  8'h00;      memory[890] <=  8'h00;      memory[891] <=  8'h00;      memory[892] <=  8'h00;      memory[893] <=  8'h00;      memory[894] <=  8'h00;      memory[895] <=  8'h00;      memory[896] <=  8'h00;      memory[897] <=  8'h00;      memory[898] <=  8'h00;      memory[899] <=  8'h00;      memory[900] <=  8'h00;      memory[901] <=  8'h00;      memory[902] <=  8'h00;      memory[903] <=  8'h00;      memory[904] <=  8'h00;      memory[905] <=  8'h00;      memory[906] <=  8'h00;      memory[907] <=  8'h00;      memory[908] <=  8'h00;      memory[909] <=  8'h00;      memory[910] <=  8'h00;      memory[911] <=  8'h00;      memory[912] <=  8'h00;      memory[913] <=  8'h00;      memory[914] <=  8'h00;      memory[915] <=  8'h00;      memory[916] <=  8'h00;      memory[917] <=  8'h00;      memory[918] <=  8'h00;      memory[919] <=  8'h00;      memory[920] <=  8'h00;      memory[921] <=  8'h00;      memory[922] <=  8'h00;      memory[923] <=  8'h00;      memory[924] <=  8'h00;      memory[925] <=  8'h00;      memory[926] <=  8'h00;      memory[927] <=  8'h00;      memory[928] <=  8'h00;      memory[929] <=  8'h00;      memory[930] <=  8'h00;      memory[931] <=  8'h00;      memory[932] <=  8'h00;      memory[933] <=  8'h00;      memory[934] <=  8'h00;      memory[935] <=  8'h00;      memory[936] <=  8'h00;      memory[937] <=  8'h00;      memory[938] <=  8'h00;      memory[939] <=  8'h00;      memory[940] <=  8'h00;      memory[941] <=  8'h00;      memory[942] <=  8'h00;      memory[943] <=  8'h00;      memory[944] <=  8'h00;      memory[945] <=  8'h00;      memory[946] <=  8'h00;      memory[947] <=  8'h00;      memory[948] <=  8'h00;      memory[949] <=  8'h00;      memory[950] <=  8'h00;      memory[951] <=  8'h00;      memory[952] <=  8'h00;      memory[953] <=  8'h00;      memory[954] <=  8'h00;      memory[955] <=  8'h00;      memory[956] <=  8'h00;      memory[957] <=  8'h00;      memory[958] <=  8'h00;      memory[959] <=  8'h00;      memory[960] <=  8'h00;      memory[961] <=  8'h00;      memory[962] <=  8'h00;      memory[963] <=  8'h00;      memory[964] <=  8'h00;      memory[965] <=  8'h00;      memory[966] <=  8'h00;      memory[967] <=  8'h00;      memory[968] <=  8'h00;      memory[969] <=  8'h00;      memory[970] <=  8'h00;      memory[971] <=  8'h00;      memory[972] <=  8'h00;      memory[973] <=  8'h00;      memory[974] <=  8'h00;      memory[975] <=  8'h00;      memory[976] <=  8'h00;      memory[977] <=  8'h00;      memory[978] <=  8'h00;      memory[979] <=  8'h00;      memory[980] <=  8'h00;      memory[981] <=  8'h00;      memory[982] <=  8'h00;      memory[983] <=  8'h00;      memory[984] <=  8'h00;      memory[985] <=  8'h00;      memory[986] <=  8'h00;      memory[987] <=  8'h00;      memory[988] <=  8'h00;      memory[989] <=  8'h00;      memory[990] <=  8'h00;      memory[991] <=  8'h00;      memory[992] <=  8'h00;      memory[993] <=  8'h00;      memory[994] <=  8'h00;      memory[995] <=  8'h00;      memory[996] <=  8'h00;      memory[997] <=  8'h00;      memory[998] <=  8'h00;      memory[999] <=  8'h00;      memory[1000] <=  8'h00;      memory[1001] <=  8'h00;      memory[1002] <=  8'h00;      memory[1003] <=  8'h00;      memory[1004] <=  8'h00;      memory[1005] <=  8'h00;      memory[1006] <=  8'h00;      memory[1007] <=  8'h00;      memory[1008] <=  8'h00;      memory[1009] <=  8'h00;      memory[1010] <=  8'h00;      memory[1011] <=  8'h00;      memory[1012] <=  8'h00;      memory[1013] <=  8'h00;      memory[1014] <=  8'h00;      memory[1015] <=  8'h00;      memory[1016] <=  8'h00;      memory[1017] <=  8'h00;      memory[1018] <=  8'h00;      memory[1019] <=  8'h00;      memory[1020] <=  8'h00;      memory[1021] <=  8'h00;      memory[1022] <=  8'h00;      memory[1023] <=  8'h00;      memory[1024] <=  8'h00;      memory[1025] <=  8'h00;      memory[1026] <=  8'h00;      memory[1027] <=  8'h00;      memory[1028] <=  8'h00;      memory[1029] <=  8'h00;      memory[1030] <=  8'h00;      memory[1031] <=  8'h00;      memory[1032] <=  8'h00;      memory[1033] <=  8'h00;      memory[1034] <=  8'h00;      memory[1035] <=  8'h00;      memory[1036] <=  8'h00;      memory[1037] <=  8'h00;      memory[1038] <=  8'h00;      memory[1039] <=  8'h00;      memory[1040] <=  8'h00;      memory[1041] <=  8'h00;      memory[1042] <=  8'h00;      memory[1043] <=  8'h00;      memory[1044] <=  8'h00;      memory[1045] <=  8'h00;      memory[1046] <=  8'h00;      memory[1047] <=  8'h00;      memory[1048] <=  8'h00;      memory[1049] <=  8'h00;      memory[1050] <=  8'h00;      memory[1051] <=  8'h00;      memory[1052] <=  8'h00;      memory[1053] <=  8'h00;      memory[1054] <=  8'h00;      memory[1055] <=  8'h00;      memory[1056] <=  8'h00;      memory[1057] <=  8'h00;      memory[1058] <=  8'h00;      memory[1059] <=  8'h00;      memory[1060] <=  8'h00;      memory[1061] <=  8'h00;      memory[1062] <=  8'h00;      memory[1063] <=  8'h00;      memory[1064] <=  8'h00;      memory[1065] <=  8'h00;      memory[1066] <=  8'h00;      memory[1067] <=  8'h00;      memory[1068] <=  8'h00;      memory[1069] <=  8'h00;      memory[1070] <=  8'h00;      memory[1071] <=  8'h00;      memory[1072] <=  8'h00;      memory[1073] <=  8'h00;      memory[1074] <=  8'h00;      memory[1075] <=  8'h00;      memory[1076] <=  8'h00;      memory[1077] <=  8'h00;      memory[1078] <=  8'h00;      memory[1079] <=  8'h00;      memory[1080] <=  8'h00;      memory[1081] <=  8'h00;      memory[1082] <=  8'h00;      memory[1083] <=  8'h00;      memory[1084] <=  8'h00;      memory[1085] <=  8'h00;      memory[1086] <=  8'h00;      memory[1087] <=  8'h00;      memory[1088] <=  8'h00;      memory[1089] <=  8'h00;      memory[1090] <=  8'h00;      memory[1091] <=  8'h00;      memory[1092] <=  8'h00;      memory[1093] <=  8'h00;      memory[1094] <=  8'h00;      memory[1095] <=  8'h00;      memory[1096] <=  8'h00;      memory[1097] <=  8'h00;      memory[1098] <=  8'h00;      memory[1099] <=  8'h00;      memory[1100] <=  8'h00;      memory[1101] <=  8'h00;      memory[1102] <=  8'h00;      memory[1103] <=  8'h00;      memory[1104] <=  8'h00;      memory[1105] <=  8'h00;      memory[1106] <=  8'h00;      memory[1107] <=  8'h00;      memory[1108] <=  8'h00;      memory[1109] <=  8'h00;      memory[1110] <=  8'h00;      memory[1111] <=  8'h00;      memory[1112] <=  8'h00;      memory[1113] <=  8'h00;      memory[1114] <=  8'h00;      memory[1115] <=  8'h00;      memory[1116] <=  8'h00;      memory[1117] <=  8'h00;      memory[1118] <=  8'h00;      memory[1119] <=  8'h00;      memory[1120] <=  8'h00;      memory[1121] <=  8'h00;      memory[1122] <=  8'h00;      memory[1123] <=  8'h00;      memory[1124] <=  8'h00;      memory[1125] <=  8'h00;      memory[1126] <=  8'h00;      memory[1127] <=  8'h00;      memory[1128] <=  8'h00;      memory[1129] <=  8'h00;      memory[1130] <=  8'h00;      memory[1131] <=  8'h00;      memory[1132] <=  8'h00;      memory[1133] <=  8'h00;      memory[1134] <=  8'h00;      memory[1135] <=  8'h00;      memory[1136] <=  8'h00;      memory[1137] <=  8'h00;      memory[1138] <=  8'h00;      memory[1139] <=  8'h00;      memory[1140] <=  8'h00;      memory[1141] <=  8'h00;      memory[1142] <=  8'h00;      memory[1143] <=  8'h00;      memory[1144] <=  8'h00;      memory[1145] <=  8'h00;      memory[1146] <=  8'h00;      memory[1147] <=  8'h00;      memory[1148] <=  8'h00;      memory[1149] <=  8'h00;      memory[1150] <=  8'h00;      memory[1151] <=  8'h00;      memory[1152] <=  8'h00;      memory[1153] <=  8'h00;      memory[1154] <=  8'h00;      memory[1155] <=  8'h00;      memory[1156] <=  8'h00;      memory[1157] <=  8'h00;      memory[1158] <=  8'h00;      memory[1159] <=  8'h00;      memory[1160] <=  8'h00;      memory[1161] <=  8'h00;      memory[1162] <=  8'h00;      memory[1163] <=  8'h00;      memory[1164] <=  8'h00;      memory[1165] <=  8'h00;      memory[1166] <=  8'h00;      memory[1167] <=  8'h00;      memory[1168] <=  8'h00;      memory[1169] <=  8'h00;      memory[1170] <=  8'h00;      memory[1171] <=  8'h00;      memory[1172] <=  8'h00;      memory[1173] <=  8'h00;      memory[1174] <=  8'h00;      memory[1175] <=  8'h00;      memory[1176] <=  8'h00;      memory[1177] <=  8'h00;      memory[1178] <=  8'h00;      memory[1179] <=  8'h00;      memory[1180] <=  8'h00;      memory[1181] <=  8'h00;      memory[1182] <=  8'h00;      memory[1183] <=  8'h00;      memory[1184] <=  8'h00;      memory[1185] <=  8'h00;      memory[1186] <=  8'h00;      memory[1187] <=  8'h00;      memory[1188] <=  8'h00;      memory[1189] <=  8'h00;      memory[1190] <=  8'h00;      memory[1191] <=  8'h00;      memory[1192] <=  8'h00;      memory[1193] <=  8'h00;      memory[1194] <=  8'h00;      memory[1195] <=  8'h00;      memory[1196] <=  8'h00;      memory[1197] <=  8'h00;      memory[1198] <=  8'h00;      memory[1199] <=  8'h00;      memory[1200] <=  8'h00;      memory[1201] <=  8'h00;      memory[1202] <=  8'h00;      memory[1203] <=  8'h00;      memory[1204] <=  8'h00;      memory[1205] <=  8'h00;      memory[1206] <=  8'h00;      memory[1207] <=  8'h00;      memory[1208] <=  8'h00;      memory[1209] <=  8'h00;      memory[1210] <=  8'h00;      memory[1211] <=  8'h00;      memory[1212] <=  8'h00;      memory[1213] <=  8'h00;      memory[1214] <=  8'h00;      memory[1215] <=  8'h00;      memory[1216] <=  8'h00;      memory[1217] <=  8'h00;      memory[1218] <=  8'h00;      memory[1219] <=  8'h00;      memory[1220] <=  8'h00;      memory[1221] <=  8'h00;      memory[1222] <=  8'h00;      memory[1223] <=  8'h00;      memory[1224] <=  8'h00;      memory[1225] <=  8'h00;      memory[1226] <=  8'h00;      memory[1227] <=  8'h00;      memory[1228] <=  8'h00;      memory[1229] <=  8'h00;      memory[1230] <=  8'h00;      memory[1231] <=  8'h00;      memory[1232] <=  8'h00;      memory[1233] <=  8'h00;      memory[1234] <=  8'h00;      memory[1235] <=  8'h00;      memory[1236] <=  8'h00;      memory[1237] <=  8'h00;      memory[1238] <=  8'h00;      memory[1239] <=  8'h00;      memory[1240] <=  8'h00;      memory[1241] <=  8'h00;      memory[1242] <=  8'h00;      memory[1243] <=  8'h00;      memory[1244] <=  8'h00;      memory[1245] <=  8'h00;      memory[1246] <=  8'h00;      memory[1247] <=  8'h00;      memory[1248] <=  8'h00;      memory[1249] <=  8'h00;      memory[1250] <=  8'h00;      memory[1251] <=  8'h00;      memory[1252] <=  8'h00;      memory[1253] <=  8'h00;      memory[1254] <=  8'h00;      memory[1255] <=  8'h00;      memory[1256] <=  8'h00;      memory[1257] <=  8'h00;      memory[1258] <=  8'h00;      memory[1259] <=  8'h00;      memory[1260] <=  8'h00;      memory[1261] <=  8'h00;      memory[1262] <=  8'h00;      memory[1263] <=  8'h00;      memory[1264] <=  8'h00;      memory[1265] <=  8'h00;      memory[1266] <=  8'h00;      memory[1267] <=  8'h00;      memory[1268] <=  8'h00;      memory[1269] <=  8'h00;      memory[1270] <=  8'h00;      memory[1271] <=  8'h00;      memory[1272] <=  8'h00;      memory[1273] <=  8'h00;      memory[1274] <=  8'h00;      memory[1275] <=  8'h00;      memory[1276] <=  8'h00;      memory[1277] <=  8'h00;      memory[1278] <=  8'h00;      memory[1279] <=  8'h00;      memory[1280] <=  8'h00;      memory[1281] <=  8'h00;      memory[1282] <=  8'h00;      memory[1283] <=  8'h00;      memory[1284] <=  8'h00;      memory[1285] <=  8'h00;      memory[1286] <=  8'h00;      memory[1287] <=  8'h00;      memory[1288] <=  8'h00;      memory[1289] <=  8'h00;      memory[1290] <=  8'h00;      memory[1291] <=  8'h00;      memory[1292] <=  8'h00;      memory[1293] <=  8'h00;      memory[1294] <=  8'h00;      memory[1295] <=  8'h00;      memory[1296] <=  8'h00;      memory[1297] <=  8'h00;      memory[1298] <=  8'h00;      memory[1299] <=  8'h00;      memory[1300] <=  8'h00;      memory[1301] <=  8'h00;      memory[1302] <=  8'h00;      memory[1303] <=  8'h00;      memory[1304] <=  8'h00;      memory[1305] <=  8'h00;      memory[1306] <=  8'h00;      memory[1307] <=  8'h00;      memory[1308] <=  8'h00;      memory[1309] <=  8'h00;      memory[1310] <=  8'h00;      memory[1311] <=  8'h00;      memory[1312] <=  8'h00;      memory[1313] <=  8'h00;      memory[1314] <=  8'h00;      memory[1315] <=  8'h00;      memory[1316] <=  8'h00;      memory[1317] <=  8'h00;      memory[1318] <=  8'h00;      memory[1319] <=  8'h00;      memory[1320] <=  8'h00;      memory[1321] <=  8'h00;      memory[1322] <=  8'h00;      memory[1323] <=  8'h00;      memory[1324] <=  8'h00;      memory[1325] <=  8'h00;      memory[1326] <=  8'h00;      memory[1327] <=  8'h00;      memory[1328] <=  8'h00;      memory[1329] <=  8'h00;      memory[1330] <=  8'h00;      memory[1331] <=  8'h00;      memory[1332] <=  8'h00;      memory[1333] <=  8'h00;      memory[1334] <=  8'h00;      memory[1335] <=  8'h00;      memory[1336] <=  8'h00;      memory[1337] <=  8'h00;      memory[1338] <=  8'h00;      memory[1339] <=  8'h00;      memory[1340] <=  8'h00;      memory[1341] <=  8'h00;      memory[1342] <=  8'h00;      memory[1343] <=  8'h00;      memory[1344] <=  8'h00;      memory[1345] <=  8'h00;      memory[1346] <=  8'h00;      memory[1347] <=  8'h00;      memory[1348] <=  8'h00;      memory[1349] <=  8'h00;      memory[1350] <=  8'h00;      memory[1351] <=  8'h00;      memory[1352] <=  8'h00;      memory[1353] <=  8'h00;      memory[1354] <=  8'h00;      memory[1355] <=  8'h00;      memory[1356] <=  8'h00;      memory[1357] <=  8'h00;      memory[1358] <=  8'h00;      memory[1359] <=  8'h00;      memory[1360] <=  8'h00;      memory[1361] <=  8'h00;      memory[1362] <=  8'h00;      memory[1363] <=  8'h00;      memory[1364] <=  8'h00;      memory[1365] <=  8'h00;      memory[1366] <=  8'h00;      memory[1367] <=  8'h00;      memory[1368] <=  8'h00;      memory[1369] <=  8'h00;      memory[1370] <=  8'h00;      memory[1371] <=  8'h00;      memory[1372] <=  8'h00;      memory[1373] <=  8'h00;      memory[1374] <=  8'h00;      memory[1375] <=  8'h00;      memory[1376] <=  8'h00;      memory[1377] <=  8'h00;      memory[1378] <=  8'h00;      memory[1379] <=  8'h00;      memory[1380] <=  8'h00;      memory[1381] <=  8'h00;      memory[1382] <=  8'h00;      memory[1383] <=  8'h00;      memory[1384] <=  8'h00;      memory[1385] <=  8'h00;      memory[1386] <=  8'h00;      memory[1387] <=  8'h00;      memory[1388] <=  8'h00;      memory[1389] <=  8'h00;      memory[1390] <=  8'h00;      memory[1391] <=  8'h00;      memory[1392] <=  8'h00;      memory[1393] <=  8'h00;      memory[1394] <=  8'h00;      memory[1395] <=  8'h00;      memory[1396] <=  8'h00;      memory[1397] <=  8'h00;      memory[1398] <=  8'h00;      memory[1399] <=  8'h00;      memory[1400] <=  8'h00;      memory[1401] <=  8'h00;      memory[1402] <=  8'h00;      memory[1403] <=  8'h00;      memory[1404] <=  8'h00;      memory[1405] <=  8'h00;      memory[1406] <=  8'h00;      memory[1407] <=  8'h00;      memory[1408] <=  8'h00;      memory[1409] <=  8'h00;      memory[1410] <=  8'h00;      memory[1411] <=  8'h00;      memory[1412] <=  8'h00;      memory[1413] <=  8'h00;      memory[1414] <=  8'h00;      memory[1415] <=  8'h00;      memory[1416] <=  8'h00;      memory[1417] <=  8'h00;      memory[1418] <=  8'h00;      memory[1419] <=  8'h00;      memory[1420] <=  8'h00;      memory[1421] <=  8'h00;      memory[1422] <=  8'h00;      memory[1423] <=  8'h00;      memory[1424] <=  8'h00;      memory[1425] <=  8'h00;      memory[1426] <=  8'h00;      memory[1427] <=  8'h00;      memory[1428] <=  8'h00;      memory[1429] <=  8'h00;      memory[1430] <=  8'h00;      memory[1431] <=  8'h00;      memory[1432] <=  8'h00;      memory[1433] <=  8'h00;      memory[1434] <=  8'h00;      memory[1435] <=  8'h00;      memory[1436] <=  8'h00;      memory[1437] <=  8'h00;      memory[1438] <=  8'h00;      memory[1439] <=  8'h00;      memory[1440] <=  8'h00;      memory[1441] <=  8'h00;      memory[1442] <=  8'h00;      memory[1443] <=  8'h00;      memory[1444] <=  8'h00;      memory[1445] <=  8'h00;      memory[1446] <=  8'h00;      memory[1447] <=  8'h00;      memory[1448] <=  8'h00;      memory[1449] <=  8'h00;      memory[1450] <=  8'h00;      memory[1451] <=  8'h00;      memory[1452] <=  8'h00;      memory[1453] <=  8'h00;      memory[1454] <=  8'h00;      memory[1455] <=  8'h00;      memory[1456] <=  8'h00;      memory[1457] <=  8'h00;      memory[1458] <=  8'h00;      memory[1459] <=  8'h00;      memory[1460] <=  8'h00;      memory[1461] <=  8'h00;      memory[1462] <=  8'h00;      memory[1463] <=  8'h00;      memory[1464] <=  8'h00;      memory[1465] <=  8'h00;      memory[1466] <=  8'h00;      memory[1467] <=  8'h00;      memory[1468] <=  8'h00;      memory[1469] <=  8'h00;      memory[1470] <=  8'h00;      memory[1471] <=  8'h00;      memory[1472] <=  8'h00;      memory[1473] <=  8'h00;      memory[1474] <=  8'h00;      memory[1475] <=  8'h00;      memory[1476] <=  8'h00;      memory[1477] <=  8'h00;      memory[1478] <=  8'h00;      memory[1479] <=  8'h00;      memory[1480] <=  8'h00;      memory[1481] <=  8'h00;      memory[1482] <=  8'h00;      memory[1483] <=  8'h00;      memory[1484] <=  8'h00;      memory[1485] <=  8'h00;      memory[1486] <=  8'h00;      memory[1487] <=  8'h00;      memory[1488] <=  8'h00;      memory[1489] <=  8'h00;      memory[1490] <=  8'h00;      memory[1491] <=  8'h00;      memory[1492] <=  8'h00;      memory[1493] <=  8'h00;      memory[1494] <=  8'h00;      memory[1495] <=  8'h00;      memory[1496] <=  8'h00;      memory[1497] <=  8'h00;      memory[1498] <=  8'h00;      memory[1499] <=  8'h00;      memory[1500] <=  8'h00;      memory[1501] <=  8'h00;      memory[1502] <=  8'h00;      memory[1503] <=  8'h00;      memory[1504] <=  8'h00;      memory[1505] <=  8'h00;      memory[1506] <=  8'h00;      memory[1507] <=  8'h00;      memory[1508] <=  8'h00;      memory[1509] <=  8'h00;      memory[1510] <=  8'h00;      memory[1511] <=  8'h00;      memory[1512] <=  8'h00;      memory[1513] <=  8'h00;      memory[1514] <=  8'h00;      memory[1515] <=  8'h00;      memory[1516] <=  8'h00;      memory[1517] <=  8'h00;      memory[1518] <=  8'h00;      memory[1519] <=  8'h00;      memory[1520] <=  8'h00;      memory[1521] <=  8'h00;      memory[1522] <=  8'h00;      memory[1523] <=  8'h00;      memory[1524] <=  8'h00;      memory[1525] <=  8'h00;      memory[1526] <=  8'h00;      memory[1527] <=  8'h00;      memory[1528] <=  8'h00;      memory[1529] <=  8'h00;      memory[1530] <=  8'h00;      memory[1531] <=  8'h00;      memory[1532] <=  8'h00;      memory[1533] <=  8'h00;      memory[1534] <=  8'h00;      memory[1535] <=  8'h00;      memory[1536] <=  8'h00;      memory[1537] <=  8'h00;      memory[1538] <=  8'h00;      memory[1539] <=  8'h00;      memory[1540] <=  8'h00;      memory[1541] <=  8'h00;      memory[1542] <=  8'h00;      memory[1543] <=  8'h00;      memory[1544] <=  8'h00;      memory[1545] <=  8'h00;      memory[1546] <=  8'h00;      memory[1547] <=  8'h00;      memory[1548] <=  8'h00;      memory[1549] <=  8'h00;      memory[1550] <=  8'h00;      memory[1551] <=  8'h00;      memory[1552] <=  8'h00;      memory[1553] <=  8'h00;      memory[1554] <=  8'h00;      memory[1555] <=  8'h00;      memory[1556] <=  8'h00;      memory[1557] <=  8'h00;      memory[1558] <=  8'h00;      memory[1559] <=  8'h00;      memory[1560] <=  8'h00;      memory[1561] <=  8'h00;      memory[1562] <=  8'h00;      memory[1563] <=  8'h00;      memory[1564] <=  8'h00;      memory[1565] <=  8'h00;      memory[1566] <=  8'h00;      memory[1567] <=  8'h00;      memory[1568] <=  8'h00;      memory[1569] <=  8'h00;      memory[1570] <=  8'h00;      memory[1571] <=  8'h00;      memory[1572] <=  8'h00;      memory[1573] <=  8'h00;      memory[1574] <=  8'h00;      memory[1575] <=  8'h00;      memory[1576] <=  8'h00;      memory[1577] <=  8'h00;      memory[1578] <=  8'h00;      memory[1579] <=  8'h00;      memory[1580] <=  8'h00;      memory[1581] <=  8'h00;      memory[1582] <=  8'h00;      memory[1583] <=  8'h00;      memory[1584] <=  8'h00;      memory[1585] <=  8'h00;      memory[1586] <=  8'h00;      memory[1587] <=  8'h00;      memory[1588] <=  8'h00;      memory[1589] <=  8'h00;      memory[1590] <=  8'h00;      memory[1591] <=  8'h00;      memory[1592] <=  8'h00;      memory[1593] <=  8'h00;      memory[1594] <=  8'h00;      memory[1595] <=  8'h00;      memory[1596] <=  8'h00;      memory[1597] <=  8'h00;      memory[1598] <=  8'h00;      memory[1599] <=  8'h00;      memory[1600] <=  8'h00;      memory[1601] <=  8'h00;      memory[1602] <=  8'h00;      memory[1603] <=  8'h00;      memory[1604] <=  8'h00;      memory[1605] <=  8'h00;      memory[1606] <=  8'h00;      memory[1607] <=  8'h00;      memory[1608] <=  8'h00;      memory[1609] <=  8'h00;      memory[1610] <=  8'h00;      memory[1611] <=  8'h00;      memory[1612] <=  8'h00;      memory[1613] <=  8'h00;      memory[1614] <=  8'h00;      memory[1615] <=  8'h00;      memory[1616] <=  8'h00;      memory[1617] <=  8'h00;      memory[1618] <=  8'h00;      memory[1619] <=  8'h00;      memory[1620] <=  8'h00;      memory[1621] <=  8'h00;      memory[1622] <=  8'h00;      memory[1623] <=  8'h00;      memory[1624] <=  8'h00;      memory[1625] <=  8'h00;      memory[1626] <=  8'h00;      memory[1627] <=  8'h00;      memory[1628] <=  8'h00;      memory[1629] <=  8'h00;      memory[1630] <=  8'h00;      memory[1631] <=  8'h00;      memory[1632] <=  8'h00;      memory[1633] <=  8'h00;      memory[1634] <=  8'h00;      memory[1635] <=  8'h00;      memory[1636] <=  8'h00;      memory[1637] <=  8'h00;      memory[1638] <=  8'h00;      memory[1639] <=  8'h00;      memory[1640] <=  8'h00;      memory[1641] <=  8'h00;      memory[1642] <=  8'h00;      memory[1643] <=  8'h00;      memory[1644] <=  8'h00;      memory[1645] <=  8'h00;      memory[1646] <=  8'h00;      memory[1647] <=  8'h00;      memory[1648] <=  8'h00;      memory[1649] <=  8'h00;      memory[1650] <=  8'h00;      memory[1651] <=  8'h00;      memory[1652] <=  8'h00;      memory[1653] <=  8'h00;      memory[1654] <=  8'h00;      memory[1655] <=  8'h00;      memory[1656] <=  8'h00;      memory[1657] <=  8'h00;      memory[1658] <=  8'h00;      memory[1659] <=  8'h00;      memory[1660] <=  8'h00;      memory[1661] <=  8'h00;      memory[1662] <=  8'h00;      memory[1663] <=  8'h00;      memory[1664] <=  8'h00;      memory[1665] <=  8'h00;      memory[1666] <=  8'h00;      memory[1667] <=  8'h00;      memory[1668] <=  8'h00;      memory[1669] <=  8'h00;      memory[1670] <=  8'h00;      memory[1671] <=  8'h00;      memory[1672] <=  8'h00;      memory[1673] <=  8'h00;      memory[1674] <=  8'h00;      memory[1675] <=  8'h00;      memory[1676] <=  8'h00;      memory[1677] <=  8'h00;      memory[1678] <=  8'h00;      memory[1679] <=  8'h00;      memory[1680] <=  8'h00;      memory[1681] <=  8'h00;      memory[1682] <=  8'h00;      memory[1683] <=  8'h00;      memory[1684] <=  8'h00;      memory[1685] <=  8'h00;      memory[1686] <=  8'h00;      memory[1687] <=  8'h00;      memory[1688] <=  8'h00;      memory[1689] <=  8'h00;      memory[1690] <=  8'h00;      memory[1691] <=  8'h00;      memory[1692] <=  8'h00;      memory[1693] <=  8'h00;      memory[1694] <=  8'h00;      memory[1695] <=  8'h00;      memory[1696] <=  8'h00;      memory[1697] <=  8'h00;      memory[1698] <=  8'h00;      memory[1699] <=  8'h00;      memory[1700] <=  8'h00;      memory[1701] <=  8'h00;      memory[1702] <=  8'h00;      memory[1703] <=  8'h00;      memory[1704] <=  8'h00;      memory[1705] <=  8'h00;      memory[1706] <=  8'h00;      memory[1707] <=  8'h00;      memory[1708] <=  8'h00;      memory[1709] <=  8'h00;      memory[1710] <=  8'h00;      memory[1711] <=  8'h00;      memory[1712] <=  8'h00;      memory[1713] <=  8'h00;      memory[1714] <=  8'h00;      memory[1715] <=  8'h00;      memory[1716] <=  8'h00;      memory[1717] <=  8'h00;      memory[1718] <=  8'h00;      memory[1719] <=  8'h00;      memory[1720] <=  8'h00;      memory[1721] <=  8'h00;      memory[1722] <=  8'h00;      memory[1723] <=  8'h00;      memory[1724] <=  8'h00;      memory[1725] <=  8'h00;      memory[1726] <=  8'h00;      memory[1727] <=  8'h00;      memory[1728] <=  8'h00;      memory[1729] <=  8'h00;      memory[1730] <=  8'h00;      memory[1731] <=  8'h00;      memory[1732] <=  8'h00;      memory[1733] <=  8'h00;      memory[1734] <=  8'h00;      memory[1735] <=  8'h00;      memory[1736] <=  8'h00;      memory[1737] <=  8'h00;      memory[1738] <=  8'h00;      memory[1739] <=  8'h00;      memory[1740] <=  8'h00;      memory[1741] <=  8'h00;      memory[1742] <=  8'h00;      memory[1743] <=  8'h00;      memory[1744] <=  8'h00;      memory[1745] <=  8'h00;      memory[1746] <=  8'h00;      memory[1747] <=  8'h00;      memory[1748] <=  8'h00;      memory[1749] <=  8'h00;      memory[1750] <=  8'h00;      memory[1751] <=  8'h00;      memory[1752] <=  8'h00;      memory[1753] <=  8'h00;      memory[1754] <=  8'h00;      memory[1755] <=  8'h00;      memory[1756] <=  8'h00;      memory[1757] <=  8'h00;      memory[1758] <=  8'h00;      memory[1759] <=  8'h00;      memory[1760] <=  8'h00;      memory[1761] <=  8'h00;      memory[1762] <=  8'h00;      memory[1763] <=  8'h00;      memory[1764] <=  8'h00;      memory[1765] <=  8'h00;      memory[1766] <=  8'h00;      memory[1767] <=  8'h00;      memory[1768] <=  8'h00;      memory[1769] <=  8'h00;      memory[1770] <=  8'h00;      memory[1771] <=  8'h00;      memory[1772] <=  8'h00;      memory[1773] <=  8'h00;      memory[1774] <=  8'h00;      memory[1775] <=  8'h00;      memory[1776] <=  8'h00;      memory[1777] <=  8'h00;      memory[1778] <=  8'h00;      memory[1779] <=  8'h00;      memory[1780] <=  8'h00;      memory[1781] <=  8'h00;      memory[1782] <=  8'h00;      memory[1783] <=  8'h00;      memory[1784] <=  8'h00;      memory[1785] <=  8'h00;      memory[1786] <=  8'h00;      memory[1787] <=  8'h00;      memory[1788] <=  8'h00;      memory[1789] <=  8'h00;      memory[1790] <=  8'h00;      memory[1791] <=  8'h00;      memory[1792] <=  8'h00;      memory[1793] <=  8'h00;      memory[1794] <=  8'h00;      memory[1795] <=  8'h00;      memory[1796] <=  8'h00;      memory[1797] <=  8'h00;      memory[1798] <=  8'h00;      memory[1799] <=  8'h00;      memory[1800] <=  8'h00;      memory[1801] <=  8'h00;      memory[1802] <=  8'h00;      memory[1803] <=  8'h00;      memory[1804] <=  8'h00;      memory[1805] <=  8'h00;      memory[1806] <=  8'h00;      memory[1807] <=  8'h00;      memory[1808] <=  8'h00;      memory[1809] <=  8'h00;      memory[1810] <=  8'h00;      memory[1811] <=  8'h00;      memory[1812] <=  8'h00;      memory[1813] <=  8'h00;      memory[1814] <=  8'h00;      memory[1815] <=  8'h00;      memory[1816] <=  8'h00;      memory[1817] <=  8'h00;      memory[1818] <=  8'h00;      memory[1819] <=  8'h00;      memory[1820] <=  8'h00;      memory[1821] <=  8'h00;      memory[1822] <=  8'h00;      memory[1823] <=  8'h00;      memory[1824] <=  8'h00;      memory[1825] <=  8'h00;      memory[1826] <=  8'h00;      memory[1827] <=  8'h00;      memory[1828] <=  8'h00;      memory[1829] <=  8'h00;      memory[1830] <=  8'h00;      memory[1831] <=  8'h00;      memory[1832] <=  8'h00;      memory[1833] <=  8'h00;      memory[1834] <=  8'h00;      memory[1835] <=  8'h00;      memory[1836] <=  8'h00;      memory[1837] <=  8'h00;      memory[1838] <=  8'h00;      memory[1839] <=  8'h00;      memory[1840] <=  8'h00;      memory[1841] <=  8'h00;      memory[1842] <=  8'h00;      memory[1843] <=  8'h00;      memory[1844] <=  8'h00;      memory[1845] <=  8'h00;      memory[1846] <=  8'h00;      memory[1847] <=  8'h00;      memory[1848] <=  8'h00;      memory[1849] <=  8'h00;      memory[1850] <=  8'h00;      memory[1851] <=  8'h00;      memory[1852] <=  8'h00;      memory[1853] <=  8'h00;      memory[1854] <=  8'h00;      memory[1855] <=  8'h00;      memory[1856] <=  8'h00;      memory[1857] <=  8'h00;      memory[1858] <=  8'h00;      memory[1859] <=  8'h00;      memory[1860] <=  8'h00;      memory[1861] <=  8'h00;      memory[1862] <=  8'h00;      memory[1863] <=  8'h00;      memory[1864] <=  8'h00;      memory[1865] <=  8'h00;      memory[1866] <=  8'h00;      memory[1867] <=  8'h00;      memory[1868] <=  8'h00;      memory[1869] <=  8'h00;      memory[1870] <=  8'h00;      memory[1871] <=  8'h00;      memory[1872] <=  8'h00;      memory[1873] <=  8'h00;      memory[1874] <=  8'h00;      memory[1875] <=  8'h00;      memory[1876] <=  8'h00;      memory[1877] <=  8'h00;      memory[1878] <=  8'h00;      memory[1879] <=  8'h00;      memory[1880] <=  8'h00;      memory[1881] <=  8'h00;      memory[1882] <=  8'h00;      memory[1883] <=  8'h00;      memory[1884] <=  8'h00;      memory[1885] <=  8'h00;      memory[1886] <=  8'h00;      memory[1887] <=  8'h00;      memory[1888] <=  8'h00;      memory[1889] <=  8'h00;      memory[1890] <=  8'h00;      memory[1891] <=  8'h00;      memory[1892] <=  8'h00;      memory[1893] <=  8'h00;      memory[1894] <=  8'h00;      memory[1895] <=  8'h00;      memory[1896] <=  8'h00;      memory[1897] <=  8'h00;      memory[1898] <=  8'h00;      memory[1899] <=  8'h00;      memory[1900] <=  8'h00;      memory[1901] <=  8'h00;      memory[1902] <=  8'h00;      memory[1903] <=  8'h00;      memory[1904] <=  8'h00;      memory[1905] <=  8'h00;      memory[1906] <=  8'h00;      memory[1907] <=  8'h00;      memory[1908] <=  8'h00;      memory[1909] <=  8'h00;      memory[1910] <=  8'h00;      memory[1911] <=  8'h00;      memory[1912] <=  8'h00;      memory[1913] <=  8'h00;      memory[1914] <=  8'h00;      memory[1915] <=  8'h00;      memory[1916] <=  8'h00;      memory[1917] <=  8'h00;      memory[1918] <=  8'h00;      memory[1919] <=  8'h00;      memory[1920] <=  8'h00;      memory[1921] <=  8'h00;      memory[1922] <=  8'h00;      memory[1923] <=  8'h00;      memory[1924] <=  8'h00;      memory[1925] <=  8'h00;      memory[1926] <=  8'h00;      memory[1927] <=  8'h00;      memory[1928] <=  8'h00;      memory[1929] <=  8'h00;      memory[1930] <=  8'h00;      memory[1931] <=  8'h00;      memory[1932] <=  8'h00;      memory[1933] <=  8'h00;      memory[1934] <=  8'h00;      memory[1935] <=  8'h00;      memory[1936] <=  8'h00;      memory[1937] <=  8'h00;      memory[1938] <=  8'h00;      memory[1939] <=  8'h00;      memory[1940] <=  8'h00;      memory[1941] <=  8'h00;      memory[1942] <=  8'h00;      memory[1943] <=  8'h00;      memory[1944] <=  8'h00;      memory[1945] <=  8'h00;      memory[1946] <=  8'h00;      memory[1947] <=  8'h00;      memory[1948] <=  8'h00;      memory[1949] <=  8'h00;      memory[1950] <=  8'h00;      memory[1951] <=  8'h00;      memory[1952] <=  8'h00;      memory[1953] <=  8'h00;      memory[1954] <=  8'h00;      memory[1955] <=  8'h00;      memory[1956] <=  8'h00;      memory[1957] <=  8'h00;      memory[1958] <=  8'h00;      memory[1959] <=  8'h00;      memory[1960] <=  8'h00;      memory[1961] <=  8'h00;      memory[1962] <=  8'h00;      memory[1963] <=  8'h00;      memory[1964] <=  8'h00;      memory[1965] <=  8'h00;      memory[1966] <=  8'h00;      memory[1967] <=  8'h00;      memory[1968] <=  8'h00;      memory[1969] <=  8'h00;      memory[1970] <=  8'h00;      memory[1971] <=  8'h00;      memory[1972] <=  8'h00;      memory[1973] <=  8'h00;      memory[1974] <=  8'h00;      memory[1975] <=  8'h00;      memory[1976] <=  8'h00;      memory[1977] <=  8'h00;      memory[1978] <=  8'h00;      memory[1979] <=  8'h00;      memory[1980] <=  8'h00;      memory[1981] <=  8'h00;      memory[1982] <=  8'h00;      memory[1983] <=  8'h00;      memory[1984] <=  8'h00;      memory[1985] <=  8'h00;      memory[1986] <=  8'h00;      memory[1987] <=  8'h00;      memory[1988] <=  8'h00;      memory[1989] <=  8'h00;      memory[1990] <=  8'h00;      memory[1991] <=  8'h00;      memory[1992] <=  8'h00;      memory[1993] <=  8'h00;      memory[1994] <=  8'h00;      memory[1995] <=  8'h00;      memory[1996] <=  8'h00;      memory[1997] <=  8'h00;      memory[1998] <=  8'h00;      memory[1999] <=  8'h00;      memory[2000] <=  8'h00;      memory[2001] <=  8'h00;      memory[2002] <=  8'h00;      memory[2003] <=  8'h00;      memory[2004] <=  8'h00;      memory[2005] <=  8'h00;      memory[2006] <=  8'h00;      memory[2007] <=  8'h00;      memory[2008] <=  8'h00;      memory[2009] <=  8'h00;      memory[2010] <=  8'h00;      memory[2011] <=  8'h00;      memory[2012] <=  8'h00;      memory[2013] <=  8'h00;      memory[2014] <=  8'h00;      memory[2015] <=  8'h00;      memory[2016] <=  8'h00;      memory[2017] <=  8'h00;      memory[2018] <=  8'h00;      memory[2019] <=  8'h00;      memory[2020] <=  8'h00;      memory[2021] <=  8'h00;      memory[2022] <=  8'h00;      memory[2023] <=  8'h00;      memory[2024] <=  8'h00;      memory[2025] <=  8'h00;      memory[2026] <=  8'h00;      memory[2027] <=  8'h00;      memory[2028] <=  8'h00;      memory[2029] <=  8'h00;      memory[2030] <=  8'h00;      memory[2031] <=  8'h00;      memory[2032] <=  8'h00;      memory[2033] <=  8'h00;      memory[2034] <=  8'h00;      memory[2035] <=  8'h00;      memory[2036] <=  8'h00;      memory[2037] <=  8'h00;      memory[2038] <=  8'h00;      memory[2039] <=  8'h00;      memory[2040] <=  8'h00;      memory[2041] <=  8'h00;      memory[2042] <=  8'h00;      memory[2043] <=  8'h00;      memory[2044] <=  8'h00;      memory[2045] <=  8'h00;      memory[2046] <=  8'h00;      memory[2047] <=  8'h00;      memory[2048] <=  8'h00;      memory[2049] <=  8'h00;      memory[2050] <=  8'h00;      memory[2051] <=  8'h00;      memory[2052] <=  8'h00;      memory[2053] <=  8'h00;      memory[2054] <=  8'h00;      memory[2055] <=  8'h00;      memory[2056] <=  8'h00;      memory[2057] <=  8'h00;      memory[2058] <=  8'h00;      memory[2059] <=  8'h00;      memory[2060] <=  8'h00;      memory[2061] <=  8'h00;      memory[2062] <=  8'h00;      memory[2063] <=  8'h00;      memory[2064] <=  8'h00;      memory[2065] <=  8'h00;      memory[2066] <=  8'h00;      memory[2067] <=  8'h00;      memory[2068] <=  8'h00;      memory[2069] <=  8'h00;      memory[2070] <=  8'h00;      memory[2071] <=  8'h00;      memory[2072] <=  8'h00;      memory[2073] <=  8'h00;      memory[2074] <=  8'h00;      memory[2075] <=  8'h00;      memory[2076] <=  8'h00;      memory[2077] <=  8'h00;      memory[2078] <=  8'h00;      memory[2079] <=  8'h00;      memory[2080] <=  8'h00;      memory[2081] <=  8'h00;      memory[2082] <=  8'h00;      memory[2083] <=  8'h00;      memory[2084] <=  8'h00;      memory[2085] <=  8'h00;      memory[2086] <=  8'h00;      memory[2087] <=  8'h00;      memory[2088] <=  8'h00;      memory[2089] <=  8'h00;      memory[2090] <=  8'h00;      memory[2091] <=  8'h00;      memory[2092] <=  8'h00;      memory[2093] <=  8'h00;      memory[2094] <=  8'h00;      memory[2095] <=  8'h00;      memory[2096] <=  8'h00;      memory[2097] <=  8'h00;      memory[2098] <=  8'h00;      memory[2099] <=  8'h00;      memory[2100] <=  8'h00;      memory[2101] <=  8'h00;      memory[2102] <=  8'h00;      memory[2103] <=  8'h00;      memory[2104] <=  8'h00;      memory[2105] <=  8'h00;      memory[2106] <=  8'h00;      memory[2107] <=  8'h00;      memory[2108] <=  8'h00;      memory[2109] <=  8'h00;      memory[2110] <=  8'h00;      memory[2111] <=  8'h00;      memory[2112] <=  8'h00;      memory[2113] <=  8'h00;      memory[2114] <=  8'h00;      memory[2115] <=  8'h00;      memory[2116] <=  8'h00;      memory[2117] <=  8'h00;      memory[2118] <=  8'h00;      memory[2119] <=  8'h00;      memory[2120] <=  8'h00;      memory[2121] <=  8'h00;      memory[2122] <=  8'h00;      memory[2123] <=  8'h00;      memory[2124] <=  8'h00;      memory[2125] <=  8'h00;      memory[2126] <=  8'h00;      memory[2127] <=  8'h00;      memory[2128] <=  8'h00;      memory[2129] <=  8'h00;      memory[2130] <=  8'h00;      memory[2131] <=  8'h00;      memory[2132] <=  8'h00;      memory[2133] <=  8'h00;      memory[2134] <=  8'h00;      memory[2135] <=  8'h00;      memory[2136] <=  8'h00;      memory[2137] <=  8'h00;      memory[2138] <=  8'h00;      memory[2139] <=  8'h00;      memory[2140] <=  8'h00;      memory[2141] <=  8'h00;      memory[2142] <=  8'h00;      memory[2143] <=  8'h00;      memory[2144] <=  8'h00;      memory[2145] <=  8'h00;      memory[2146] <=  8'h00;      memory[2147] <=  8'h00;      memory[2148] <=  8'h00;      memory[2149] <=  8'h00;      memory[2150] <=  8'h00;      memory[2151] <=  8'h00;      memory[2152] <=  8'h00;      memory[2153] <=  8'h00;      memory[2154] <=  8'h00;      memory[2155] <=  8'h00;      memory[2156] <=  8'h00;      memory[2157] <=  8'h00;      memory[2158] <=  8'h00;      memory[2159] <=  8'h00;      memory[2160] <=  8'h00;      memory[2161] <=  8'h00;      memory[2162] <=  8'h00;      memory[2163] <=  8'h00;      memory[2164] <=  8'h00;      memory[2165] <=  8'h00;      memory[2166] <=  8'h00;      memory[2167] <=  8'h00;      memory[2168] <=  8'h00;      memory[2169] <=  8'h00;      memory[2170] <=  8'h00;      memory[2171] <=  8'h00;      memory[2172] <=  8'h00;      memory[2173] <=  8'h00;      memory[2174] <=  8'h00;      memory[2175] <=  8'h00;      memory[2176] <=  8'h00;      memory[2177] <=  8'h00;      memory[2178] <=  8'h00;      memory[2179] <=  8'h00;      memory[2180] <=  8'h00;      memory[2181] <=  8'h00;      memory[2182] <=  8'h00;      memory[2183] <=  8'h00;      memory[2184] <=  8'h00;      memory[2185] <=  8'h00;      memory[2186] <=  8'h00;      memory[2187] <=  8'h00;      memory[2188] <=  8'h00;      memory[2189] <=  8'h00;      memory[2190] <=  8'h00;      memory[2191] <=  8'h00;      memory[2192] <=  8'h00;      memory[2193] <=  8'h00;      memory[2194] <=  8'h00;      memory[2195] <=  8'h00;      memory[2196] <=  8'h00;      memory[2197] <=  8'h00;      memory[2198] <=  8'h00;      memory[2199] <=  8'h00;      memory[2200] <=  8'h00;      memory[2201] <=  8'h00;      memory[2202] <=  8'h00;      memory[2203] <=  8'h00;      memory[2204] <=  8'h00;      memory[2205] <=  8'h00;      memory[2206] <=  8'h00;      memory[2207] <=  8'h00;      memory[2208] <=  8'h00;      memory[2209] <=  8'h00;      memory[2210] <=  8'h00;      memory[2211] <=  8'h00;      memory[2212] <=  8'h00;      memory[2213] <=  8'h00;      memory[2214] <=  8'h00;      memory[2215] <=  8'h00;      memory[2216] <=  8'h00;      memory[2217] <=  8'h00;      memory[2218] <=  8'h00;      memory[2219] <=  8'h00;      memory[2220] <=  8'h00;      memory[2221] <=  8'h00;      memory[2222] <=  8'h00;      memory[2223] <=  8'h00;      memory[2224] <=  8'h00;      memory[2225] <=  8'h00;      memory[2226] <=  8'h00;      memory[2227] <=  8'h00;      memory[2228] <=  8'h00;      memory[2229] <=  8'h00;      memory[2230] <=  8'h00;      memory[2231] <=  8'h00;      memory[2232] <=  8'h00;      memory[2233] <=  8'h00;      memory[2234] <=  8'h00;      memory[2235] <=  8'h00;      memory[2236] <=  8'h00;      memory[2237] <=  8'h00;      memory[2238] <=  8'h00;      memory[2239] <=  8'h00;      memory[2240] <=  8'h00;      memory[2241] <=  8'h00;      memory[2242] <=  8'h00;      memory[2243] <=  8'h00;      memory[2244] <=  8'h00;      memory[2245] <=  8'h00;      memory[2246] <=  8'h00;      memory[2247] <=  8'h00;      memory[2248] <=  8'h00;      memory[2249] <=  8'h00;      memory[2250] <=  8'h00;      memory[2251] <=  8'h00;      memory[2252] <=  8'h00;      memory[2253] <=  8'h00;      memory[2254] <=  8'h00;      memory[2255] <=  8'h00;      memory[2256] <=  8'h00;      memory[2257] <=  8'h00;      memory[2258] <=  8'h00;      memory[2259] <=  8'h00;      memory[2260] <=  8'h00;      memory[2261] <=  8'h00;      memory[2262] <=  8'h00;      memory[2263] <=  8'h00;      memory[2264] <=  8'h00;      memory[2265] <=  8'h00;      memory[2266] <=  8'h00;      memory[2267] <=  8'h00;      memory[2268] <=  8'h00;      memory[2269] <=  8'h00;      memory[2270] <=  8'h00;      memory[2271] <=  8'h00;      memory[2272] <=  8'h00;      memory[2273] <=  8'h00;      memory[2274] <=  8'h00;      memory[2275] <=  8'h00;      memory[2276] <=  8'h00;      memory[2277] <=  8'h00;      memory[2278] <=  8'h00;      memory[2279] <=  8'h00;      memory[2280] <=  8'h00;      memory[2281] <=  8'h00;      memory[2282] <=  8'h00;      memory[2283] <=  8'h00;      memory[2284] <=  8'h00;      memory[2285] <=  8'h00;      memory[2286] <=  8'h00;      memory[2287] <=  8'h00;      memory[2288] <=  8'h00;      memory[2289] <=  8'h00;      memory[2290] <=  8'h00;      memory[2291] <=  8'h00;      memory[2292] <=  8'h00;      memory[2293] <=  8'h00;      memory[2294] <=  8'h00;      memory[2295] <=  8'h00;      memory[2296] <=  8'h00;      memory[2297] <=  8'h00;      memory[2298] <=  8'h00;      memory[2299] <=  8'h00;      memory[2300] <=  8'h00;      memory[2301] <=  8'h00;      memory[2302] <=  8'h00;      memory[2303] <=  8'h00;      memory[2304] <=  8'h00;      memory[2305] <=  8'h00;      memory[2306] <=  8'h00;      memory[2307] <=  8'h00;      memory[2308] <=  8'h00;      memory[2309] <=  8'h00;      memory[2310] <=  8'h00;      memory[2311] <=  8'h00;      memory[2312] <=  8'h00;      memory[2313] <=  8'h00;      memory[2314] <=  8'h00;      memory[2315] <=  8'h00;      memory[2316] <=  8'h00;      memory[2317] <=  8'h00;      memory[2318] <=  8'h00;      memory[2319] <=  8'h00;      memory[2320] <=  8'h00;      memory[2321] <=  8'h00;      memory[2322] <=  8'h00;      memory[2323] <=  8'h00;      memory[2324] <=  8'h00;      memory[2325] <=  8'h00;      memory[2326] <=  8'h00;      memory[2327] <=  8'h00;      memory[2328] <=  8'h00;      memory[2329] <=  8'h00;      memory[2330] <=  8'h00;      memory[2331] <=  8'h00;      memory[2332] <=  8'h00;      memory[2333] <=  8'h00;      memory[2334] <=  8'h00;      memory[2335] <=  8'h00;      memory[2336] <=  8'h00;      memory[2337] <=  8'h00;      memory[2338] <=  8'h00;      memory[2339] <=  8'h00;      memory[2340] <=  8'h00;      memory[2341] <=  8'h00;      memory[2342] <=  8'h00;      memory[2343] <=  8'h00;      memory[2344] <=  8'h00;      memory[2345] <=  8'h00;      memory[2346] <=  8'h00;      memory[2347] <=  8'h00;      memory[2348] <=  8'h00;      memory[2349] <=  8'h00;      memory[2350] <=  8'h00;      memory[2351] <=  8'h00;      memory[2352] <=  8'h00;      memory[2353] <=  8'h00;      memory[2354] <=  8'h00;      memory[2355] <=  8'h00;      memory[2356] <=  8'h00;      memory[2357] <=  8'h00;      memory[2358] <=  8'h00;      memory[2359] <=  8'h00;      memory[2360] <=  8'h00;      memory[2361] <=  8'h00;      memory[2362] <=  8'h00;      memory[2363] <=  8'h00;      memory[2364] <=  8'h00;      memory[2365] <=  8'h00;      memory[2366] <=  8'h00;      memory[2367] <=  8'h00;      memory[2368] <=  8'h00;      memory[2369] <=  8'h00;      memory[2370] <=  8'h00;      memory[2371] <=  8'h00;      memory[2372] <=  8'h00;      memory[2373] <=  8'h00;      memory[2374] <=  8'h00;      memory[2375] <=  8'h00;      memory[2376] <=  8'h00;      memory[2377] <=  8'h00;      memory[2378] <=  8'h00;      memory[2379] <=  8'h00;      memory[2380] <=  8'h00;      memory[2381] <=  8'h00;      memory[2382] <=  8'h00;      memory[2383] <=  8'h00;      memory[2384] <=  8'h00;      memory[2385] <=  8'h00;      memory[2386] <=  8'h00;      memory[2387] <=  8'h00;      memory[2388] <=  8'h00;      memory[2389] <=  8'h00;      memory[2390] <=  8'h00;      memory[2391] <=  8'h00;      memory[2392] <=  8'h00;      memory[2393] <=  8'h00;      memory[2394] <=  8'h00;      memory[2395] <=  8'h00;      memory[2396] <=  8'h00;      memory[2397] <=  8'h00;      memory[2398] <=  8'h00;      memory[2399] <=  8'h00;      memory[2400] <=  8'h00;      memory[2401] <=  8'h00;      memory[2402] <=  8'h00;      memory[2403] <=  8'h00;      memory[2404] <=  8'h00;      memory[2405] <=  8'h00;      memory[2406] <=  8'h00;      memory[2407] <=  8'h00;      memory[2408] <=  8'h00;      memory[2409] <=  8'h00;      memory[2410] <=  8'h00;      memory[2411] <=  8'h00;      memory[2412] <=  8'h00;      memory[2413] <=  8'h00;      memory[2414] <=  8'h00;      memory[2415] <=  8'h00;      memory[2416] <=  8'h00;      memory[2417] <=  8'h00;      memory[2418] <=  8'h00;      memory[2419] <=  8'h00;      memory[2420] <=  8'h00;      memory[2421] <=  8'h00;      memory[2422] <=  8'h00;      memory[2423] <=  8'h00;      memory[2424] <=  8'h00;      memory[2425] <=  8'h00;      memory[2426] <=  8'h00;      memory[2427] <=  8'h00;      memory[2428] <=  8'h00;      memory[2429] <=  8'h00;      memory[2430] <=  8'h00;      memory[2431] <=  8'h00;      memory[2432] <=  8'h00;      memory[2433] <=  8'h00;      memory[2434] <=  8'h00;      memory[2435] <=  8'h00;      memory[2436] <=  8'h00;      memory[2437] <=  8'h00;      memory[2438] <=  8'h00;      memory[2439] <=  8'h00;      memory[2440] <=  8'h00;      memory[2441] <=  8'h00;      memory[2442] <=  8'h00;      memory[2443] <=  8'h00;      memory[2444] <=  8'h00;      memory[2445] <=  8'h00;      memory[2446] <=  8'h00;      memory[2447] <=  8'h00;      memory[2448] <=  8'h00;      memory[2449] <=  8'h00;      memory[2450] <=  8'h00;      memory[2451] <=  8'h00;      memory[2452] <=  8'h00;      memory[2453] <=  8'h00;      memory[2454] <=  8'h00;      memory[2455] <=  8'h00;      memory[2456] <=  8'h00;      memory[2457] <=  8'h00;      memory[2458] <=  8'h00;      memory[2459] <=  8'h00;      memory[2460] <=  8'h00;      memory[2461] <=  8'h00;      memory[2462] <=  8'h00;      memory[2463] <=  8'h00;      memory[2464] <=  8'h00;      memory[2465] <=  8'h00;      memory[2466] <=  8'h00;      memory[2467] <=  8'h00;      memory[2468] <=  8'h00;      memory[2469] <=  8'h00;      memory[2470] <=  8'h00;      memory[2471] <=  8'h00;      memory[2472] <=  8'h00;      memory[2473] <=  8'h00;      memory[2474] <=  8'h00;      memory[2475] <=  8'h00;      memory[2476] <=  8'h00;      memory[2477] <=  8'h00;      memory[2478] <=  8'h00;      memory[2479] <=  8'h00;      memory[2480] <=  8'h00;      memory[2481] <=  8'h00;      memory[2482] <=  8'h00;      memory[2483] <=  8'h00;      memory[2484] <=  8'h00;      memory[2485] <=  8'h00;      memory[2486] <=  8'h00;      memory[2487] <=  8'h00;      memory[2488] <=  8'h00;      memory[2489] <=  8'h00;      memory[2490] <=  8'h00;      memory[2491] <=  8'h00;      memory[2492] <=  8'h00;      memory[2493] <=  8'h00;      memory[2494] <=  8'h00;      memory[2495] <=  8'h00;      memory[2496] <=  8'h00;      memory[2497] <=  8'h00;      memory[2498] <=  8'h00;      memory[2499] <=  8'h00;      memory[2500] <=  8'h00;      memory[2501] <=  8'h00;      memory[2502] <=  8'h00;      memory[2503] <=  8'h00;      memory[2504] <=  8'h00;      memory[2505] <=  8'h00;      memory[2506] <=  8'h00;      memory[2507] <=  8'h00;      memory[2508] <=  8'h00;      memory[2509] <=  8'h00;      memory[2510] <=  8'h00;      memory[2511] <=  8'h00;      memory[2512] <=  8'h00;      memory[2513] <=  8'h00;      memory[2514] <=  8'h00;      memory[2515] <=  8'h00;      memory[2516] <=  8'h00;      memory[2517] <=  8'h00;      memory[2518] <=  8'h00;      memory[2519] <=  8'h00;      memory[2520] <=  8'h00;      memory[2521] <=  8'h00;      memory[2522] <=  8'h00;      memory[2523] <=  8'h00;      memory[2524] <=  8'h00;      memory[2525] <=  8'h00;      memory[2526] <=  8'h00;      memory[2527] <=  8'h00;      memory[2528] <=  8'h00;      memory[2529] <=  8'h00;      memory[2530] <=  8'h00;      memory[2531] <=  8'h00;      memory[2532] <=  8'h00;      memory[2533] <=  8'h00;      memory[2534] <=  8'h00;      memory[2535] <=  8'h00;      memory[2536] <=  8'h00;      memory[2537] <=  8'h00;      memory[2538] <=  8'h00;      memory[2539] <=  8'h00;      memory[2540] <=  8'h00;      memory[2541] <=  8'h00;      memory[2542] <=  8'h00;      memory[2543] <=  8'h00;      memory[2544] <=  8'h00;      memory[2545] <=  8'h00;      memory[2546] <=  8'h00;      memory[2547] <=  8'h00;      memory[2548] <=  8'h00;      memory[2549] <=  8'h00;      memory[2550] <=  8'h00;      memory[2551] <=  8'h00;      memory[2552] <=  8'h00;      memory[2553] <=  8'h00;      memory[2554] <=  8'h00;      memory[2555] <=  8'h00;      memory[2556] <=  8'h00;      memory[2557] <=  8'h00;      memory[2558] <=  8'h00;      memory[2559] <=  8'h00;      memory[2560] <=  8'h00;      memory[2561] <=  8'h00;      memory[2562] <=  8'h00;      memory[2563] <=  8'h00;      memory[2564] <=  8'h00;      memory[2565] <=  8'h00;      memory[2566] <=  8'h00;      memory[2567] <=  8'h00;      memory[2568] <=  8'h00;      memory[2569] <=  8'h00;      memory[2570] <=  8'h00;      memory[2571] <=  8'h00;      memory[2572] <=  8'h00;      memory[2573] <=  8'h00;      memory[2574] <=  8'h00;      memory[2575] <=  8'h00;      memory[2576] <=  8'h00;      memory[2577] <=  8'h00;      memory[2578] <=  8'h00;      memory[2579] <=  8'h00;      memory[2580] <=  8'h00;      memory[2581] <=  8'h00;      memory[2582] <=  8'h00;      memory[2583] <=  8'h00;      memory[2584] <=  8'h00;      memory[2585] <=  8'h00;      memory[2586] <=  8'h00;      memory[2587] <=  8'h00;      memory[2588] <=  8'h00;      memory[2589] <=  8'h00;      memory[2590] <=  8'h00;      memory[2591] <=  8'h00;      memory[2592] <=  8'h00;      memory[2593] <=  8'h00;      memory[2594] <=  8'h00;      memory[2595] <=  8'h00;      memory[2596] <=  8'h00;      memory[2597] <=  8'h00;      memory[2598] <=  8'h00;      memory[2599] <=  8'h00;      memory[2600] <=  8'h00;      memory[2601] <=  8'h00;      memory[2602] <=  8'h00;      memory[2603] <=  8'h00;      memory[2604] <=  8'h00;      memory[2605] <=  8'h00;      memory[2606] <=  8'h00;      memory[2607] <=  8'h00;      memory[2608] <=  8'h00;      memory[2609] <=  8'h00;      memory[2610] <=  8'h00;      memory[2611] <=  8'h00;      memory[2612] <=  8'h00;      memory[2613] <=  8'h00;      memory[2614] <=  8'h00;      memory[2615] <=  8'h00;      memory[2616] <=  8'h00;      memory[2617] <=  8'h00;      memory[2618] <=  8'h00;      memory[2619] <=  8'h00;      memory[2620] <=  8'h00;      memory[2621] <=  8'h00;      memory[2622] <=  8'h00;      memory[2623] <=  8'h00;      memory[2624] <=  8'h00;      memory[2625] <=  8'h00;      memory[2626] <=  8'h00;      memory[2627] <=  8'h00;      memory[2628] <=  8'h00;      memory[2629] <=  8'h00;      memory[2630] <=  8'h00;      memory[2631] <=  8'h00;      memory[2632] <=  8'h00;      memory[2633] <=  8'h00;      memory[2634] <=  8'h00;      memory[2635] <=  8'h00;      memory[2636] <=  8'h00;      memory[2637] <=  8'h00;      memory[2638] <=  8'h00;      memory[2639] <=  8'h00;      memory[2640] <=  8'h00;      memory[2641] <=  8'h00;      memory[2642] <=  8'h00;      memory[2643] <=  8'h00;      memory[2644] <=  8'h00;      memory[2645] <=  8'h00;      memory[2646] <=  8'h00;      memory[2647] <=  8'h00;      memory[2648] <=  8'h00;      memory[2649] <=  8'h00;      memory[2650] <=  8'h00;      memory[2651] <=  8'h00;      memory[2652] <=  8'h00;      memory[2653] <=  8'h00;      memory[2654] <=  8'h00;      memory[2655] <=  8'h00;      memory[2656] <=  8'h00;      memory[2657] <=  8'h00;      memory[2658] <=  8'h00;      memory[2659] <=  8'h00;      memory[2660] <=  8'h00;      memory[2661] <=  8'h00;      memory[2662] <=  8'h00;      memory[2663] <=  8'h00;      memory[2664] <=  8'h00;      memory[2665] <=  8'h00;      memory[2666] <=  8'h00;      memory[2667] <=  8'h00;      memory[2668] <=  8'h00;      memory[2669] <=  8'h00;      memory[2670] <=  8'h00;      memory[2671] <=  8'h00;      memory[2672] <=  8'h00;      memory[2673] <=  8'h00;      memory[2674] <=  8'h00;      memory[2675] <=  8'h00;      memory[2676] <=  8'h00;      memory[2677] <=  8'h00;      memory[2678] <=  8'h00;      memory[2679] <=  8'h00;      memory[2680] <=  8'h00;      memory[2681] <=  8'h00;      memory[2682] <=  8'h00;      memory[2683] <=  8'h00;      memory[2684] <=  8'h00;      memory[2685] <=  8'h00;      memory[2686] <=  8'h00;      memory[2687] <=  8'h00;      memory[2688] <=  8'h00;      memory[2689] <=  8'h00;      memory[2690] <=  8'h00;      memory[2691] <=  8'h00;      memory[2692] <=  8'h00;      memory[2693] <=  8'h00;      memory[2694] <=  8'h00;      memory[2695] <=  8'h00;      memory[2696] <=  8'h00;      memory[2697] <=  8'h00;      memory[2698] <=  8'h00;      memory[2699] <=  8'h00;      memory[2700] <=  8'h00;      memory[2701] <=  8'h00;      memory[2702] <=  8'h00;      memory[2703] <=  8'h00;      memory[2704] <=  8'h00;      memory[2705] <=  8'h00;      memory[2706] <=  8'h00;      memory[2707] <=  8'h00;      memory[2708] <=  8'h00;      memory[2709] <=  8'h00;      memory[2710] <=  8'h00;      memory[2711] <=  8'h00;      memory[2712] <=  8'h00;      memory[2713] <=  8'h00;      memory[2714] <=  8'h00;      memory[2715] <=  8'h00;      memory[2716] <=  8'h00;      memory[2717] <=  8'h00;      memory[2718] <=  8'h00;      memory[2719] <=  8'h00;      memory[2720] <=  8'h00;      memory[2721] <=  8'h00;      memory[2722] <=  8'h00;      memory[2723] <=  8'h00;      memory[2724] <=  8'h00;      memory[2725] <=  8'h00;      memory[2726] <=  8'h00;      memory[2727] <=  8'h00;      memory[2728] <=  8'h00;      memory[2729] <=  8'h00;      memory[2730] <=  8'h00;      memory[2731] <=  8'h00;      memory[2732] <=  8'h00;      memory[2733] <=  8'h00;      memory[2734] <=  8'h00;      memory[2735] <=  8'h00;      memory[2736] <=  8'h00;      memory[2737] <=  8'h00;      memory[2738] <=  8'h00;      memory[2739] <=  8'h00;      memory[2740] <=  8'h00;      memory[2741] <=  8'h00;      memory[2742] <=  8'h00;      memory[2743] <=  8'h00;      memory[2744] <=  8'h00;      memory[2745] <=  8'h00;      memory[2746] <=  8'h00;      memory[2747] <=  8'h00;      memory[2748] <=  8'h00;      memory[2749] <=  8'h00;      memory[2750] <=  8'h00;      memory[2751] <=  8'h00;      memory[2752] <=  8'h00;      memory[2753] <=  8'h00;      memory[2754] <=  8'h00;      memory[2755] <=  8'h00;      memory[2756] <=  8'h00;      memory[2757] <=  8'h00;      memory[2758] <=  8'h00;      memory[2759] <=  8'h00;      memory[2760] <=  8'h00;      memory[2761] <=  8'h00;      memory[2762] <=  8'h00;      memory[2763] <=  8'h00;      memory[2764] <=  8'h00;      memory[2765] <=  8'h00;      memory[2766] <=  8'h00;      memory[2767] <=  8'h00;      memory[2768] <=  8'h00;      memory[2769] <=  8'h00;      memory[2770] <=  8'h00;      memory[2771] <=  8'h00;      memory[2772] <=  8'h00;      memory[2773] <=  8'h00;      memory[2774] <=  8'h00;      memory[2775] <=  8'h00;      memory[2776] <=  8'h00;      memory[2777] <=  8'h00;      memory[2778] <=  8'h00;      memory[2779] <=  8'h00;      memory[2780] <=  8'h00;      memory[2781] <=  8'h00;      memory[2782] <=  8'h00;      memory[2783] <=  8'h00;      memory[2784] <=  8'h00;      memory[2785] <=  8'h00;      memory[2786] <=  8'h00;      memory[2787] <=  8'h00;      memory[2788] <=  8'h00;      memory[2789] <=  8'h00;      memory[2790] <=  8'h00;      memory[2791] <=  8'h00;      memory[2792] <=  8'h00;      memory[2793] <=  8'h00;      memory[2794] <=  8'h00;      memory[2795] <=  8'h00;      memory[2796] <=  8'h00;      memory[2797] <=  8'h00;      memory[2798] <=  8'h00;      memory[2799] <=  8'h00;      memory[2800] <=  8'h00;      memory[2801] <=  8'h00;      memory[2802] <=  8'h00;      memory[2803] <=  8'h00;      memory[2804] <=  8'h00;      memory[2805] <=  8'h00;      memory[2806] <=  8'h00;      memory[2807] <=  8'h00;      memory[2808] <=  8'h00;      memory[2809] <=  8'h00;      memory[2810] <=  8'h00;      memory[2811] <=  8'h00;      memory[2812] <=  8'h00;      memory[2813] <=  8'h00;      memory[2814] <=  8'h00;      memory[2815] <=  8'h00;      memory[2816] <=  8'h00;      memory[2817] <=  8'h00;      memory[2818] <=  8'h00;      memory[2819] <=  8'h00;      memory[2820] <=  8'h00;      memory[2821] <=  8'h00;      memory[2822] <=  8'h00;      memory[2823] <=  8'h00;      memory[2824] <=  8'h00;      memory[2825] <=  8'h00;      memory[2826] <=  8'h00;      memory[2827] <=  8'h00;      memory[2828] <=  8'h00;      memory[2829] <=  8'h00;      memory[2830] <=  8'h00;      memory[2831] <=  8'h00;      memory[2832] <=  8'h00;      memory[2833] <=  8'h00;      memory[2834] <=  8'h00;      memory[2835] <=  8'h00;      memory[2836] <=  8'h00;      memory[2837] <=  8'h00;      memory[2838] <=  8'h00;      memory[2839] <=  8'h00;      memory[2840] <=  8'h00;      memory[2841] <=  8'h00;      memory[2842] <=  8'h00;      memory[2843] <=  8'h00;      memory[2844] <=  8'h00;      memory[2845] <=  8'h00;      memory[2846] <=  8'h00;      memory[2847] <=  8'h00;      memory[2848] <=  8'h00;      memory[2849] <=  8'h00;      memory[2850] <=  8'h00;      memory[2851] <=  8'h00;      memory[2852] <=  8'h00;      memory[2853] <=  8'h00;      memory[2854] <=  8'h00;      memory[2855] <=  8'h00;      memory[2856] <=  8'h00;      memory[2857] <=  8'h00;      memory[2858] <=  8'h00;      memory[2859] <=  8'h00;      memory[2860] <=  8'h00;      memory[2861] <=  8'h00;      memory[2862] <=  8'h00;      memory[2863] <=  8'h00;      memory[2864] <=  8'h00;      memory[2865] <=  8'h00;      memory[2866] <=  8'h00;      memory[2867] <=  8'h00;      memory[2868] <=  8'h00;      memory[2869] <=  8'h00;      memory[2870] <=  8'h00;      memory[2871] <=  8'h00;      memory[2872] <=  8'h00;      memory[2873] <=  8'h00;      memory[2874] <=  8'h00;      memory[2875] <=  8'h00;      memory[2876] <=  8'h00;      memory[2877] <=  8'h00;      memory[2878] <=  8'h00;      memory[2879] <=  8'h00;      memory[2880] <=  8'h00;      memory[2881] <=  8'h00;      memory[2882] <=  8'h00;      memory[2883] <=  8'h00;      memory[2884] <=  8'h00;      memory[2885] <=  8'h00;      memory[2886] <=  8'h00;      memory[2887] <=  8'h00;      memory[2888] <=  8'h00;      memory[2889] <=  8'h00;      memory[2890] <=  8'h00;      memory[2891] <=  8'h00;      memory[2892] <=  8'h00;      memory[2893] <=  8'h00;      memory[2894] <=  8'h00;      memory[2895] <=  8'h00;      memory[2896] <=  8'h00;      memory[2897] <=  8'h00;      memory[2898] <=  8'h00;      memory[2899] <=  8'h00;      memory[2900] <=  8'h00;      memory[2901] <=  8'h00;      memory[2902] <=  8'h00;      memory[2903] <=  8'h00;      memory[2904] <=  8'h00;      memory[2905] <=  8'h00;      memory[2906] <=  8'h00;      memory[2907] <=  8'h00;      memory[2908] <=  8'h00;      memory[2909] <=  8'h00;      memory[2910] <=  8'h00;      memory[2911] <=  8'h00;      memory[2912] <=  8'h00;      memory[2913] <=  8'h00;      memory[2914] <=  8'h00;      memory[2915] <=  8'h00;      memory[2916] <=  8'h00;      memory[2917] <=  8'h00;      memory[2918] <=  8'h00;      memory[2919] <=  8'h00;      memory[2920] <=  8'h00;      memory[2921] <=  8'h00;      memory[2922] <=  8'h00;      memory[2923] <=  8'h00;      memory[2924] <=  8'h00;      memory[2925] <=  8'h00;      memory[2926] <=  8'h00;      memory[2927] <=  8'h00;      memory[2928] <=  8'h00;      memory[2929] <=  8'h00;      memory[2930] <=  8'h00;      memory[2931] <=  8'h00;      memory[2932] <=  8'h00;      memory[2933] <=  8'h00;      memory[2934] <=  8'h00;      memory[2935] <=  8'h00;      memory[2936] <=  8'h00;      memory[2937] <=  8'h00;      memory[2938] <=  8'h00;      memory[2939] <=  8'h00;      memory[2940] <=  8'h00;      memory[2941] <=  8'h00;      memory[2942] <=  8'h00;      memory[2943] <=  8'h00;      memory[2944] <=  8'h00;      memory[2945] <=  8'h00;      memory[2946] <=  8'h00;      memory[2947] <=  8'h00;      memory[2948] <=  8'h00;      memory[2949] <=  8'h00;      memory[2950] <=  8'h00;      memory[2951] <=  8'h00;      memory[2952] <=  8'h00;      memory[2953] <=  8'h00;      memory[2954] <=  8'h00;      memory[2955] <=  8'h00;      memory[2956] <=  8'h00;      memory[2957] <=  8'h00;      memory[2958] <=  8'h00;      memory[2959] <=  8'h00;      memory[2960] <=  8'h00;      memory[2961] <=  8'h00;      memory[2962] <=  8'h00;      memory[2963] <=  8'h00;      memory[2964] <=  8'h00;      memory[2965] <=  8'h00;      memory[2966] <=  8'h00;      memory[2967] <=  8'h00;      memory[2968] <=  8'h00;      memory[2969] <=  8'h00;      memory[2970] <=  8'h00;      memory[2971] <=  8'h00;      memory[2972] <=  8'h00;      memory[2973] <=  8'h00;      memory[2974] <=  8'h00;      memory[2975] <=  8'h00;      memory[2976] <=  8'h00;      memory[2977] <=  8'h00;      memory[2978] <=  8'h00;      memory[2979] <=  8'h00;      memory[2980] <=  8'h00;      memory[2981] <=  8'h00;      memory[2982] <=  8'h00;      memory[2983] <=  8'h00;      memory[2984] <=  8'h00;      memory[2985] <=  8'h00;      memory[2986] <=  8'h00;      memory[2987] <=  8'h00;      memory[2988] <=  8'h00;      memory[2989] <=  8'h00;      memory[2990] <=  8'h00;      memory[2991] <=  8'h00;      memory[2992] <=  8'h00;      memory[2993] <=  8'h00;      memory[2994] <=  8'h00;      memory[2995] <=  8'h00;      memory[2996] <=  8'h00;      memory[2997] <=  8'h00;      memory[2998] <=  8'h00;      memory[2999] <=  8'h00;      memory[3000] <=  8'h00;      memory[3001] <=  8'h00;      memory[3002] <=  8'h00;      memory[3003] <=  8'h00;      memory[3004] <=  8'h00;      memory[3005] <=  8'h00;      memory[3006] <=  8'h00;      memory[3007] <=  8'h00;      memory[3008] <=  8'h00;      memory[3009] <=  8'h00;      memory[3010] <=  8'h00;      memory[3011] <=  8'h00;      memory[3012] <=  8'h00;      memory[3013] <=  8'h00;      memory[3014] <=  8'h00;      memory[3015] <=  8'h00;      memory[3016] <=  8'h00;      memory[3017] <=  8'h00;      memory[3018] <=  8'h00;      memory[3019] <=  8'h00;      memory[3020] <=  8'h00;      memory[3021] <=  8'h00;      memory[3022] <=  8'h00;      memory[3023] <=  8'h00;      memory[3024] <=  8'h00;      memory[3025] <=  8'h00;      memory[3026] <=  8'h00;      memory[3027] <=  8'h00;      memory[3028] <=  8'h00;      memory[3029] <=  8'h00;      memory[3030] <=  8'h00;      memory[3031] <=  8'h00;      memory[3032] <=  8'h00;      memory[3033] <=  8'h00;      memory[3034] <=  8'h00;      memory[3035] <=  8'h00;      memory[3036] <=  8'h00;      memory[3037] <=  8'h00;      memory[3038] <=  8'h00;      memory[3039] <=  8'h00;      memory[3040] <=  8'h00;      memory[3041] <=  8'h00;      memory[3042] <=  8'h00;      memory[3043] <=  8'h00;      memory[3044] <=  8'h00;      memory[3045] <=  8'h00;      memory[3046] <=  8'h00;      memory[3047] <=  8'h00;      memory[3048] <=  8'h00;      memory[3049] <=  8'h00;      memory[3050] <=  8'h00;      memory[3051] <=  8'h00;      memory[3052] <=  8'h00;      memory[3053] <=  8'h00;      memory[3054] <=  8'h00;      memory[3055] <=  8'h00;      memory[3056] <=  8'h00;      memory[3057] <=  8'h00;      memory[3058] <=  8'h00;      memory[3059] <=  8'h00;      memory[3060] <=  8'h00;      memory[3061] <=  8'h00;      memory[3062] <=  8'h00;      memory[3063] <=  8'h00;      memory[3064] <=  8'h00;      memory[3065] <=  8'h00;      memory[3066] <=  8'h00;      memory[3067] <=  8'h00;      memory[3068] <=  8'h00;      memory[3069] <=  8'h00;      memory[3070] <=  8'h00;      memory[3071] <=  8'h00;      memory[3072] <=  8'h00;      memory[3073] <=  8'h00;      memory[3074] <=  8'h00;      memory[3075] <=  8'h00;      memory[3076] <=  8'h00;      memory[3077] <=  8'h00;      memory[3078] <=  8'h00;      memory[3079] <=  8'h00;      memory[3080] <=  8'h00;      memory[3081] <=  8'h00;      memory[3082] <=  8'h00;      memory[3083] <=  8'h00;      memory[3084] <=  8'h00;      memory[3085] <=  8'h00;      memory[3086] <=  8'h00;      memory[3087] <=  8'h00;      memory[3088] <=  8'h00;      memory[3089] <=  8'h00;      memory[3090] <=  8'h00;      memory[3091] <=  8'h00;      memory[3092] <=  8'h00;      memory[3093] <=  8'h00;      memory[3094] <=  8'h00;      memory[3095] <=  8'h00;      memory[3096] <=  8'h00;      memory[3097] <=  8'h00;      memory[3098] <=  8'h00;      memory[3099] <=  8'h00;      memory[3100] <=  8'h00;      memory[3101] <=  8'h00;      memory[3102] <=  8'h00;      memory[3103] <=  8'h00;      memory[3104] <=  8'h00;      memory[3105] <=  8'h00;      memory[3106] <=  8'h00;      memory[3107] <=  8'h00;      memory[3108] <=  8'h00;      memory[3109] <=  8'h00;      memory[3110] <=  8'h00;      memory[3111] <=  8'h00;      memory[3112] <=  8'h00;      memory[3113] <=  8'h00;      memory[3114] <=  8'h00;      memory[3115] <=  8'h00;      memory[3116] <=  8'h00;      memory[3117] <=  8'h00;      memory[3118] <=  8'h00;      memory[3119] <=  8'h00;      memory[3120] <=  8'h00;      memory[3121] <=  8'h00;      memory[3122] <=  8'h00;      memory[3123] <=  8'h00;      memory[3124] <=  8'h00;      memory[3125] <=  8'h00;      memory[3126] <=  8'h00;      memory[3127] <=  8'h00;      memory[3128] <=  8'h00;      memory[3129] <=  8'h00;      memory[3130] <=  8'h00;      memory[3131] <=  8'h00;      memory[3132] <=  8'h00;      memory[3133] <=  8'h00;      memory[3134] <=  8'h00;      memory[3135] <=  8'h00;      memory[3136] <=  8'h00;      memory[3137] <=  8'h00;      memory[3138] <=  8'h00;      memory[3139] <=  8'h00;      memory[3140] <=  8'h00;      memory[3141] <=  8'h00;      memory[3142] <=  8'h00;      memory[3143] <=  8'h00;      memory[3144] <=  8'h00;      memory[3145] <=  8'h00;      memory[3146] <=  8'h00;      memory[3147] <=  8'h00;      memory[3148] <=  8'h00;      memory[3149] <=  8'h00;      memory[3150] <=  8'h00;      memory[3151] <=  8'h00;      memory[3152] <=  8'h00;      memory[3153] <=  8'h00;      memory[3154] <=  8'h00;      memory[3155] <=  8'h00;      memory[3156] <=  8'h00;      memory[3157] <=  8'h00;      memory[3158] <=  8'h00;      memory[3159] <=  8'h00;      memory[3160] <=  8'h00;      memory[3161] <=  8'h00;      memory[3162] <=  8'h00;      memory[3163] <=  8'h00;      memory[3164] <=  8'h00;      memory[3165] <=  8'h00;      memory[3166] <=  8'h00;      memory[3167] <=  8'h00;      memory[3168] <=  8'h00;      memory[3169] <=  8'h00;      memory[3170] <=  8'h00;      memory[3171] <=  8'h00;      memory[3172] <=  8'h00;      memory[3173] <=  8'h00;      memory[3174] <=  8'h00;      memory[3175] <=  8'h00;      memory[3176] <=  8'h00;      memory[3177] <=  8'h00;      memory[3178] <=  8'h00;      memory[3179] <=  8'h00;      memory[3180] <=  8'h00;      memory[3181] <=  8'h00;      memory[3182] <=  8'h00;      memory[3183] <=  8'h00;      memory[3184] <=  8'h00;      memory[3185] <=  8'h00;      memory[3186] <=  8'h00;      memory[3187] <=  8'h00;      memory[3188] <=  8'h00;      memory[3189] <=  8'h00;      memory[3190] <=  8'h00;      memory[3191] <=  8'h00;      memory[3192] <=  8'h00;      memory[3193] <=  8'h00;      memory[3194] <=  8'h00;      memory[3195] <=  8'h00;      memory[3196] <=  8'h00;      memory[3197] <=  8'h00;      memory[3198] <=  8'h00;      memory[3199] <=  8'h00;      memory[3200] <=  8'h00;      memory[3201] <=  8'h00;      memory[3202] <=  8'h00;      memory[3203] <=  8'h00;      memory[3204] <=  8'h00;      memory[3205] <=  8'h00;      memory[3206] <=  8'h00;      memory[3207] <=  8'h00;      memory[3208] <=  8'h00;      memory[3209] <=  8'h00;      memory[3210] <=  8'h00;      memory[3211] <=  8'h00;      memory[3212] <=  8'h00;      memory[3213] <=  8'h00;      memory[3214] <=  8'h00;      memory[3215] <=  8'h00;      memory[3216] <=  8'h00;      memory[3217] <=  8'h00;      memory[3218] <=  8'h00;      memory[3219] <=  8'h00;      memory[3220] <=  8'h00;      memory[3221] <=  8'h00;      memory[3222] <=  8'h00;      memory[3223] <=  8'h00;      memory[3224] <=  8'h00;      memory[3225] <=  8'h00;      memory[3226] <=  8'h00;      memory[3227] <=  8'h00;      memory[3228] <=  8'h00;      memory[3229] <=  8'h00;      memory[3230] <=  8'h00;      memory[3231] <=  8'h00;      memory[3232] <=  8'h00;      memory[3233] <=  8'h00;      memory[3234] <=  8'h00;      memory[3235] <=  8'h00;      memory[3236] <=  8'h00;      memory[3237] <=  8'h00;      memory[3238] <=  8'h00;      memory[3239] <=  8'h00;      memory[3240] <=  8'h00;      memory[3241] <=  8'h00;      memory[3242] <=  8'h00;      memory[3243] <=  8'h00;      memory[3244] <=  8'h00;      memory[3245] <=  8'h00;      memory[3246] <=  8'h00;      memory[3247] <=  8'h00;      memory[3248] <=  8'h00;      memory[3249] <=  8'h00;      memory[3250] <=  8'h00;      memory[3251] <=  8'h00;      memory[3252] <=  8'h00;      memory[3253] <=  8'h00;      memory[3254] <=  8'h00;      memory[3255] <=  8'h00;      memory[3256] <=  8'h00;      memory[3257] <=  8'h00;      memory[3258] <=  8'h00;      memory[3259] <=  8'h00;      memory[3260] <=  8'h00;      memory[3261] <=  8'h00;      memory[3262] <=  8'h00;      memory[3263] <=  8'h00;      memory[3264] <=  8'h00;      memory[3265] <=  8'h00;      memory[3266] <=  8'h00;      memory[3267] <=  8'h00;      memory[3268] <=  8'h00;      memory[3269] <=  8'h00;      memory[3270] <=  8'h00;      memory[3271] <=  8'h00;      memory[3272] <=  8'h00;      memory[3273] <=  8'h00;      memory[3274] <=  8'h00;      memory[3275] <=  8'h00;      memory[3276] <=  8'h00;      memory[3277] <=  8'h00;      memory[3278] <=  8'h00;      memory[3279] <=  8'h00;      memory[3280] <=  8'h00;      memory[3281] <=  8'h00;      memory[3282] <=  8'h00;      memory[3283] <=  8'h00;      memory[3284] <=  8'h00;      memory[3285] <=  8'h00;      memory[3286] <=  8'h00;      memory[3287] <=  8'h00;      memory[3288] <=  8'h00;      memory[3289] <=  8'h00;      memory[3290] <=  8'h00;      memory[3291] <=  8'h00;      memory[3292] <=  8'h00;      memory[3293] <=  8'h00;      memory[3294] <=  8'h00;      memory[3295] <=  8'h00;      memory[3296] <=  8'h00;      memory[3297] <=  8'h00;      memory[3298] <=  8'h00;      memory[3299] <=  8'h00;      memory[3300] <=  8'h00;      memory[3301] <=  8'h00;      memory[3302] <=  8'h00;      memory[3303] <=  8'h00;      memory[3304] <=  8'h00;      memory[3305] <=  8'h00;      memory[3306] <=  8'h00;      memory[3307] <=  8'h00;      memory[3308] <=  8'h00;      memory[3309] <=  8'h00;      memory[3310] <=  8'h00;      memory[3311] <=  8'h00;      memory[3312] <=  8'h00;      memory[3313] <=  8'h00;      memory[3314] <=  8'h00;      memory[3315] <=  8'h00;      memory[3316] <=  8'h00;      memory[3317] <=  8'h00;      memory[3318] <=  8'h00;      memory[3319] <=  8'h00;      memory[3320] <=  8'h00;      memory[3321] <=  8'h00;      memory[3322] <=  8'h00;      memory[3323] <=  8'h00;      memory[3324] <=  8'h00;      memory[3325] <=  8'h00;      memory[3326] <=  8'h00;      memory[3327] <=  8'h00;      memory[3328] <=  8'h00;      memory[3329] <=  8'h00;      memory[3330] <=  8'h00;      memory[3331] <=  8'h00;      memory[3332] <=  8'h00;      memory[3333] <=  8'h00;      memory[3334] <=  8'h00;      memory[3335] <=  8'h00;      memory[3336] <=  8'h00;      memory[3337] <=  8'h00;      memory[3338] <=  8'h00;      memory[3339] <=  8'h00;      memory[3340] <=  8'h00;      memory[3341] <=  8'h00;      memory[3342] <=  8'h00;      memory[3343] <=  8'h00;      memory[3344] <=  8'h00;      memory[3345] <=  8'h00;      memory[3346] <=  8'h00;      memory[3347] <=  8'h00;      memory[3348] <=  8'h00;      memory[3349] <=  8'h00;      memory[3350] <=  8'h00;      memory[3351] <=  8'h00;      memory[3352] <=  8'h00;      memory[3353] <=  8'h00;      memory[3354] <=  8'h00;      memory[3355] <=  8'h00;      memory[3356] <=  8'h00;      memory[3357] <=  8'h00;      memory[3358] <=  8'h00;      memory[3359] <=  8'h00;      memory[3360] <=  8'h00;      memory[3361] <=  8'h00;      memory[3362] <=  8'h00;      memory[3363] <=  8'h00;      memory[3364] <=  8'h00;      memory[3365] <=  8'h00;      memory[3366] <=  8'h00;      memory[3367] <=  8'h00;      memory[3368] <=  8'h00;      memory[3369] <=  8'h00;      memory[3370] <=  8'h00;      memory[3371] <=  8'h00;      memory[3372] <=  8'h00;      memory[3373] <=  8'h00;      memory[3374] <=  8'h00;      memory[3375] <=  8'h00;      memory[3376] <=  8'h00;      memory[3377] <=  8'h00;      memory[3378] <=  8'h00;      memory[3379] <=  8'h00;      memory[3380] <=  8'h00;      memory[3381] <=  8'h00;      memory[3382] <=  8'h00;      memory[3383] <=  8'h00;      memory[3384] <=  8'h00;      memory[3385] <=  8'h00;      memory[3386] <=  8'h00;      memory[3387] <=  8'h00;      memory[3388] <=  8'h00;      memory[3389] <=  8'h00;      memory[3390] <=  8'h00;      memory[3391] <=  8'h00;      memory[3392] <=  8'h00;      memory[3393] <=  8'h00;      memory[3394] <=  8'h00;      memory[3395] <=  8'h00;      memory[3396] <=  8'h00;      memory[3397] <=  8'h00;      memory[3398] <=  8'h00;      memory[3399] <=  8'h00;      memory[3400] <=  8'h00;      memory[3401] <=  8'h00;      memory[3402] <=  8'h00;      memory[3403] <=  8'h00;      memory[3404] <=  8'h00;      memory[3405] <=  8'h00;      memory[3406] <=  8'h00;      memory[3407] <=  8'h00;      memory[3408] <=  8'h00;      memory[3409] <=  8'h00;      memory[3410] <=  8'h00;      memory[3411] <=  8'h00;      memory[3412] <=  8'h00;      memory[3413] <=  8'h00;      memory[3414] <=  8'h00;      memory[3415] <=  8'h00;      memory[3416] <=  8'h00;      memory[3417] <=  8'h00;      memory[3418] <=  8'h00;      memory[3419] <=  8'h00;      memory[3420] <=  8'h00;      memory[3421] <=  8'h00;      memory[3422] <=  8'h00;      memory[3423] <=  8'h00;      memory[3424] <=  8'h00;      memory[3425] <=  8'h00;      memory[3426] <=  8'h00;      memory[3427] <=  8'h00;      memory[3428] <=  8'h00;      memory[3429] <=  8'h00;      memory[3430] <=  8'h00;      memory[3431] <=  8'h00;      memory[3432] <=  8'h00;      memory[3433] <=  8'h00;      memory[3434] <=  8'h00;      memory[3435] <=  8'h00;      memory[3436] <=  8'h00;      memory[3437] <=  8'h00;      memory[3438] <=  8'h00;      memory[3439] <=  8'h00;      memory[3440] <=  8'h00;      memory[3441] <=  8'h00;      memory[3442] <=  8'h00;      memory[3443] <=  8'h00;      memory[3444] <=  8'h00;      memory[3445] <=  8'h00;      memory[3446] <=  8'h00;      memory[3447] <=  8'h00;      memory[3448] <=  8'h00;      memory[3449] <=  8'h00;      memory[3450] <=  8'h00;      memory[3451] <=  8'h00;      memory[3452] <=  8'h00;      memory[3453] <=  8'h00;      memory[3454] <=  8'h00;      memory[3455] <=  8'h00;      memory[3456] <=  8'h00;      memory[3457] <=  8'h00;      memory[3458] <=  8'h00;      memory[3459] <=  8'h00;      memory[3460] <=  8'h00;      memory[3461] <=  8'h00;      memory[3462] <=  8'h00;      memory[3463] <=  8'h00;      memory[3464] <=  8'h00;      memory[3465] <=  8'h00;      memory[3466] <=  8'h00;      memory[3467] <=  8'h00;      memory[3468] <=  8'h00;      memory[3469] <=  8'h00;      memory[3470] <=  8'h00;      memory[3471] <=  8'h00;      memory[3472] <=  8'h00;      memory[3473] <=  8'h00;      memory[3474] <=  8'h00;      memory[3475] <=  8'h00;      memory[3476] <=  8'h00;      memory[3477] <=  8'h00;      memory[3478] <=  8'h00;      memory[3479] <=  8'h00;      memory[3480] <=  8'h00;      memory[3481] <=  8'h00;      memory[3482] <=  8'h00;      memory[3483] <=  8'h00;      memory[3484] <=  8'h00;      memory[3485] <=  8'h00;      memory[3486] <=  8'h00;      memory[3487] <=  8'h00;      memory[3488] <=  8'h00;      memory[3489] <=  8'h00;      memory[3490] <=  8'h00;      memory[3491] <=  8'h00;      memory[3492] <=  8'h00;      memory[3493] <=  8'h00;      memory[3494] <=  8'h00;      memory[3495] <=  8'h00;      memory[3496] <=  8'h00;      memory[3497] <=  8'h00;      memory[3498] <=  8'h00;      memory[3499] <=  8'h00;      memory[3500] <=  8'h00;      memory[3501] <=  8'h00;      memory[3502] <=  8'h00;      memory[3503] <=  8'h00;      memory[3504] <=  8'h00;      memory[3505] <=  8'h00;      memory[3506] <=  8'h00;      memory[3507] <=  8'h00;      memory[3508] <=  8'h00;      memory[3509] <=  8'h00;      memory[3510] <=  8'h00;      memory[3511] <=  8'h00;      memory[3512] <=  8'h00;      memory[3513] <=  8'h00;      memory[3514] <=  8'h00;      memory[3515] <=  8'h00;      memory[3516] <=  8'h00;      memory[3517] <=  8'h00;      memory[3518] <=  8'h00;      memory[3519] <=  8'h00;      memory[3520] <=  8'h00;      memory[3521] <=  8'h00;      memory[3522] <=  8'h00;      memory[3523] <=  8'h00;      memory[3524] <=  8'h00;      memory[3525] <=  8'h00;      memory[3526] <=  8'h00;      memory[3527] <=  8'h00;      memory[3528] <=  8'h00;      memory[3529] <=  8'h00;      memory[3530] <=  8'h00;      memory[3531] <=  8'h00;      memory[3532] <=  8'h00;      memory[3533] <=  8'h00;      memory[3534] <=  8'h00;      memory[3535] <=  8'h00;      memory[3536] <=  8'h00;      memory[3537] <=  8'h00;      memory[3538] <=  8'h00;      memory[3539] <=  8'h00;      memory[3540] <=  8'h00;      memory[3541] <=  8'h00;      memory[3542] <=  8'h00;      memory[3543] <=  8'h00;      memory[3544] <=  8'h00;      memory[3545] <=  8'h00;      memory[3546] <=  8'h00;      memory[3547] <=  8'h00;      memory[3548] <=  8'h00;      memory[3549] <=  8'h00;      memory[3550] <=  8'h00;      memory[3551] <=  8'h00;      memory[3552] <=  8'h00;      memory[3553] <=  8'h00;      memory[3554] <=  8'h00;      memory[3555] <=  8'h00;      memory[3556] <=  8'h00;      memory[3557] <=  8'h00;      memory[3558] <=  8'h00;      memory[3559] <=  8'h00;      memory[3560] <=  8'h00;      memory[3561] <=  8'h00;      memory[3562] <=  8'h00;      memory[3563] <=  8'h00;      memory[3564] <=  8'h00;      memory[3565] <=  8'h00;      memory[3566] <=  8'h00;      memory[3567] <=  8'h00;      memory[3568] <=  8'h00;      memory[3569] <=  8'h00;      memory[3570] <=  8'h00;      memory[3571] <=  8'h00;      memory[3572] <=  8'h00;      memory[3573] <=  8'h00;      memory[3574] <=  8'h00;      memory[3575] <=  8'h00;      memory[3576] <=  8'h00;      memory[3577] <=  8'h00;      memory[3578] <=  8'h00;      memory[3579] <=  8'h00;      memory[3580] <=  8'h00;      memory[3581] <=  8'h00;      memory[3582] <=  8'h00;      memory[3583] <=  8'h00;      memory[3584] <=  8'h00;      memory[3585] <=  8'h00;      memory[3586] <=  8'h00;      memory[3587] <=  8'h00;      memory[3588] <=  8'h00;      memory[3589] <=  8'h00;      memory[3590] <=  8'h00;      memory[3591] <=  8'h00;      memory[3592] <=  8'h00;      memory[3593] <=  8'h00;      memory[3594] <=  8'h00;      memory[3595] <=  8'h00;      memory[3596] <=  8'h00;      memory[3597] <=  8'h00;      memory[3598] <=  8'h00;      memory[3599] <=  8'h00;      memory[3600] <=  8'h00;      memory[3601] <=  8'h00;      memory[3602] <=  8'h00;      memory[3603] <=  8'h00;      memory[3604] <=  8'h00;      memory[3605] <=  8'h00;      memory[3606] <=  8'h00;      memory[3607] <=  8'h00;      memory[3608] <=  8'h00;      memory[3609] <=  8'h00;      memory[3610] <=  8'h00;      memory[3611] <=  8'h00;      memory[3612] <=  8'h00;      memory[3613] <=  8'h00;      memory[3614] <=  8'h00;      memory[3615] <=  8'h00;      memory[3616] <=  8'h00;      memory[3617] <=  8'h00;      memory[3618] <=  8'h00;      memory[3619] <=  8'h00;      memory[3620] <=  8'h00;      memory[3621] <=  8'h00;      memory[3622] <=  8'h00;      memory[3623] <=  8'h00;      memory[3624] <=  8'h00;      memory[3625] <=  8'h00;      memory[3626] <=  8'h00;      memory[3627] <=  8'h00;      memory[3628] <=  8'h00;      memory[3629] <=  8'h00;      memory[3630] <=  8'h00;      memory[3631] <=  8'h00;      memory[3632] <=  8'h00;      memory[3633] <=  8'h00;      memory[3634] <=  8'h00;      memory[3635] <=  8'h00;      memory[3636] <=  8'h00;      memory[3637] <=  8'h00;      memory[3638] <=  8'h00;      memory[3639] <=  8'h00;      memory[3640] <=  8'h00;      memory[3641] <=  8'h00;      memory[3642] <=  8'h00;      memory[3643] <=  8'h00;      memory[3644] <=  8'h00;      memory[3645] <=  8'h00;      memory[3646] <=  8'h00;      memory[3647] <=  8'h00;      memory[3648] <=  8'h00;      memory[3649] <=  8'h00;      memory[3650] <=  8'h00;      memory[3651] <=  8'h00;      memory[3652] <=  8'h00;      memory[3653] <=  8'h00;      memory[3654] <=  8'h00;      memory[3655] <=  8'h00;      memory[3656] <=  8'h00;      memory[3657] <=  8'h00;      memory[3658] <=  8'h00;      memory[3659] <=  8'h00;      memory[3660] <=  8'h00;      memory[3661] <=  8'h00;      memory[3662] <=  8'h00;      memory[3663] <=  8'h00;      memory[3664] <=  8'h00;      memory[3665] <=  8'h00;      memory[3666] <=  8'h00;      memory[3667] <=  8'h00;      memory[3668] <=  8'h00;      memory[3669] <=  8'h00;      memory[3670] <=  8'h00;      memory[3671] <=  8'h00;      memory[3672] <=  8'h00;      memory[3673] <=  8'h00;      memory[3674] <=  8'h00;      memory[3675] <=  8'h00;      memory[3676] <=  8'h00;      memory[3677] <=  8'h00;      memory[3678] <=  8'h00;      memory[3679] <=  8'h00;      memory[3680] <=  8'h00;      memory[3681] <=  8'h00;      memory[3682] <=  8'h00;      memory[3683] <=  8'h00;      memory[3684] <=  8'h00;      memory[3685] <=  8'h00;      memory[3686] <=  8'h00;      memory[3687] <=  8'h00;      memory[3688] <=  8'h00;      memory[3689] <=  8'h00;      memory[3690] <=  8'h00;      memory[3691] <=  8'h00;      memory[3692] <=  8'h00;      memory[3693] <=  8'h00;      memory[3694] <=  8'h00;      memory[3695] <=  8'h00;      memory[3696] <=  8'h00;      memory[3697] <=  8'h00;      memory[3698] <=  8'h00;      memory[3699] <=  8'h00;      memory[3700] <=  8'h00;      memory[3701] <=  8'h00;      memory[3702] <=  8'h00;      memory[3703] <=  8'h00;      memory[3704] <=  8'h00;      memory[3705] <=  8'h00;      memory[3706] <=  8'h00;      memory[3707] <=  8'h00;      memory[3708] <=  8'h00;      memory[3709] <=  8'h00;      memory[3710] <=  8'h00;      memory[3711] <=  8'h00;      memory[3712] <=  8'h00;      memory[3713] <=  8'h00;      memory[3714] <=  8'h00;      memory[3715] <=  8'h00;      memory[3716] <=  8'h00;      memory[3717] <=  8'h00;      memory[3718] <=  8'h00;      memory[3719] <=  8'h00;      memory[3720] <=  8'h00;      memory[3721] <=  8'h00;      memory[3722] <=  8'h00;      memory[3723] <=  8'h00;      memory[3724] <=  8'h00;      memory[3725] <=  8'h00;      memory[3726] <=  8'h00;      memory[3727] <=  8'h00;      memory[3728] <=  8'h00;      memory[3729] <=  8'h00;      memory[3730] <=  8'h00;      memory[3731] <=  8'h00;      memory[3732] <=  8'h00;      memory[3733] <=  8'h00;      memory[3734] <=  8'h00;      memory[3735] <=  8'h00;      memory[3736] <=  8'h00;      memory[3737] <=  8'h00;      memory[3738] <=  8'h00;      memory[3739] <=  8'h00;      memory[3740] <=  8'h00;      memory[3741] <=  8'h00;      memory[3742] <=  8'h00;      memory[3743] <=  8'h00;      memory[3744] <=  8'h00;      memory[3745] <=  8'h00;      memory[3746] <=  8'h00;      memory[3747] <=  8'h00;      memory[3748] <=  8'h00;      memory[3749] <=  8'h00;      memory[3750] <=  8'h00;      memory[3751] <=  8'h00;      memory[3752] <=  8'h00;      memory[3753] <=  8'h00;      memory[3754] <=  8'h00;      memory[3755] <=  8'h00;      memory[3756] <=  8'h00;      memory[3757] <=  8'h00;      memory[3758] <=  8'h00;      memory[3759] <=  8'h00;      memory[3760] <=  8'h00;      memory[3761] <=  8'h00;      memory[3762] <=  8'h00;      memory[3763] <=  8'h00;      memory[3764] <=  8'h00;      memory[3765] <=  8'h00;      memory[3766] <=  8'h00;      memory[3767] <=  8'h00;      memory[3768] <=  8'h00;      memory[3769] <=  8'h00;      memory[3770] <=  8'h00;      memory[3771] <=  8'h00;      memory[3772] <=  8'h00;      memory[3773] <=  8'h00;      memory[3774] <=  8'h00;      memory[3775] <=  8'h00;      memory[3776] <=  8'h00;      memory[3777] <=  8'h00;      memory[3778] <=  8'h00;      memory[3779] <=  8'h00;      memory[3780] <=  8'h00;      memory[3781] <=  8'h00;      memory[3782] <=  8'h00;      memory[3783] <=  8'h00;      memory[3784] <=  8'h00;      memory[3785] <=  8'h00;      memory[3786] <=  8'h00;      memory[3787] <=  8'h00;      memory[3788] <=  8'h00;      memory[3789] <=  8'h00;      memory[3790] <=  8'h00;      memory[3791] <=  8'h00;      memory[3792] <=  8'h00;      memory[3793] <=  8'h00;      memory[3794] <=  8'h00;      memory[3795] <=  8'h00;      memory[3796] <=  8'h00;      memory[3797] <=  8'h00;      memory[3798] <=  8'h00;      memory[3799] <=  8'h00;      memory[3800] <=  8'h00;      memory[3801] <=  8'h00;      memory[3802] <=  8'h00;      memory[3803] <=  8'h00;      memory[3804] <=  8'h00;      memory[3805] <=  8'h00;      memory[3806] <=  8'h00;      memory[3807] <=  8'h00;      memory[3808] <=  8'h00;      memory[3809] <=  8'h00;      memory[3810] <=  8'h00;      memory[3811] <=  8'h00;      memory[3812] <=  8'h00;      memory[3813] <=  8'h00;      memory[3814] <=  8'h00;      memory[3815] <=  8'h00;      memory[3816] <=  8'h00;      memory[3817] <=  8'h00;      memory[3818] <=  8'h00;      memory[3819] <=  8'h00;      memory[3820] <=  8'h00;      memory[3821] <=  8'h00;      memory[3822] <=  8'h00;      memory[3823] <=  8'h00;      memory[3824] <=  8'h00;      memory[3825] <=  8'h00;      memory[3826] <=  8'h00;      memory[3827] <=  8'h00;      memory[3828] <=  8'h00;      memory[3829] <=  8'h00;      memory[3830] <=  8'h00;      memory[3831] <=  8'h00;      memory[3832] <=  8'h00;      memory[3833] <=  8'h00;      memory[3834] <=  8'h00;      memory[3835] <=  8'h00;      memory[3836] <=  8'h00;      memory[3837] <=  8'h00;      memory[3838] <=  8'h00;      memory[3839] <=  8'h00;      memory[3840] <=  8'h00;      memory[3841] <=  8'h00;      memory[3842] <=  8'h00;      memory[3843] <=  8'h00;      memory[3844] <=  8'h00;      memory[3845] <=  8'h00;      memory[3846] <=  8'h00;      memory[3847] <=  8'h00;      memory[3848] <=  8'h00;      memory[3849] <=  8'h00;      memory[3850] <=  8'h00;      memory[3851] <=  8'h00;      memory[3852] <=  8'h00;      memory[3853] <=  8'h00;      memory[3854] <=  8'h00;      memory[3855] <=  8'h00;      memory[3856] <=  8'h00;      memory[3857] <=  8'h00;      memory[3858] <=  8'h00;      memory[3859] <=  8'h00;      memory[3860] <=  8'h00;      memory[3861] <=  8'h00;      memory[3862] <=  8'h00;      memory[3863] <=  8'h00;      memory[3864] <=  8'h00;      memory[3865] <=  8'h00;      memory[3866] <=  8'h00;      memory[3867] <=  8'h00;      memory[3868] <=  8'h00;      memory[3869] <=  8'h00;      memory[3870] <=  8'h00;      memory[3871] <=  8'h00;      memory[3872] <=  8'h00;      memory[3873] <=  8'h00;      memory[3874] <=  8'h00;      memory[3875] <=  8'h00;      memory[3876] <=  8'h00;      memory[3877] <=  8'h00;      memory[3878] <=  8'h00;      memory[3879] <=  8'h00;      memory[3880] <=  8'h00;      memory[3881] <=  8'h00;      memory[3882] <=  8'h00;      memory[3883] <=  8'h00;      memory[3884] <=  8'h00;      memory[3885] <=  8'h00;      memory[3886] <=  8'h00;      memory[3887] <=  8'h00;      memory[3888] <=  8'h00;      memory[3889] <=  8'h00;      memory[3890] <=  8'h00;      memory[3891] <=  8'h00;      memory[3892] <=  8'h00;      memory[3893] <=  8'h00;      memory[3894] <=  8'h00;      memory[3895] <=  8'h00;      memory[3896] <=  8'h00;      memory[3897] <=  8'h00;      memory[3898] <=  8'h00;      memory[3899] <=  8'h00;      memory[3900] <=  8'h00;      memory[3901] <=  8'h00;      memory[3902] <=  8'h00;      memory[3903] <=  8'h00;      memory[3904] <=  8'h00;      memory[3905] <=  8'h00;      memory[3906] <=  8'h00;      memory[3907] <=  8'h00;      memory[3908] <=  8'h00;      memory[3909] <=  8'h00;      memory[3910] <=  8'h00;      memory[3911] <=  8'h00;      memory[3912] <=  8'h00;      memory[3913] <=  8'h00;      memory[3914] <=  8'h00;      memory[3915] <=  8'h00;      memory[3916] <=  8'h00;      memory[3917] <=  8'h00;      memory[3918] <=  8'h00;      memory[3919] <=  8'h00;      memory[3920] <=  8'h00;      memory[3921] <=  8'h00;      memory[3922] <=  8'h00;      memory[3923] <=  8'h00;      memory[3924] <=  8'h00;      memory[3925] <=  8'h00;      memory[3926] <=  8'h00;      memory[3927] <=  8'h00;      memory[3928] <=  8'h00;      memory[3929] <=  8'h00;      memory[3930] <=  8'h00;      memory[3931] <=  8'h00;      memory[3932] <=  8'h00;      memory[3933] <=  8'h00;      memory[3934] <=  8'h00;      memory[3935] <=  8'h00;      memory[3936] <=  8'h00;      memory[3937] <=  8'h00;      memory[3938] <=  8'h00;      memory[3939] <=  8'h00;      memory[3940] <=  8'h00;      memory[3941] <=  8'h00;      memory[3942] <=  8'h00;      memory[3943] <=  8'h00;      memory[3944] <=  8'h00;      memory[3945] <=  8'h00;      memory[3946] <=  8'h00;      memory[3947] <=  8'h00;      memory[3948] <=  8'h00;      memory[3949] <=  8'h00;      memory[3950] <=  8'h00;      memory[3951] <=  8'h00;      memory[3952] <=  8'h00;      memory[3953] <=  8'h00;      memory[3954] <=  8'h00;      memory[3955] <=  8'h00;      memory[3956] <=  8'h00;      memory[3957] <=  8'h00;      memory[3958] <=  8'h00;      memory[3959] <=  8'h00;      memory[3960] <=  8'h00;      memory[3961] <=  8'h00;      memory[3962] <=  8'h00;      memory[3963] <=  8'h00;      memory[3964] <=  8'h00;      memory[3965] <=  8'h00;      memory[3966] <=  8'h00;      memory[3967] <=  8'h00;      memory[3968] <=  8'h00;      memory[3969] <=  8'h00;      memory[3970] <=  8'h00;      memory[3971] <=  8'h00;      memory[3972] <=  8'h00;      memory[3973] <=  8'h00;      memory[3974] <=  8'h00;      memory[3975] <=  8'h00;      memory[3976] <=  8'h00;      memory[3977] <=  8'h00;      memory[3978] <=  8'h00;      memory[3979] <=  8'h00;      memory[3980] <=  8'h00;      memory[3981] <=  8'h00;      memory[3982] <=  8'h00;      memory[3983] <=  8'h00;      memory[3984] <=  8'h00;      memory[3985] <=  8'h00;      memory[3986] <=  8'h00;      memory[3987] <=  8'h00;      memory[3988] <=  8'h00;      memory[3989] <=  8'h00;      memory[3990] <=  8'h00;      memory[3991] <=  8'h00;      memory[3992] <=  8'h00;      memory[3993] <=  8'h00;      memory[3994] <=  8'h00;      memory[3995] <=  8'h00;      memory[3996] <=  8'h00;      memory[3997] <=  8'h00;      memory[3998] <=  8'h00;      memory[3999] <=  8'h00;      memory[4000] <=  8'h00;      memory[4001] <=  8'h00;      memory[4002] <=  8'h00;      memory[4003] <=  8'h00;      memory[4004] <=  8'h00;      memory[4005] <=  8'h00;      memory[4006] <=  8'h00;      memory[4007] <=  8'h00;      memory[4008] <=  8'h00;      memory[4009] <=  8'h00;      memory[4010] <=  8'h00;      memory[4011] <=  8'h00;      memory[4012] <=  8'h00;      memory[4013] <=  8'h00;      memory[4014] <=  8'h00;      memory[4015] <=  8'h00;      memory[4016] <=  8'h00;      memory[4017] <=  8'h00;      memory[4018] <=  8'h00;      memory[4019] <=  8'h00;      memory[4020] <=  8'h00;      memory[4021] <=  8'h00;      memory[4022] <=  8'h00;      memory[4023] <=  8'h00;      memory[4024] <=  8'h00;      memory[4025] <=  8'h00;      memory[4026] <=  8'h00;      memory[4027] <=  8'h00;      memory[4028] <=  8'h00;      memory[4029] <=  8'h00;      memory[4030] <=  8'h00;      memory[4031] <=  8'h00;      memory[4032] <=  8'h00;      memory[4033] <=  8'h00;      memory[4034] <=  8'h00;      memory[4035] <=  8'h00;      memory[4036] <=  8'h00;      memory[4037] <=  8'h00;      memory[4038] <=  8'h00;      memory[4039] <=  8'h00;      memory[4040] <=  8'h00;      memory[4041] <=  8'h00;      memory[4042] <=  8'h00;      memory[4043] <=  8'h00;      memory[4044] <=  8'h00;      memory[4045] <=  8'h00;      memory[4046] <=  8'h00;      memory[4047] <=  8'h00;      memory[4048] <=  8'h00;      memory[4049] <=  8'h00;      memory[4050] <=  8'h00;      memory[4051] <=  8'h00;      memory[4052] <=  8'h00;      memory[4053] <=  8'h00;      memory[4054] <=  8'h00;      memory[4055] <=  8'h00;      memory[4056] <=  8'h00;      memory[4057] <=  8'h00;      memory[4058] <=  8'h00;      memory[4059] <=  8'h00;      memory[4060] <=  8'h00;      memory[4061] <=  8'h00;      memory[4062] <=  8'h00;      memory[4063] <=  8'h00;      memory[4064] <=  8'h00;      memory[4065] <=  8'h00;      memory[4066] <=  8'h00;      memory[4067] <=  8'h00;      memory[4068] <=  8'h00;      memory[4069] <=  8'h00;      memory[4070] <=  8'h00;      memory[4071] <=  8'h00;      memory[4072] <=  8'h00;      memory[4073] <=  8'h00;      memory[4074] <=  8'h00;      memory[4075] <=  8'h00;      memory[4076] <=  8'h00;      memory[4077] <=  8'h00;      memory[4078] <=  8'h00;      memory[4079] <=  8'h00;      memory[4080] <=  8'h00;      memory[4081] <=  8'h00;      memory[4082] <=  8'h00;      memory[4083] <=  8'h00;      memory[4084] <=  8'h00;      memory[4085] <=  8'h00;      memory[4086] <=  8'h00;      memory[4087] <=  8'h00;      memory[4088] <=  8'h00;      memory[4089] <=  8'h00;      memory[4090] <=  8'h00;      memory[4091] <=  8'h00;      memory[4092] <=  8'h00;      memory[4093] <=  8'h00;      memory[4094] <=  8'h00;      memory[4095] <=  8'h00;      memory[4096] <=  8'h00;      memory[4097] <=  8'h00;      memory[4098] <=  8'h00;      memory[4099] <=  8'h00;      memory[4100] <=  8'h00;      memory[4101] <=  8'h00;      memory[4102] <=  8'h00;      memory[4103] <=  8'h00;      memory[4104] <=  8'h00;      memory[4105] <=  8'h00;      memory[4106] <=  8'h00;      memory[4107] <=  8'h00;      memory[4108] <=  8'h00;      memory[4109] <=  8'h00;      memory[4110] <=  8'h00;      memory[4111] <=  8'h00;      memory[4112] <=  8'h00;      memory[4113] <=  8'h00;      memory[4114] <=  8'h00;      memory[4115] <=  8'h00;      memory[4116] <=  8'h00;      memory[4117] <=  8'h00;      memory[4118] <=  8'h00;      memory[4119] <=  8'h00;      memory[4120] <=  8'h00;      memory[4121] <=  8'h00;      memory[4122] <=  8'h00;      memory[4123] <=  8'h00;      memory[4124] <=  8'h00;      memory[4125] <=  8'h00;      memory[4126] <=  8'h00;      memory[4127] <=  8'h00;      memory[4128] <=  8'h00;      memory[4129] <=  8'h00;      memory[4130] <=  8'h00;      memory[4131] <=  8'h00;      memory[4132] <=  8'h00;      memory[4133] <=  8'h00;      memory[4134] <=  8'h00;      memory[4135] <=  8'h00;      memory[4136] <=  8'h00;      memory[4137] <=  8'h00;      memory[4138] <=  8'h00;      memory[4139] <=  8'h00;      memory[4140] <=  8'h00;      memory[4141] <=  8'h00;      memory[4142] <=  8'h00;      memory[4143] <=  8'h00;      memory[4144] <=  8'h00;      memory[4145] <=  8'h00;      memory[4146] <=  8'h00;      memory[4147] <=  8'h00;      memory[4148] <=  8'h00;      memory[4149] <=  8'h00;      memory[4150] <=  8'h00;      memory[4151] <=  8'h00;      memory[4152] <=  8'h00;      memory[4153] <=  8'h00;      memory[4154] <=  8'h00;      memory[4155] <=  8'h00;      memory[4156] <=  8'h00;      memory[4157] <=  8'h00;      memory[4158] <=  8'h00;      memory[4159] <=  8'h00;      memory[4160] <=  8'h00;      memory[4161] <=  8'h00;      memory[4162] <=  8'h00;      memory[4163] <=  8'h00;      memory[4164] <=  8'h00;      memory[4165] <=  8'h00;      memory[4166] <=  8'h00;      memory[4167] <=  8'h00;      memory[4168] <=  8'h00;      memory[4169] <=  8'h00;      memory[4170] <=  8'h00;      memory[4171] <=  8'h00;      memory[4172] <=  8'h00;      memory[4173] <=  8'h00;      memory[4174] <=  8'h00;      memory[4175] <=  8'h00;      memory[4176] <=  8'h00;      memory[4177] <=  8'h00;      memory[4178] <=  8'h00;      memory[4179] <=  8'h00;      memory[4180] <=  8'h00;      memory[4181] <=  8'h00;      memory[4182] <=  8'h00;      memory[4183] <=  8'h00;      memory[4184] <=  8'h00;      memory[4185] <=  8'h00;      memory[4186] <=  8'h00;      memory[4187] <=  8'h00;      memory[4188] <=  8'h00;      memory[4189] <=  8'h00;      memory[4190] <=  8'h00;      memory[4191] <=  8'h00;      memory[4192] <=  8'h00;      memory[4193] <=  8'h00;      memory[4194] <=  8'h00;      memory[4195] <=  8'h00;      memory[4196] <=  8'h00;      memory[4197] <=  8'h00;      memory[4198] <=  8'h00;      memory[4199] <=  8'h00;      memory[4200] <=  8'h00;      memory[4201] <=  8'h00;      memory[4202] <=  8'h00;      memory[4203] <=  8'h00;      memory[4204] <=  8'h00;      memory[4205] <=  8'h00;      memory[4206] <=  8'h00;      memory[4207] <=  8'h00;      memory[4208] <=  8'h00;      memory[4209] <=  8'h00;      memory[4210] <=  8'h00;      memory[4211] <=  8'h00;      memory[4212] <=  8'h00;      memory[4213] <=  8'h00;      memory[4214] <=  8'h00;      memory[4215] <=  8'h00;      memory[4216] <=  8'h00;      memory[4217] <=  8'h00;      memory[4218] <=  8'h00;      memory[4219] <=  8'h00;      memory[4220] <=  8'h00;      memory[4221] <=  8'h00;      memory[4222] <=  8'h00;      memory[4223] <=  8'h00;      memory[4224] <=  8'h00;      memory[4225] <=  8'h00;      memory[4226] <=  8'h00;      memory[4227] <=  8'h00;      memory[4228] <=  8'h00;      memory[4229] <=  8'h00;      memory[4230] <=  8'h00;      memory[4231] <=  8'h00;      memory[4232] <=  8'h00;      memory[4233] <=  8'h00;      memory[4234] <=  8'h00;      memory[4235] <=  8'h00;      memory[4236] <=  8'h00;      memory[4237] <=  8'h00;      memory[4238] <=  8'h00;      memory[4239] <=  8'h00;      memory[4240] <=  8'h00;      memory[4241] <=  8'h00;      memory[4242] <=  8'h00;      memory[4243] <=  8'h00;      memory[4244] <=  8'h00;      memory[4245] <=  8'h00;      memory[4246] <=  8'h00;      memory[4247] <=  8'h00;      memory[4248] <=  8'h00;      memory[4249] <=  8'h00;      memory[4250] <=  8'h00;      memory[4251] <=  8'h00;      memory[4252] <=  8'h00;      memory[4253] <=  8'h00;      memory[4254] <=  8'h00;      memory[4255] <=  8'h00;      memory[4256] <=  8'h00;      memory[4257] <=  8'h00;      memory[4258] <=  8'h00;      memory[4259] <=  8'h00;      memory[4260] <=  8'h00;      memory[4261] <=  8'h00;      memory[4262] <=  8'h00;      memory[4263] <=  8'h00;      memory[4264] <=  8'h00;      memory[4265] <=  8'h00;      memory[4266] <=  8'h00;      memory[4267] <=  8'h00;      memory[4268] <=  8'h00;      memory[4269] <=  8'h00;      memory[4270] <=  8'h00;      memory[4271] <=  8'h00;      memory[4272] <=  8'h00;      memory[4273] <=  8'h00;      memory[4274] <=  8'h00;      memory[4275] <=  8'h00;      memory[4276] <=  8'h00;      memory[4277] <=  8'h00;      memory[4278] <=  8'h00;      memory[4279] <=  8'h00;      memory[4280] <=  8'h00;      memory[4281] <=  8'h00;      memory[4282] <=  8'h00;      memory[4283] <=  8'h00;      memory[4284] <=  8'h00;      memory[4285] <=  8'h00;      memory[4286] <=  8'h00;      memory[4287] <=  8'h00;      memory[4288] <=  8'h00;      memory[4289] <=  8'h00;      memory[4290] <=  8'h00;      memory[4291] <=  8'h00;      memory[4292] <=  8'h00;      memory[4293] <=  8'h00;      memory[4294] <=  8'h00;      memory[4295] <=  8'h00;      memory[4296] <=  8'h00;      memory[4297] <=  8'h00;      memory[4298] <=  8'h00;      memory[4299] <=  8'h00;      memory[4300] <=  8'h00;      memory[4301] <=  8'h00;      memory[4302] <=  8'h00;      memory[4303] <=  8'h00;      memory[4304] <=  8'h00;      memory[4305] <=  8'h00;      memory[4306] <=  8'h00;      memory[4307] <=  8'h00;      memory[4308] <=  8'h00;      memory[4309] <=  8'h00;      memory[4310] <=  8'h00;      memory[4311] <=  8'h00;      memory[4312] <=  8'h00;      memory[4313] <=  8'h00;      memory[4314] <=  8'h00;      memory[4315] <=  8'h00;      memory[4316] <=  8'h00;      memory[4317] <=  8'h00;      memory[4318] <=  8'h00;      memory[4319] <=  8'h00;      memory[4320] <=  8'h00;      memory[4321] <=  8'h00;      memory[4322] <=  8'h00;      memory[4323] <=  8'h00;      memory[4324] <=  8'h00;      memory[4325] <=  8'h00;      memory[4326] <=  8'h00;      memory[4327] <=  8'h00;      memory[4328] <=  8'h00;      memory[4329] <=  8'h00;      memory[4330] <=  8'h00;      memory[4331] <=  8'h00;      memory[4332] <=  8'h00;      memory[4333] <=  8'h00;      memory[4334] <=  8'h00;      memory[4335] <=  8'h00;      memory[4336] <=  8'h00;      memory[4337] <=  8'h00;      memory[4338] <=  8'h00;      memory[4339] <=  8'h00;      memory[4340] <=  8'h00;      memory[4341] <=  8'h00;      memory[4342] <=  8'h00;      memory[4343] <=  8'h00;      memory[4344] <=  8'h00;      memory[4345] <=  8'h00;      memory[4346] <=  8'h00;      memory[4347] <=  8'h00;      memory[4348] <=  8'h00;      memory[4349] <=  8'h00;      memory[4350] <=  8'h00;      memory[4351] <=  8'h00;      memory[4352] <=  8'h00;      memory[4353] <=  8'h00;      memory[4354] <=  8'h00;      memory[4355] <=  8'h00;      memory[4356] <=  8'h00;      memory[4357] <=  8'h00;      memory[4358] <=  8'h00;      memory[4359] <=  8'h00;      memory[4360] <=  8'h00;      memory[4361] <=  8'h00;      memory[4362] <=  8'h00;      memory[4363] <=  8'h00;      memory[4364] <=  8'h00;      memory[4365] <=  8'h00;      memory[4366] <=  8'h00;      memory[4367] <=  8'h00;      memory[4368] <=  8'h00;      memory[4369] <=  8'h00;      memory[4370] <=  8'h00;      memory[4371] <=  8'h00;      memory[4372] <=  8'h00;      memory[4373] <=  8'h00;      memory[4374] <=  8'h00;      memory[4375] <=  8'h00;      memory[4376] <=  8'h00;      memory[4377] <=  8'h00;      memory[4378] <=  8'h00;      memory[4379] <=  8'h00;      memory[4380] <=  8'h00;      memory[4381] <=  8'h00;      memory[4382] <=  8'h00;      memory[4383] <=  8'h00;      memory[4384] <=  8'h00;      memory[4385] <=  8'h00;      memory[4386] <=  8'h00;      memory[4387] <=  8'h00;      memory[4388] <=  8'h00;      memory[4389] <=  8'h00;      memory[4390] <=  8'h00;      memory[4391] <=  8'h00;      memory[4392] <=  8'h00;      memory[4393] <=  8'h00;      memory[4394] <=  8'h00;      memory[4395] <=  8'h00;      memory[4396] <=  8'h00;      memory[4397] <=  8'h00;      memory[4398] <=  8'h00;      memory[4399] <=  8'h00;      memory[4400] <=  8'h00;      memory[4401] <=  8'h00;      memory[4402] <=  8'h00;      memory[4403] <=  8'h00;      memory[4404] <=  8'h00;      memory[4405] <=  8'h00;      memory[4406] <=  8'h00;      memory[4407] <=  8'h00;      memory[4408] <=  8'h00;      memory[4409] <=  8'h00;      memory[4410] <=  8'h00;      memory[4411] <=  8'h00;      memory[4412] <=  8'h00;      memory[4413] <=  8'h00;      memory[4414] <=  8'h00;      memory[4415] <=  8'h00;      memory[4416] <=  8'h00;      memory[4417] <=  8'h00;      memory[4418] <=  8'h00;      memory[4419] <=  8'h00;      memory[4420] <=  8'h00;      memory[4421] <=  8'h00;      memory[4422] <=  8'h00;      memory[4423] <=  8'h00;      memory[4424] <=  8'h00;      memory[4425] <=  8'h00;      memory[4426] <=  8'h00;      memory[4427] <=  8'h00;      memory[4428] <=  8'h00;      memory[4429] <=  8'h00;      memory[4430] <=  8'h00;      memory[4431] <=  8'h00;      memory[4432] <=  8'h00;      memory[4433] <=  8'h00;      memory[4434] <=  8'h00;      memory[4435] <=  8'h00;      memory[4436] <=  8'h00;      memory[4437] <=  8'h00;      memory[4438] <=  8'h00;      memory[4439] <=  8'h00;      memory[4440] <=  8'h00;      memory[4441] <=  8'h00;      memory[4442] <=  8'h00;      memory[4443] <=  8'h00;      memory[4444] <=  8'h00;      memory[4445] <=  8'h00;      memory[4446] <=  8'h00;      memory[4447] <=  8'h00;      memory[4448] <=  8'h00;      memory[4449] <=  8'h00;      memory[4450] <=  8'h00;      memory[4451] <=  8'h00;      memory[4452] <=  8'h00;      memory[4453] <=  8'h00;      memory[4454] <=  8'h00;      memory[4455] <=  8'h00;      memory[4456] <=  8'h00;      memory[4457] <=  8'h00;      memory[4458] <=  8'h00;      memory[4459] <=  8'h00;      memory[4460] <=  8'h00;      memory[4461] <=  8'h00;      memory[4462] <=  8'h00;      memory[4463] <=  8'h00;      memory[4464] <=  8'h00;      memory[4465] <=  8'h00;      memory[4466] <=  8'h00;      memory[4467] <=  8'h00;      memory[4468] <=  8'h00;      memory[4469] <=  8'h00;      memory[4470] <=  8'h00;      memory[4471] <=  8'h00;      memory[4472] <=  8'h00;      memory[4473] <=  8'h00;      memory[4474] <=  8'h00;      memory[4475] <=  8'h00;      memory[4476] <=  8'h00;      memory[4477] <=  8'h00;      memory[4478] <=  8'h00;      memory[4479] <=  8'h00;      memory[4480] <=  8'h00;      memory[4481] <=  8'h00;      memory[4482] <=  8'h00;      memory[4483] <=  8'h00;      memory[4484] <=  8'h00;      memory[4485] <=  8'h00;      memory[4486] <=  8'h00;      memory[4487] <=  8'h00;      memory[4488] <=  8'h00;      memory[4489] <=  8'h00;      memory[4490] <=  8'h00;      memory[4491] <=  8'h00;      memory[4492] <=  8'h00;      memory[4493] <=  8'h00;      memory[4494] <=  8'h00;      memory[4495] <=  8'h00;      memory[4496] <=  8'h00;      memory[4497] <=  8'h00;      memory[4498] <=  8'h00;      memory[4499] <=  8'h00;      memory[4500] <=  8'h00;      memory[4501] <=  8'h00;      memory[4502] <=  8'h00;      memory[4503] <=  8'h00;      memory[4504] <=  8'h00;      memory[4505] <=  8'h00;      memory[4506] <=  8'h00;      memory[4507] <=  8'h00;      memory[4508] <=  8'h00;      memory[4509] <=  8'h00;      memory[4510] <=  8'h00;      memory[4511] <=  8'h00;      memory[4512] <=  8'h00;      memory[4513] <=  8'h00;      memory[4514] <=  8'h00;      memory[4515] <=  8'h00;      memory[4516] <=  8'h00;      memory[4517] <=  8'h00;      memory[4518] <=  8'h00;      memory[4519] <=  8'h00;      memory[4520] <=  8'h00;      memory[4521] <=  8'h00;      memory[4522] <=  8'h00;      memory[4523] <=  8'h00;      memory[4524] <=  8'h00;      memory[4525] <=  8'h00;      memory[4526] <=  8'h00;      memory[4527] <=  8'h00;      memory[4528] <=  8'h00;      memory[4529] <=  8'h00;      memory[4530] <=  8'h00;      memory[4531] <=  8'h00;      memory[4532] <=  8'h00;      memory[4533] <=  8'h00;      memory[4534] <=  8'h00;      memory[4535] <=  8'h00;      memory[4536] <=  8'h00;      memory[4537] <=  8'h00;      memory[4538] <=  8'h00;      memory[4539] <=  8'h00;      memory[4540] <=  8'h00;      memory[4541] <=  8'h00;      memory[4542] <=  8'h00;      memory[4543] <=  8'h00;      memory[4544] <=  8'h00;      memory[4545] <=  8'h00;      memory[4546] <=  8'h00;      memory[4547] <=  8'h00;      memory[4548] <=  8'h00;      memory[4549] <=  8'h00;      memory[4550] <=  8'h00;      memory[4551] <=  8'h00;      memory[4552] <=  8'h00;      memory[4553] <=  8'h00;      memory[4554] <=  8'h00;      memory[4555] <=  8'h00;      memory[4556] <=  8'h00;      memory[4557] <=  8'h00;      memory[4558] <=  8'h00;      memory[4559] <=  8'h00;      memory[4560] <=  8'h00;      memory[4561] <=  8'h00;      memory[4562] <=  8'h00;      memory[4563] <=  8'h00;      memory[4564] <=  8'h00;      memory[4565] <=  8'h00;      memory[4566] <=  8'h00;      memory[4567] <=  8'h00;      memory[4568] <=  8'h00;      memory[4569] <=  8'h00;      memory[4570] <=  8'h00;      memory[4571] <=  8'h00;      memory[4572] <=  8'h00;      memory[4573] <=  8'h00;      memory[4574] <=  8'h00;      memory[4575] <=  8'h00;      memory[4576] <=  8'h00;      memory[4577] <=  8'h00;      memory[4578] <=  8'h00;      memory[4579] <=  8'h00;      memory[4580] <=  8'h00;      memory[4581] <=  8'h00;      memory[4582] <=  8'h00;      memory[4583] <=  8'h00;      memory[4584] <=  8'h00;      memory[4585] <=  8'h00;      memory[4586] <=  8'h00;      memory[4587] <=  8'h00;      memory[4588] <=  8'h00;      memory[4589] <=  8'h00;      memory[4590] <=  8'h00;      memory[4591] <=  8'h00;      memory[4592] <=  8'h00;      memory[4593] <=  8'h00;      memory[4594] <=  8'h00;      memory[4595] <=  8'h00;      memory[4596] <=  8'h00;      memory[4597] <=  8'h00;      memory[4598] <=  8'h00;      memory[4599] <=  8'h00;      memory[4600] <=  8'h00;      memory[4601] <=  8'h00;      memory[4602] <=  8'h00;      memory[4603] <=  8'h00;      memory[4604] <=  8'h00;      memory[4605] <=  8'h00;      memory[4606] <=  8'h00;      memory[4607] <=  8'h00;      memory[4608] <=  8'h00;      memory[4609] <=  8'h00;      memory[4610] <=  8'h00;      memory[4611] <=  8'h00;      memory[4612] <=  8'h00;      memory[4613] <=  8'h00;      memory[4614] <=  8'h00;      memory[4615] <=  8'h00;      memory[4616] <=  8'h00;      memory[4617] <=  8'h00;      memory[4618] <=  8'h00;      memory[4619] <=  8'h00;      memory[4620] <=  8'h00;      memory[4621] <=  8'h00;      memory[4622] <=  8'h00;      memory[4623] <=  8'h00;      memory[4624] <=  8'h00;      memory[4625] <=  8'h00;      memory[4626] <=  8'h00;      memory[4627] <=  8'h00;      memory[4628] <=  8'h00;      memory[4629] <=  8'h00;      memory[4630] <=  8'h00;      memory[4631] <=  8'h00;      memory[4632] <=  8'h00;      memory[4633] <=  8'h00;      memory[4634] <=  8'h00;      memory[4635] <=  8'h00;      memory[4636] <=  8'h00;      memory[4637] <=  8'h00;      memory[4638] <=  8'h00;      memory[4639] <=  8'h00;      memory[4640] <=  8'h00;      memory[4641] <=  8'h00;      memory[4642] <=  8'h00;      memory[4643] <=  8'h00;      memory[4644] <=  8'h00;      memory[4645] <=  8'h00;      memory[4646] <=  8'h00;      memory[4647] <=  8'h00;      memory[4648] <=  8'h00;      memory[4649] <=  8'h00;      memory[4650] <=  8'h00;      memory[4651] <=  8'h00;      memory[4652] <=  8'h00;      memory[4653] <=  8'h00;      memory[4654] <=  8'h00;      memory[4655] <=  8'h00;      memory[4656] <=  8'h00;      memory[4657] <=  8'h00;      memory[4658] <=  8'h00;      memory[4659] <=  8'h00;      memory[4660] <=  8'h00;      memory[4661] <=  8'h00;      memory[4662] <=  8'h00;      memory[4663] <=  8'h00;      memory[4664] <=  8'h00;      memory[4665] <=  8'h00;      memory[4666] <=  8'h00;      memory[4667] <=  8'h00;      memory[4668] <=  8'h00;      memory[4669] <=  8'h00;      memory[4670] <=  8'h00;      memory[4671] <=  8'h00;      memory[4672] <=  8'h00;      memory[4673] <=  8'h00;      memory[4674] <=  8'h00;      memory[4675] <=  8'h00;      memory[4676] <=  8'h00;      memory[4677] <=  8'h00;      memory[4678] <=  8'h00;      memory[4679] <=  8'h00;      memory[4680] <=  8'h00;      memory[4681] <=  8'h00;      memory[4682] <=  8'h00;      memory[4683] <=  8'h00;      memory[4684] <=  8'h00;      memory[4685] <=  8'h00;      memory[4686] <=  8'h00;      memory[4687] <=  8'h00;      memory[4688] <=  8'h00;      memory[4689] <=  8'h00;      memory[4690] <=  8'h00;      memory[4691] <=  8'h00;      memory[4692] <=  8'h00;      memory[4693] <=  8'h00;      memory[4694] <=  8'h00;      memory[4695] <=  8'h00;      memory[4696] <=  8'h00;      memory[4697] <=  8'h00;      memory[4698] <=  8'h00;      memory[4699] <=  8'h00;      memory[4700] <=  8'h00;      memory[4701] <=  8'h00;      memory[4702] <=  8'h00;      memory[4703] <=  8'h00;      memory[4704] <=  8'h00;      memory[4705] <=  8'h00;      memory[4706] <=  8'h00;      memory[4707] <=  8'h00;      memory[4708] <=  8'h00;      memory[4709] <=  8'h00;      memory[4710] <=  8'h00;      memory[4711] <=  8'h00;      memory[4712] <=  8'h00;      memory[4713] <=  8'h00;      memory[4714] <=  8'h00;      memory[4715] <=  8'h00;      memory[4716] <=  8'h00;      memory[4717] <=  8'h00;      memory[4718] <=  8'h00;      memory[4719] <=  8'h00;      memory[4720] <=  8'h00;      memory[4721] <=  8'h00;      memory[4722] <=  8'h00;      memory[4723] <=  8'h00;      memory[4724] <=  8'h00;      memory[4725] <=  8'h00;      memory[4726] <=  8'h00;      memory[4727] <=  8'h00;      memory[4728] <=  8'h00;      memory[4729] <=  8'h00;      memory[4730] <=  8'h00;      memory[4731] <=  8'h00;      memory[4732] <=  8'h00;      memory[4733] <=  8'h00;      memory[4734] <=  8'h00;      memory[4735] <=  8'h00;      memory[4736] <=  8'h00;      memory[4737] <=  8'h00;      memory[4738] <=  8'h00;      memory[4739] <=  8'h00;      memory[4740] <=  8'h00;      memory[4741] <=  8'h00;      memory[4742] <=  8'h00;      memory[4743] <=  8'h00;      memory[4744] <=  8'h00;      memory[4745] <=  8'h00;      memory[4746] <=  8'h00;      memory[4747] <=  8'h00;      memory[4748] <=  8'h00;      memory[4749] <=  8'h00;      memory[4750] <=  8'h00;      memory[4751] <=  8'h00;      memory[4752] <=  8'h00;      memory[4753] <=  8'h00;      memory[4754] <=  8'h00;      memory[4755] <=  8'h00;      memory[4756] <=  8'h00;      memory[4757] <=  8'h00;      memory[4758] <=  8'h00;      memory[4759] <=  8'h00;      memory[4760] <=  8'h00;      memory[4761] <=  8'h00;      memory[4762] <=  8'h00;      memory[4763] <=  8'h00;      memory[4764] <=  8'h00;      memory[4765] <=  8'h00;      memory[4766] <=  8'h00;      memory[4767] <=  8'h00;      memory[4768] <=  8'h00;      memory[4769] <=  8'h00;      memory[4770] <=  8'h00;      memory[4771] <=  8'h00;      memory[4772] <=  8'h00;      memory[4773] <=  8'h00;      memory[4774] <=  8'h00;      memory[4775] <=  8'h00;      memory[4776] <=  8'h00;      memory[4777] <=  8'h00;      memory[4778] <=  8'h00;      memory[4779] <=  8'h00;      memory[4780] <=  8'h00;      memory[4781] <=  8'h00;      memory[4782] <=  8'h00;      memory[4783] <=  8'h00;      memory[4784] <=  8'h00;      memory[4785] <=  8'h00;      memory[4786] <=  8'h00;      memory[4787] <=  8'h00;      memory[4788] <=  8'h00;      memory[4789] <=  8'h00;      memory[4790] <=  8'h00;      memory[4791] <=  8'h00;      memory[4792] <=  8'h00;      memory[4793] <=  8'h00;      memory[4794] <=  8'h00;      memory[4795] <=  8'h00;      memory[4796] <=  8'h00;      memory[4797] <=  8'h00;      memory[4798] <=  8'h00;      memory[4799] <=  8'h00;      memory[4800] <=  8'h00;      memory[4801] <=  8'h00;      memory[4802] <=  8'h00;      memory[4803] <=  8'h00;      memory[4804] <=  8'h00;      memory[4805] <=  8'h00;      memory[4806] <=  8'h00;      memory[4807] <=  8'h00;      memory[4808] <=  8'h00;      memory[4809] <=  8'h00;      memory[4810] <=  8'h00;      memory[4811] <=  8'h00;      memory[4812] <=  8'h00;      memory[4813] <=  8'h00;      memory[4814] <=  8'h00;      memory[4815] <=  8'h00;      memory[4816] <=  8'h00;      memory[4817] <=  8'h00;      memory[4818] <=  8'h00;      memory[4819] <=  8'h00;      memory[4820] <=  8'h00;      memory[4821] <=  8'h00;      memory[4822] <=  8'h00;      memory[4823] <=  8'h00;      memory[4824] <=  8'h00;      memory[4825] <=  8'h00;      memory[4826] <=  8'h00;      memory[4827] <=  8'h00;      memory[4828] <=  8'h00;      memory[4829] <=  8'h00;      memory[4830] <=  8'h00;      memory[4831] <=  8'h00;      memory[4832] <=  8'h00;      memory[4833] <=  8'h00;      memory[4834] <=  8'h00;      memory[4835] <=  8'h00;      memory[4836] <=  8'h00;      memory[4837] <=  8'h00;      memory[4838] <=  8'h00;      memory[4839] <=  8'h00;      memory[4840] <=  8'h00;      memory[4841] <=  8'h00;      memory[4842] <=  8'h00;      memory[4843] <=  8'h00;      memory[4844] <=  8'h00;      memory[4845] <=  8'h00;      memory[4846] <=  8'h00;      memory[4847] <=  8'h00;      memory[4848] <=  8'h00;      memory[4849] <=  8'h00;      memory[4850] <=  8'h00;      memory[4851] <=  8'h00;      memory[4852] <=  8'h00;      memory[4853] <=  8'h00;      memory[4854] <=  8'h00;      memory[4855] <=  8'h00;      memory[4856] <=  8'h00;      memory[4857] <=  8'h00;      memory[4858] <=  8'h00;      memory[4859] <=  8'h00;      memory[4860] <=  8'h00;      memory[4861] <=  8'h00;      memory[4862] <=  8'h00;      memory[4863] <=  8'h00;      memory[4864] <=  8'h00;      memory[4865] <=  8'h00;      memory[4866] <=  8'h00;      memory[4867] <=  8'h00;      memory[4868] <=  8'h00;      memory[4869] <=  8'h00;      memory[4870] <=  8'h00;      memory[4871] <=  8'h00;      memory[4872] <=  8'h00;      memory[4873] <=  8'h00;      memory[4874] <=  8'h00;      memory[4875] <=  8'h00;      memory[4876] <=  8'h00;      memory[4877] <=  8'h00;      memory[4878] <=  8'h00;      memory[4879] <=  8'h00;      memory[4880] <=  8'h00;      memory[4881] <=  8'h00;      memory[4882] <=  8'h00;      memory[4883] <=  8'h00;      memory[4884] <=  8'h00;      memory[4885] <=  8'h00;      memory[4886] <=  8'h00;      memory[4887] <=  8'h00;      memory[4888] <=  8'h00;      memory[4889] <=  8'h00;      memory[4890] <=  8'h00;      memory[4891] <=  8'h00;      memory[4892] <=  8'h00;      memory[4893] <=  8'h00;      memory[4894] <=  8'h00;      memory[4895] <=  8'h00;      memory[4896] <=  8'h00;      memory[4897] <=  8'h00;      memory[4898] <=  8'h00;      memory[4899] <=  8'h00;      memory[4900] <=  8'h00;      memory[4901] <=  8'h00;      memory[4902] <=  8'h00;      memory[4903] <=  8'h00;      memory[4904] <=  8'h00;      memory[4905] <=  8'h00;      memory[4906] <=  8'h00;      memory[4907] <=  8'h00;      memory[4908] <=  8'h00;      memory[4909] <=  8'h00;      memory[4910] <=  8'h00;      memory[4911] <=  8'h00;      memory[4912] <=  8'h00;      memory[4913] <=  8'h00;      memory[4914] <=  8'h00;      memory[4915] <=  8'h00;      memory[4916] <=  8'h00;      memory[4917] <=  8'h00;      memory[4918] <=  8'h00;      memory[4919] <=  8'h00;      memory[4920] <=  8'h00;      memory[4921] <=  8'h00;      memory[4922] <=  8'h00;      memory[4923] <=  8'h00;      memory[4924] <=  8'h00;      memory[4925] <=  8'h00;      memory[4926] <=  8'h00;      memory[4927] <=  8'h00;      memory[4928] <=  8'h00;      memory[4929] <=  8'h00;      memory[4930] <=  8'h00;      memory[4931] <=  8'h00;      memory[4932] <=  8'h00;      memory[4933] <=  8'h00;      memory[4934] <=  8'h00;      memory[4935] <=  8'h00;      memory[4936] <=  8'h00;      memory[4937] <=  8'h00;      memory[4938] <=  8'h00;      memory[4939] <=  8'h00;      memory[4940] <=  8'h00;      memory[4941] <=  8'h00;      memory[4942] <=  8'h00;      memory[4943] <=  8'h00;      memory[4944] <=  8'h00;      memory[4945] <=  8'h00;      memory[4946] <=  8'h00;      memory[4947] <=  8'h00;      memory[4948] <=  8'h00;      memory[4949] <=  8'h00;      memory[4950] <=  8'h00;      memory[4951] <=  8'h00;      memory[4952] <=  8'h00;      memory[4953] <=  8'h00;      memory[4954] <=  8'h00;      memory[4955] <=  8'h00;      memory[4956] <=  8'h00;      memory[4957] <=  8'h00;      memory[4958] <=  8'h00;      memory[4959] <=  8'h00;      memory[4960] <=  8'h00;      memory[4961] <=  8'h00;      memory[4962] <=  8'h00;      memory[4963] <=  8'h00;      memory[4964] <=  8'h00;      memory[4965] <=  8'h00;      memory[4966] <=  8'h00;      memory[4967] <=  8'h00;      memory[4968] <=  8'h00;      memory[4969] <=  8'h00;      memory[4970] <=  8'h00;      memory[4971] <=  8'h00;      memory[4972] <=  8'h00;      memory[4973] <=  8'h00;      memory[4974] <=  8'h00;      memory[4975] <=  8'h00;      memory[4976] <=  8'h00;      memory[4977] <=  8'h00;      memory[4978] <=  8'h00;      memory[4979] <=  8'h00;      memory[4980] <=  8'h00;      memory[4981] <=  8'h00;      memory[4982] <=  8'h00;      memory[4983] <=  8'h00;      memory[4984] <=  8'h00;      memory[4985] <=  8'h00;      memory[4986] <=  8'h00;      memory[4987] <=  8'h00;      memory[4988] <=  8'h00;      memory[4989] <=  8'h00;      memory[4990] <=  8'h00;      memory[4991] <=  8'h00;      memory[4992] <=  8'h00;      memory[4993] <=  8'h00;      memory[4994] <=  8'h00;      memory[4995] <=  8'h00;      memory[4996] <=  8'h00;      memory[4997] <=  8'h00;      memory[4998] <=  8'h00;      memory[4999] <=  8'h00;      memory[5000] <=  8'h00;      memory[5001] <=  8'h00;      memory[5002] <=  8'h00;      memory[5003] <=  8'h00;      memory[5004] <=  8'h00;      memory[5005] <=  8'h00;      memory[5006] <=  8'h00;      memory[5007] <=  8'h00;      memory[5008] <=  8'h00;      memory[5009] <=  8'h00;      memory[5010] <=  8'h00;      memory[5011] <=  8'h00;      memory[5012] <=  8'h00;      memory[5013] <=  8'h00;      memory[5014] <=  8'h00;      memory[5015] <=  8'h00;      memory[5016] <=  8'h00;      memory[5017] <=  8'h00;      memory[5018] <=  8'h00;      memory[5019] <=  8'h00;      memory[5020] <=  8'h00;      memory[5021] <=  8'h00;      memory[5022] <=  8'h00;      memory[5023] <=  8'h00;      memory[5024] <=  8'h00;      memory[5025] <=  8'h00;      memory[5026] <=  8'h00;      memory[5027] <=  8'h00;      memory[5028] <=  8'h00;      memory[5029] <=  8'h00;      memory[5030] <=  8'h00;      memory[5031] <=  8'h00;      memory[5032] <=  8'h00;      memory[5033] <=  8'h00;      memory[5034] <=  8'h00;      memory[5035] <=  8'h00;      memory[5036] <=  8'h00;      memory[5037] <=  8'h00;      memory[5038] <=  8'h00;      memory[5039] <=  8'h00;      memory[5040] <=  8'h00;      memory[5041] <=  8'h00;      memory[5042] <=  8'h00;      memory[5043] <=  8'h00;      memory[5044] <=  8'h00;      memory[5045] <=  8'h00;      memory[5046] <=  8'h00;      memory[5047] <=  8'h00;      memory[5048] <=  8'h00;      memory[5049] <=  8'h00;      memory[5050] <=  8'h00;      memory[5051] <=  8'h00;      memory[5052] <=  8'h00;      memory[5053] <=  8'h00;      memory[5054] <=  8'h00;      memory[5055] <=  8'h00;      memory[5056] <=  8'h00;      memory[5057] <=  8'h00;      memory[5058] <=  8'h00;      memory[5059] <=  8'h00;      memory[5060] <=  8'h00;      memory[5061] <=  8'h00;      memory[5062] <=  8'h00;      memory[5063] <=  8'h00;      memory[5064] <=  8'h00;      memory[5065] <=  8'h00;      memory[5066] <=  8'h00;      memory[5067] <=  8'h00;      memory[5068] <=  8'h00;      memory[5069] <=  8'h00;      memory[5070] <=  8'h00;      memory[5071] <=  8'h00;      memory[5072] <=  8'h00;      memory[5073] <=  8'h00;      memory[5074] <=  8'h00;      memory[5075] <=  8'h00;      memory[5076] <=  8'h00;      memory[5077] <=  8'h00;      memory[5078] <=  8'h00;      memory[5079] <=  8'h00;      memory[5080] <=  8'h00;      memory[5081] <=  8'h00;      memory[5082] <=  8'h00;      memory[5083] <=  8'h00;      memory[5084] <=  8'h00;      memory[5085] <=  8'h00;      memory[5086] <=  8'h00;      memory[5087] <=  8'h00;      memory[5088] <=  8'h00;      memory[5089] <=  8'h00;      memory[5090] <=  8'h00;      memory[5091] <=  8'h00;      memory[5092] <=  8'h00;      memory[5093] <=  8'h00;      memory[5094] <=  8'h00;      memory[5095] <=  8'h00;      memory[5096] <=  8'h00;      memory[5097] <=  8'h00;      memory[5098] <=  8'h00;      memory[5099] <=  8'h00;      memory[5100] <=  8'h00;      memory[5101] <=  8'h00;      memory[5102] <=  8'h00;      memory[5103] <=  8'h00;      memory[5104] <=  8'h00;      memory[5105] <=  8'h00;      memory[5106] <=  8'h00;      memory[5107] <=  8'h00;      memory[5108] <=  8'h00;      memory[5109] <=  8'h00;      memory[5110] <=  8'h00;      memory[5111] <=  8'h00;      memory[5112] <=  8'h00;      memory[5113] <=  8'h00;      memory[5114] <=  8'h00;      memory[5115] <=  8'h00;      memory[5116] <=  8'h00;      memory[5117] <=  8'h00;      memory[5118] <=  8'h00;      memory[5119] <=  8'h00;      memory[5120] <=  8'h00;      memory[5121] <=  8'h00;      memory[5122] <=  8'h00;      memory[5123] <=  8'h00;      memory[5124] <=  8'h00;      memory[5125] <=  8'h00;      memory[5126] <=  8'h00;      memory[5127] <=  8'h00;      memory[5128] <=  8'h00;      memory[5129] <=  8'h00;      memory[5130] <=  8'h00;      memory[5131] <=  8'h00;      memory[5132] <=  8'h00;      memory[5133] <=  8'h00;      memory[5134] <=  8'h00;      memory[5135] <=  8'h00;      memory[5136] <=  8'h00;      memory[5137] <=  8'h00;      memory[5138] <=  8'h00;      memory[5139] <=  8'h00;      memory[5140] <=  8'h00;      memory[5141] <=  8'h00;      memory[5142] <=  8'h00;      memory[5143] <=  8'h00;      memory[5144] <=  8'h00;      memory[5145] <=  8'h00;      memory[5146] <=  8'h00;      memory[5147] <=  8'h00;      memory[5148] <=  8'h00;      memory[5149] <=  8'h00;      memory[5150] <=  8'h00;      memory[5151] <=  8'h00;      memory[5152] <=  8'h00;      memory[5153] <=  8'h00;      memory[5154] <=  8'h00;      memory[5155] <=  8'h00;      memory[5156] <=  8'h00;      memory[5157] <=  8'h00;      memory[5158] <=  8'h00;      memory[5159] <=  8'h00;      memory[5160] <=  8'h00;      memory[5161] <=  8'h00;      memory[5162] <=  8'h00;      memory[5163] <=  8'h00;      memory[5164] <=  8'h00;      memory[5165] <=  8'h00;      memory[5166] <=  8'h00;      memory[5167] <=  8'h00;      memory[5168] <=  8'h00;      memory[5169] <=  8'h00;      memory[5170] <=  8'h00;      memory[5171] <=  8'h00;      memory[5172] <=  8'h00;      memory[5173] <=  8'h00;      memory[5174] <=  8'h00;      memory[5175] <=  8'h00;      memory[5176] <=  8'h00;      memory[5177] <=  8'h00;      memory[5178] <=  8'h00;      memory[5179] <=  8'h00;      memory[5180] <=  8'h00;      memory[5181] <=  8'h00;      memory[5182] <=  8'h00;      memory[5183] <=  8'h00;      memory[5184] <=  8'h00;      memory[5185] <=  8'h00;      memory[5186] <=  8'h00;      memory[5187] <=  8'h00;      memory[5188] <=  8'h00;      memory[5189] <=  8'h00;      memory[5190] <=  8'h00;      memory[5191] <=  8'h00;      memory[5192] <=  8'h00;      memory[5193] <=  8'h00;      memory[5194] <=  8'h00;      memory[5195] <=  8'h00;      memory[5196] <=  8'h00;      memory[5197] <=  8'h00;      memory[5198] <=  8'h00;      memory[5199] <=  8'h00;      memory[5200] <=  8'h00;      memory[5201] <=  8'h00;      memory[5202] <=  8'h00;      memory[5203] <=  8'h00;      memory[5204] <=  8'h00;      memory[5205] <=  8'h00;      memory[5206] <=  8'h00;      memory[5207] <=  8'h00;      memory[5208] <=  8'h00;      memory[5209] <=  8'h00;      memory[5210] <=  8'h00;      memory[5211] <=  8'h00;      memory[5212] <=  8'h00;      memory[5213] <=  8'h00;      memory[5214] <=  8'h00;      memory[5215] <=  8'h00;      memory[5216] <=  8'h00;      memory[5217] <=  8'h00;      memory[5218] <=  8'h00;      memory[5219] <=  8'h00;      memory[5220] <=  8'h00;      memory[5221] <=  8'h00;      memory[5222] <=  8'h00;      memory[5223] <=  8'h00;      memory[5224] <=  8'h00;      memory[5225] <=  8'h00;      memory[5226] <=  8'h00;      memory[5227] <=  8'h00;      memory[5228] <=  8'h00;      memory[5229] <=  8'h00;      memory[5230] <=  8'h00;      memory[5231] <=  8'h00;      memory[5232] <=  8'h00;      memory[5233] <=  8'h00;      memory[5234] <=  8'h00;      memory[5235] <=  8'h00;      memory[5236] <=  8'h00;      memory[5237] <=  8'h00;      memory[5238] <=  8'h00;      memory[5239] <=  8'h00;      memory[5240] <=  8'h00;      memory[5241] <=  8'h00;      memory[5242] <=  8'h00;      memory[5243] <=  8'h00;      memory[5244] <=  8'h00;      memory[5245] <=  8'h00;      memory[5246] <=  8'h00;      memory[5247] <=  8'h00;      memory[5248] <=  8'h00;      memory[5249] <=  8'h00;      memory[5250] <=  8'h00;      memory[5251] <=  8'h00;      memory[5252] <=  8'h00;      memory[5253] <=  8'h00;      memory[5254] <=  8'h00;      memory[5255] <=  8'h00;      memory[5256] <=  8'h00;      memory[5257] <=  8'h00;      memory[5258] <=  8'h00;      memory[5259] <=  8'h00;      memory[5260] <=  8'h00;      memory[5261] <=  8'h00;      memory[5262] <=  8'h00;      memory[5263] <=  8'h00;      memory[5264] <=  8'h00;      memory[5265] <=  8'h00;      memory[5266] <=  8'h00;      memory[5267] <=  8'h00;      memory[5268] <=  8'h00;      memory[5269] <=  8'h00;      memory[5270] <=  8'h00;      memory[5271] <=  8'h00;      memory[5272] <=  8'h00;      memory[5273] <=  8'h00;      memory[5274] <=  8'h00;      memory[5275] <=  8'h00;      memory[5276] <=  8'h00;      memory[5277] <=  8'h00;      memory[5278] <=  8'h00;      memory[5279] <=  8'h00;      memory[5280] <=  8'h00;      memory[5281] <=  8'h00;      memory[5282] <=  8'h00;      memory[5283] <=  8'h00;      memory[5284] <=  8'h00;      memory[5285] <=  8'h00;      memory[5286] <=  8'h00;      memory[5287] <=  8'h00;      memory[5288] <=  8'h00;      memory[5289] <=  8'h00;      memory[5290] <=  8'h00;      memory[5291] <=  8'h00;      memory[5292] <=  8'h00;      memory[5293] <=  8'h00;      memory[5294] <=  8'h00;      memory[5295] <=  8'h00;      memory[5296] <=  8'h00;      memory[5297] <=  8'h00;      memory[5298] <=  8'h00;      memory[5299] <=  8'h00;      memory[5300] <=  8'h00;      memory[5301] <=  8'h00;      memory[5302] <=  8'h00;      memory[5303] <=  8'h00;      memory[5304] <=  8'h00;      memory[5305] <=  8'h00;      memory[5306] <=  8'h00;      memory[5307] <=  8'h00;      memory[5308] <=  8'h00;      memory[5309] <=  8'h00;      memory[5310] <=  8'h00;      memory[5311] <=  8'h00;      memory[5312] <=  8'h00;      memory[5313] <=  8'h00;      memory[5314] <=  8'h00;      memory[5315] <=  8'h00;      memory[5316] <=  8'h00;      memory[5317] <=  8'h00;      memory[5318] <=  8'h00;      memory[5319] <=  8'h00;      memory[5320] <=  8'h00;      memory[5321] <=  8'h00;      memory[5322] <=  8'h00;      memory[5323] <=  8'h00;      memory[5324] <=  8'h00;      memory[5325] <=  8'h00;      memory[5326] <=  8'h00;      memory[5327] <=  8'h00;      memory[5328] <=  8'h00;      memory[5329] <=  8'h00;      memory[5330] <=  8'h00;      memory[5331] <=  8'h00;      memory[5332] <=  8'h00;      memory[5333] <=  8'h00;      memory[5334] <=  8'h00;      memory[5335] <=  8'h00;      memory[5336] <=  8'h00;      memory[5337] <=  8'h00;      memory[5338] <=  8'h00;      memory[5339] <=  8'h00;      memory[5340] <=  8'h00;      memory[5341] <=  8'h00;      memory[5342] <=  8'h00;      memory[5343] <=  8'h00;      memory[5344] <=  8'h00;      memory[5345] <=  8'h00;      memory[5346] <=  8'h00;      memory[5347] <=  8'h00;      memory[5348] <=  8'h00;      memory[5349] <=  8'h00;      memory[5350] <=  8'h00;      memory[5351] <=  8'h00;      memory[5352] <=  8'h00;      memory[5353] <=  8'h00;      memory[5354] <=  8'h00;      memory[5355] <=  8'h00;      memory[5356] <=  8'h00;      memory[5357] <=  8'h00;      memory[5358] <=  8'h00;      memory[5359] <=  8'h00;      memory[5360] <=  8'h00;      memory[5361] <=  8'h00;      memory[5362] <=  8'h00;      memory[5363] <=  8'h00;      memory[5364] <=  8'h00;      memory[5365] <=  8'h00;      memory[5366] <=  8'h00;      memory[5367] <=  8'h00;      memory[5368] <=  8'h00;      memory[5369] <=  8'h00;      memory[5370] <=  8'h00;      memory[5371] <=  8'h00;      memory[5372] <=  8'h00;      memory[5373] <=  8'h00;      memory[5374] <=  8'h00;      memory[5375] <=  8'h00;      memory[5376] <=  8'h00;      memory[5377] <=  8'h00;      memory[5378] <=  8'h00;      memory[5379] <=  8'h00;      memory[5380] <=  8'h00;      memory[5381] <=  8'h00;      memory[5382] <=  8'h00;      memory[5383] <=  8'h00;      memory[5384] <=  8'h00;      memory[5385] <=  8'h00;      memory[5386] <=  8'h00;      memory[5387] <=  8'h00;      memory[5388] <=  8'h00;      memory[5389] <=  8'h00;      memory[5390] <=  8'h00;      memory[5391] <=  8'h00;      memory[5392] <=  8'h00;      memory[5393] <=  8'h00;      memory[5394] <=  8'h00;      memory[5395] <=  8'h00;      memory[5396] <=  8'h00;      memory[5397] <=  8'h00;      memory[5398] <=  8'h00;      memory[5399] <=  8'h00;      memory[5400] <=  8'h00;      memory[5401] <=  8'h00;      memory[5402] <=  8'h00;      memory[5403] <=  8'h00;      memory[5404] <=  8'h00;      memory[5405] <=  8'h00;      memory[5406] <=  8'h00;      memory[5407] <=  8'h00;      memory[5408] <=  8'h00;      memory[5409] <=  8'h00;      memory[5410] <=  8'h00;      memory[5411] <=  8'h00;      memory[5412] <=  8'h00;      memory[5413] <=  8'h00;      memory[5414] <=  8'h00;      memory[5415] <=  8'h00;      memory[5416] <=  8'h00;      memory[5417] <=  8'h00;      memory[5418] <=  8'h00;      memory[5419] <=  8'h00;      memory[5420] <=  8'h00;      memory[5421] <=  8'h00;      memory[5422] <=  8'h00;      memory[5423] <=  8'h00;      memory[5424] <=  8'h00;      memory[5425] <=  8'h00;      memory[5426] <=  8'h00;      memory[5427] <=  8'h00;      memory[5428] <=  8'h00;      memory[5429] <=  8'h00;      memory[5430] <=  8'h00;      memory[5431] <=  8'h00;      memory[5432] <=  8'h00;      memory[5433] <=  8'h00;      memory[5434] <=  8'h00;      memory[5435] <=  8'h00;      memory[5436] <=  8'h00;      memory[5437] <=  8'h00;      memory[5438] <=  8'h00;      memory[5439] <=  8'h00;      memory[5440] <=  8'h00;      memory[5441] <=  8'h00;      memory[5442] <=  8'h00;      memory[5443] <=  8'h00;      memory[5444] <=  8'h00;      memory[5445] <=  8'h00;      memory[5446] <=  8'h00;      memory[5447] <=  8'h00;      memory[5448] <=  8'h00;      memory[5449] <=  8'h00;      memory[5450] <=  8'h00;      memory[5451] <=  8'h00;      memory[5452] <=  8'h00;      memory[5453] <=  8'h00;      memory[5454] <=  8'h00;      memory[5455] <=  8'h00;      memory[5456] <=  8'h00;      memory[5457] <=  8'h00;      memory[5458] <=  8'h00;      memory[5459] <=  8'h00;      memory[5460] <=  8'h00;      memory[5461] <=  8'h00;      memory[5462] <=  8'h00;      memory[5463] <=  8'h00;      memory[5464] <=  8'h00;      memory[5465] <=  8'h00;      memory[5466] <=  8'h00;      memory[5467] <=  8'h00;      memory[5468] <=  8'h00;      memory[5469] <=  8'h00;      memory[5470] <=  8'h00;      memory[5471] <=  8'h00;      memory[5472] <=  8'h00;      memory[5473] <=  8'h00;      memory[5474] <=  8'h00;      memory[5475] <=  8'h00;      memory[5476] <=  8'h00;      memory[5477] <=  8'h00;      memory[5478] <=  8'h00;      memory[5479] <=  8'h00;      memory[5480] <=  8'h00;      memory[5481] <=  8'h00;      memory[5482] <=  8'h00;      memory[5483] <=  8'h00;      memory[5484] <=  8'h00;      memory[5485] <=  8'h00;      memory[5486] <=  8'h00;      memory[5487] <=  8'h00;      memory[5488] <=  8'h00;      memory[5489] <=  8'h00;      memory[5490] <=  8'h00;      memory[5491] <=  8'h00;      memory[5492] <=  8'h00;      memory[5493] <=  8'h00;      memory[5494] <=  8'h00;      memory[5495] <=  8'h00;      memory[5496] <=  8'h00;      memory[5497] <=  8'h00;      memory[5498] <=  8'h00;      memory[5499] <=  8'h00;      memory[5500] <=  8'h00;      memory[5501] <=  8'h00;      memory[5502] <=  8'h00;      memory[5503] <=  8'h00;      memory[5504] <=  8'h00;      memory[5505] <=  8'h00;      memory[5506] <=  8'h00;      memory[5507] <=  8'h00;      memory[5508] <=  8'h00;      memory[5509] <=  8'h00;      memory[5510] <=  8'h00;      memory[5511] <=  8'h00;      memory[5512] <=  8'h00;      memory[5513] <=  8'h00;      memory[5514] <=  8'h00;      memory[5515] <=  8'h00;      memory[5516] <=  8'h00;      memory[5517] <=  8'h00;      memory[5518] <=  8'h00;      memory[5519] <=  8'h00;      memory[5520] <=  8'h00;      memory[5521] <=  8'h00;      memory[5522] <=  8'h00;      memory[5523] <=  8'h00;      memory[5524] <=  8'h00;      memory[5525] <=  8'h00;      memory[5526] <=  8'h00;      memory[5527] <=  8'h00;      memory[5528] <=  8'h00;      memory[5529] <=  8'h00;      memory[5530] <=  8'h00;      memory[5531] <=  8'h00;      memory[5532] <=  8'h00;      memory[5533] <=  8'h00;      memory[5534] <=  8'h00;      memory[5535] <=  8'h00;      memory[5536] <=  8'h00;      memory[5537] <=  8'h00;      memory[5538] <=  8'h00;      memory[5539] <=  8'h00;      memory[5540] <=  8'h00;      memory[5541] <=  8'h00;      memory[5542] <=  8'h00;      memory[5543] <=  8'h00;      memory[5544] <=  8'h00;      memory[5545] <=  8'h00;      memory[5546] <=  8'h00;      memory[5547] <=  8'h00;      memory[5548] <=  8'h00;      memory[5549] <=  8'h00;      memory[5550] <=  8'h00;      memory[5551] <=  8'h00;      memory[5552] <=  8'h00;      memory[5553] <=  8'h00;      memory[5554] <=  8'h00;      memory[5555] <=  8'h00;      memory[5556] <=  8'h00;      memory[5557] <=  8'h00;      memory[5558] <=  8'h00;      memory[5559] <=  8'h00;      memory[5560] <=  8'h00;      memory[5561] <=  8'h00;      memory[5562] <=  8'h00;      memory[5563] <=  8'h00;      memory[5564] <=  8'h00;      memory[5565] <=  8'h00;      memory[5566] <=  8'h00;      memory[5567] <=  8'h00;      memory[5568] <=  8'h00;      memory[5569] <=  8'h00;      memory[5570] <=  8'h00;      memory[5571] <=  8'h00;      memory[5572] <=  8'h00;      memory[5573] <=  8'h00;      memory[5574] <=  8'h00;      memory[5575] <=  8'h00;      memory[5576] <=  8'h00;      memory[5577] <=  8'h00;      memory[5578] <=  8'h00;      memory[5579] <=  8'h00;      memory[5580] <=  8'h00;      memory[5581] <=  8'h00;      memory[5582] <=  8'h00;      memory[5583] <=  8'h00;      memory[5584] <=  8'h00;      memory[5585] <=  8'h00;      memory[5586] <=  8'h00;      memory[5587] <=  8'h00;      memory[5588] <=  8'h00;      memory[5589] <=  8'h00;      memory[5590] <=  8'h00;      memory[5591] <=  8'h00;      memory[5592] <=  8'h00;      memory[5593] <=  8'h00;      memory[5594] <=  8'h00;      memory[5595] <=  8'h00;      memory[5596] <=  8'h00;      memory[5597] <=  8'h00;      memory[5598] <=  8'h00;      memory[5599] <=  8'h00;      memory[5600] <=  8'h00;      memory[5601] <=  8'h00;      memory[5602] <=  8'h00;      memory[5603] <=  8'h00;      memory[5604] <=  8'h00;      memory[5605] <=  8'h00;      memory[5606] <=  8'h00;      memory[5607] <=  8'h00;      memory[5608] <=  8'h00;      memory[5609] <=  8'h00;      memory[5610] <=  8'h00;      memory[5611] <=  8'h00;      memory[5612] <=  8'h00;      memory[5613] <=  8'h00;      memory[5614] <=  8'h00;      memory[5615] <=  8'h00;      memory[5616] <=  8'h00;      memory[5617] <=  8'h00;      memory[5618] <=  8'h00;      memory[5619] <=  8'h00;      memory[5620] <=  8'h00;      memory[5621] <=  8'h00;      memory[5622] <=  8'h00;      memory[5623] <=  8'h00;      memory[5624] <=  8'h00;      memory[5625] <=  8'h00;      memory[5626] <=  8'h00;      memory[5627] <=  8'h00;      memory[5628] <=  8'h00;      memory[5629] <=  8'h00;      memory[5630] <=  8'h00;      memory[5631] <=  8'h00;      memory[5632] <=  8'h00;      memory[5633] <=  8'h00;      memory[5634] <=  8'h00;      memory[5635] <=  8'h00;      memory[5636] <=  8'h00;      memory[5637] <=  8'h00;      memory[5638] <=  8'h00;      memory[5639] <=  8'h00;      memory[5640] <=  8'h00;      memory[5641] <=  8'h00;      memory[5642] <=  8'h00;      memory[5643] <=  8'h00;      memory[5644] <=  8'h00;      memory[5645] <=  8'h00;      memory[5646] <=  8'h00;      memory[5647] <=  8'h00;      memory[5648] <=  8'h00;      memory[5649] <=  8'h00;      memory[5650] <=  8'h00;      memory[5651] <=  8'h00;      memory[5652] <=  8'h00;      memory[5653] <=  8'h00;      memory[5654] <=  8'h00;      memory[5655] <=  8'h00;      memory[5656] <=  8'h00;      memory[5657] <=  8'h00;      memory[5658] <=  8'h00;      memory[5659] <=  8'h00;      memory[5660] <=  8'h00;      memory[5661] <=  8'h00;      memory[5662] <=  8'h00;      memory[5663] <=  8'h00;      memory[5664] <=  8'h00;      memory[5665] <=  8'h00;      memory[5666] <=  8'h00;      memory[5667] <=  8'h00;      memory[5668] <=  8'h00;      memory[5669] <=  8'h00;      memory[5670] <=  8'h00;      memory[5671] <=  8'h00;      memory[5672] <=  8'h00;      memory[5673] <=  8'h00;      memory[5674] <=  8'h00;      memory[5675] <=  8'h00;      memory[5676] <=  8'h00;      memory[5677] <=  8'h00;      memory[5678] <=  8'h00;      memory[5679] <=  8'h00;      memory[5680] <=  8'h00;      memory[5681] <=  8'h00;      memory[5682] <=  8'h00;      memory[5683] <=  8'h00;      memory[5684] <=  8'h00;      memory[5685] <=  8'h00;      memory[5686] <=  8'h00;      memory[5687] <=  8'h00;      memory[5688] <=  8'h00;      memory[5689] <=  8'h00;      memory[5690] <=  8'h00;      memory[5691] <=  8'h00;      memory[5692] <=  8'h00;      memory[5693] <=  8'h00;      memory[5694] <=  8'h00;      memory[5695] <=  8'h00;      memory[5696] <=  8'h00;      memory[5697] <=  8'h00;      memory[5698] <=  8'h00;      memory[5699] <=  8'h00;      memory[5700] <=  8'h00;      memory[5701] <=  8'h00;      memory[5702] <=  8'h00;      memory[5703] <=  8'h00;      memory[5704] <=  8'h00;      memory[5705] <=  8'h00;      memory[5706] <=  8'h00;      memory[5707] <=  8'h00;      memory[5708] <=  8'h00;      memory[5709] <=  8'h00;      memory[5710] <=  8'h00;      memory[5711] <=  8'h00;      memory[5712] <=  8'h00;      memory[5713] <=  8'h00;      memory[5714] <=  8'h00;      memory[5715] <=  8'h00;      memory[5716] <=  8'h00;      memory[5717] <=  8'h00;      memory[5718] <=  8'h00;      memory[5719] <=  8'h00;      memory[5720] <=  8'h00;      memory[5721] <=  8'h00;      memory[5722] <=  8'h00;      memory[5723] <=  8'h00;      memory[5724] <=  8'h00;      memory[5725] <=  8'h00;      memory[5726] <=  8'h00;      memory[5727] <=  8'h00;      memory[5728] <=  8'h00;      memory[5729] <=  8'h00;      memory[5730] <=  8'h00;      memory[5731] <=  8'h00;      memory[5732] <=  8'h00;      memory[5733] <=  8'h00;      memory[5734] <=  8'h00;      memory[5735] <=  8'h00;      memory[5736] <=  8'h00;      memory[5737] <=  8'h00;      memory[5738] <=  8'h00;      memory[5739] <=  8'h00;      memory[5740] <=  8'h00;      memory[5741] <=  8'h00;      memory[5742] <=  8'h00;      memory[5743] <=  8'h00;      memory[5744] <=  8'h00;      memory[5745] <=  8'h00;      memory[5746] <=  8'h00;      memory[5747] <=  8'h00;      memory[5748] <=  8'h00;      memory[5749] <=  8'h00;      memory[5750] <=  8'h00;      memory[5751] <=  8'h00;      memory[5752] <=  8'h00;      memory[5753] <=  8'h00;      memory[5754] <=  8'h00;      memory[5755] <=  8'h00;      memory[5756] <=  8'h00;      memory[5757] <=  8'h00;      memory[5758] <=  8'h00;      memory[5759] <=  8'h00;      memory[5760] <=  8'h00;      memory[5761] <=  8'h00;      memory[5762] <=  8'h00;      memory[5763] <=  8'h00;      memory[5764] <=  8'h00;      memory[5765] <=  8'h00;      memory[5766] <=  8'h00;      memory[5767] <=  8'h00;      memory[5768] <=  8'h00;      memory[5769] <=  8'h00;      memory[5770] <=  8'h00;      memory[5771] <=  8'h00;      memory[5772] <=  8'h00;      memory[5773] <=  8'h00;      memory[5774] <=  8'h00;      memory[5775] <=  8'h00;      memory[5776] <=  8'h00;      memory[5777] <=  8'h00;      memory[5778] <=  8'h00;      memory[5779] <=  8'h00;      memory[5780] <=  8'h00;      memory[5781] <=  8'h00;      memory[5782] <=  8'h00;      memory[5783] <=  8'h00;      memory[5784] <=  8'h00;      memory[5785] <=  8'h00;      memory[5786] <=  8'h00;      memory[5787] <=  8'h00;      memory[5788] <=  8'h00;      memory[5789] <=  8'h00;      memory[5790] <=  8'h00;      memory[5791] <=  8'h00;      memory[5792] <=  8'h00;      memory[5793] <=  8'h00;      memory[5794] <=  8'h00;      memory[5795] <=  8'h00;      memory[5796] <=  8'h00;      memory[5797] <=  8'h00;      memory[5798] <=  8'h00;      memory[5799] <=  8'h00;      memory[5800] <=  8'h00;      memory[5801] <=  8'h00;      memory[5802] <=  8'h00;      memory[5803] <=  8'h00;      memory[5804] <=  8'h00;      memory[5805] <=  8'h00;      memory[5806] <=  8'h00;      memory[5807] <=  8'h00;      memory[5808] <=  8'h00;      memory[5809] <=  8'h00;      memory[5810] <=  8'h00;      memory[5811] <=  8'h00;      memory[5812] <=  8'h00;      memory[5813] <=  8'h00;      memory[5814] <=  8'h00;      memory[5815] <=  8'h00;      memory[5816] <=  8'h00;      memory[5817] <=  8'h00;      memory[5818] <=  8'h00;      memory[5819] <=  8'h00;      memory[5820] <=  8'h00;      memory[5821] <=  8'h00;      memory[5822] <=  8'h00;      memory[5823] <=  8'h00;      memory[5824] <=  8'h00;      memory[5825] <=  8'h00;      memory[5826] <=  8'h00;      memory[5827] <=  8'h00;      memory[5828] <=  8'h00;      memory[5829] <=  8'h00;      memory[5830] <=  8'h00;      memory[5831] <=  8'h00;      memory[5832] <=  8'h00;      memory[5833] <=  8'h00;      memory[5834] <=  8'h00;      memory[5835] <=  8'h00;      memory[5836] <=  8'h00;      memory[5837] <=  8'h00;      memory[5838] <=  8'h00;      memory[5839] <=  8'h00;      memory[5840] <=  8'h00;      memory[5841] <=  8'h00;      memory[5842] <=  8'h00;      memory[5843] <=  8'h00;      memory[5844] <=  8'h00;      memory[5845] <=  8'h00;      memory[5846] <=  8'h00;      memory[5847] <=  8'h00;      memory[5848] <=  8'h00;      memory[5849] <=  8'h00;      memory[5850] <=  8'h00;      memory[5851] <=  8'h00;      memory[5852] <=  8'h00;      memory[5853] <=  8'h00;      memory[5854] <=  8'h00;      memory[5855] <=  8'h00;      memory[5856] <=  8'h00;      memory[5857] <=  8'h00;      memory[5858] <=  8'h00;      memory[5859] <=  8'h00;      memory[5860] <=  8'h00;      memory[5861] <=  8'h00;      memory[5862] <=  8'h00;      memory[5863] <=  8'h00;      memory[5864] <=  8'h00;      memory[5865] <=  8'h00;      memory[5866] <=  8'h00;      memory[5867] <=  8'h00;      memory[5868] <=  8'h00;      memory[5869] <=  8'h00;      memory[5870] <=  8'h00;      memory[5871] <=  8'h00;      memory[5872] <=  8'h00;      memory[5873] <=  8'h00;      memory[5874] <=  8'h00;      memory[5875] <=  8'h00;      memory[5876] <=  8'h00;      memory[5877] <=  8'h00;      memory[5878] <=  8'h00;      memory[5879] <=  8'h00;      memory[5880] <=  8'h00;      memory[5881] <=  8'h00;      memory[5882] <=  8'h00;      memory[5883] <=  8'h00;      memory[5884] <=  8'h00;      memory[5885] <=  8'h00;      memory[5886] <=  8'h00;      memory[5887] <=  8'h00;      memory[5888] <=  8'h00;      memory[5889] <=  8'h00;      memory[5890] <=  8'h00;      memory[5891] <=  8'h00;      memory[5892] <=  8'h00;      memory[5893] <=  8'h00;      memory[5894] <=  8'h00;      memory[5895] <=  8'h00;      memory[5896] <=  8'h00;      memory[5897] <=  8'h00;      memory[5898] <=  8'h00;      memory[5899] <=  8'h00;      memory[5900] <=  8'h00;      memory[5901] <=  8'h00;      memory[5902] <=  8'h00;      memory[5903] <=  8'h00;      memory[5904] <=  8'h00;      memory[5905] <=  8'h00;      memory[5906] <=  8'h00;      memory[5907] <=  8'h00;      memory[5908] <=  8'h00;      memory[5909] <=  8'h00;      memory[5910] <=  8'h00;      memory[5911] <=  8'h00;      memory[5912] <=  8'h00;      memory[5913] <=  8'h00;      memory[5914] <=  8'h00;      memory[5915] <=  8'h00;      memory[5916] <=  8'h00;      memory[5917] <=  8'h00;      memory[5918] <=  8'h00;      memory[5919] <=  8'h00;      memory[5920] <=  8'h00;      memory[5921] <=  8'h00;      memory[5922] <=  8'h00;      memory[5923] <=  8'h00;      memory[5924] <=  8'h00;      memory[5925] <=  8'h00;      memory[5926] <=  8'h00;      memory[5927] <=  8'h00;      memory[5928] <=  8'h00;      memory[5929] <=  8'h00;      memory[5930] <=  8'h00;      memory[5931] <=  8'h00;      memory[5932] <=  8'h00;      memory[5933] <=  8'h00;      memory[5934] <=  8'h00;      memory[5935] <=  8'h00;      memory[5936] <=  8'h00;      memory[5937] <=  8'h00;      memory[5938] <=  8'h00;      memory[5939] <=  8'h00;      memory[5940] <=  8'h00;      memory[5941] <=  8'h00;      memory[5942] <=  8'h00;      memory[5943] <=  8'h00;      memory[5944] <=  8'h00;      memory[5945] <=  8'h00;      memory[5946] <=  8'h00;      memory[5947] <=  8'h00;      memory[5948] <=  8'h00;      memory[5949] <=  8'h00;      memory[5950] <=  8'h00;      memory[5951] <=  8'h00;      memory[5952] <=  8'h00;      memory[5953] <=  8'h00;      memory[5954] <=  8'h00;      memory[5955] <=  8'h00;      memory[5956] <=  8'h00;      memory[5957] <=  8'h00;      memory[5958] <=  8'h00;      memory[5959] <=  8'h00;      memory[5960] <=  8'h00;      memory[5961] <=  8'h00;      memory[5962] <=  8'h00;      memory[5963] <=  8'h00;      memory[5964] <=  8'h00;      memory[5965] <=  8'h00;      memory[5966] <=  8'h00;      memory[5967] <=  8'h00;      memory[5968] <=  8'h00;      memory[5969] <=  8'h00;      memory[5970] <=  8'h00;      memory[5971] <=  8'h00;      memory[5972] <=  8'h00;      memory[5973] <=  8'h00;      memory[5974] <=  8'h00;      memory[5975] <=  8'h00;      memory[5976] <=  8'h00;      memory[5977] <=  8'h00;      memory[5978] <=  8'h00;      memory[5979] <=  8'h00;      memory[5980] <=  8'h00;      memory[5981] <=  8'h00;      memory[5982] <=  8'h00;      memory[5983] <=  8'h00;      memory[5984] <=  8'h00;      memory[5985] <=  8'h00;      memory[5986] <=  8'h00;      memory[5987] <=  8'h00;      memory[5988] <=  8'h00;      memory[5989] <=  8'h00;      memory[5990] <=  8'h00;      memory[5991] <=  8'h00;      memory[5992] <=  8'h00;      memory[5993] <=  8'h00;      memory[5994] <=  8'h00;      memory[5995] <=  8'h00;      memory[5996] <=  8'h00;      memory[5997] <=  8'h00;      memory[5998] <=  8'h00;      memory[5999] <=  8'h00;      memory[6000] <=  8'h00;      memory[6001] <=  8'h00;      memory[6002] <=  8'h00;      memory[6003] <=  8'h00;      memory[6004] <=  8'h00;      memory[6005] <=  8'h00;      memory[6006] <=  8'h00;      memory[6007] <=  8'h00;      memory[6008] <=  8'h00;      memory[6009] <=  8'h00;      memory[6010] <=  8'h00;      memory[6011] <=  8'h00;      memory[6012] <=  8'h00;      memory[6013] <=  8'h00;      memory[6014] <=  8'h00;      memory[6015] <=  8'h00;      memory[6016] <=  8'h00;      memory[6017] <=  8'h00;      memory[6018] <=  8'h00;      memory[6019] <=  8'h00;      memory[6020] <=  8'h00;      memory[6021] <=  8'h00;      memory[6022] <=  8'h00;      memory[6023] <=  8'h00;      memory[6024] <=  8'h00;      memory[6025] <=  8'h00;      memory[6026] <=  8'h00;      memory[6027] <=  8'h00;      memory[6028] <=  8'h00;      memory[6029] <=  8'h00;      memory[6030] <=  8'h00;      memory[6031] <=  8'h00;      memory[6032] <=  8'h00;      memory[6033] <=  8'h00;      memory[6034] <=  8'h00;      memory[6035] <=  8'h00;      memory[6036] <=  8'h00;      memory[6037] <=  8'h00;      memory[6038] <=  8'h00;      memory[6039] <=  8'h00;      memory[6040] <=  8'h00;      memory[6041] <=  8'h00;      memory[6042] <=  8'h00;      memory[6043] <=  8'h00;      memory[6044] <=  8'h00;      memory[6045] <=  8'h00;      memory[6046] <=  8'h00;      memory[6047] <=  8'h00;      memory[6048] <=  8'h00;      memory[6049] <=  8'h00;      memory[6050] <=  8'h00;      memory[6051] <=  8'h00;      memory[6052] <=  8'h00;      memory[6053] <=  8'h00;      memory[6054] <=  8'h00;      memory[6055] <=  8'h00;      memory[6056] <=  8'h00;      memory[6057] <=  8'h00;      memory[6058] <=  8'h00;      memory[6059] <=  8'h00;      memory[6060] <=  8'h00;      memory[6061] <=  8'h00;      memory[6062] <=  8'h00;      memory[6063] <=  8'h00;      memory[6064] <=  8'h00;      memory[6065] <=  8'h00;      memory[6066] <=  8'h00;      memory[6067] <=  8'h00;      memory[6068] <=  8'h00;      memory[6069] <=  8'h00;      memory[6070] <=  8'h00;      memory[6071] <=  8'h00;      memory[6072] <=  8'h00;      memory[6073] <=  8'h00;      memory[6074] <=  8'h00;      memory[6075] <=  8'h00;      memory[6076] <=  8'h00;      memory[6077] <=  8'h00;      memory[6078] <=  8'h00;      memory[6079] <=  8'h00;      memory[6080] <=  8'h00;      memory[6081] <=  8'h00;      memory[6082] <=  8'h00;      memory[6083] <=  8'h00;      memory[6084] <=  8'h00;      memory[6085] <=  8'h00;      memory[6086] <=  8'h00;      memory[6087] <=  8'h00;      memory[6088] <=  8'h00;      memory[6089] <=  8'h00;      memory[6090] <=  8'h00;      memory[6091] <=  8'h00;      memory[6092] <=  8'h00;      memory[6093] <=  8'h00;      memory[6094] <=  8'h00;      memory[6095] <=  8'h00;      memory[6096] <=  8'h00;      memory[6097] <=  8'h00;      memory[6098] <=  8'h00;      memory[6099] <=  8'h00;      memory[6100] <=  8'h00;      memory[6101] <=  8'h00;      memory[6102] <=  8'h00;      memory[6103] <=  8'h00;      memory[6104] <=  8'h00;      memory[6105] <=  8'h00;      memory[6106] <=  8'h00;      memory[6107] <=  8'h00;      memory[6108] <=  8'h00;      memory[6109] <=  8'h00;      memory[6110] <=  8'h00;      memory[6111] <=  8'h00;      memory[6112] <=  8'h00;      memory[6113] <=  8'h00;      memory[6114] <=  8'h00;      memory[6115] <=  8'h00;      memory[6116] <=  8'h00;      memory[6117] <=  8'h00;      memory[6118] <=  8'h00;      memory[6119] <=  8'h00;      memory[6120] <=  8'h00;      memory[6121] <=  8'h00;      memory[6122] <=  8'h00;      memory[6123] <=  8'h00;      memory[6124] <=  8'h00;      memory[6125] <=  8'h00;      memory[6126] <=  8'h00;      memory[6127] <=  8'h00;      memory[6128] <=  8'h00;      memory[6129] <=  8'h00;      memory[6130] <=  8'h00;      memory[6131] <=  8'h00;      memory[6132] <=  8'h00;      memory[6133] <=  8'h00;      memory[6134] <=  8'h00;      memory[6135] <=  8'h00;      memory[6136] <=  8'h00;      memory[6137] <=  8'h00;      memory[6138] <=  8'h00;      memory[6139] <=  8'h00;      memory[6140] <=  8'h00;      memory[6141] <=  8'h00;      memory[6142] <=  8'h00;      memory[6143] <=  8'h00;      memory[6144] <=  8'h00;      memory[6145] <=  8'h00;      memory[6146] <=  8'h00;      memory[6147] <=  8'h00;      memory[6148] <=  8'h00;      memory[6149] <=  8'h00;      memory[6150] <=  8'h00;      memory[6151] <=  8'h00;      memory[6152] <=  8'h00;      memory[6153] <=  8'h00;      memory[6154] <=  8'h00;      memory[6155] <=  8'h00;      memory[6156] <=  8'h00;      memory[6157] <=  8'h00;      memory[6158] <=  8'h00;      memory[6159] <=  8'h00;      memory[6160] <=  8'h00;      memory[6161] <=  8'h00;      memory[6162] <=  8'h00;      memory[6163] <=  8'h00;      memory[6164] <=  8'h00;      memory[6165] <=  8'h00;      memory[6166] <=  8'h00;      memory[6167] <=  8'h00;      memory[6168] <=  8'h00;      memory[6169] <=  8'h00;      memory[6170] <=  8'h00;      memory[6171] <=  8'h00;      memory[6172] <=  8'h00;      memory[6173] <=  8'h00;      memory[6174] <=  8'h00;      memory[6175] <=  8'h00;      memory[6176] <=  8'h00;      memory[6177] <=  8'h00;      memory[6178] <=  8'h00;      memory[6179] <=  8'h00;      memory[6180] <=  8'h00;      memory[6181] <=  8'h00;      memory[6182] <=  8'h00;      memory[6183] <=  8'h00;      memory[6184] <=  8'h00;      memory[6185] <=  8'h00;      memory[6186] <=  8'h00;      memory[6187] <=  8'h00;      memory[6188] <=  8'h00;      memory[6189] <=  8'h00;      memory[6190] <=  8'h00;      memory[6191] <=  8'h00;      memory[6192] <=  8'h00;      memory[6193] <=  8'h00;      memory[6194] <=  8'h00;      memory[6195] <=  8'h00;      memory[6196] <=  8'h00;      memory[6197] <=  8'h00;      memory[6198] <=  8'h00;      memory[6199] <=  8'h00;      memory[6200] <=  8'h00;      memory[6201] <=  8'h00;      memory[6202] <=  8'h00;      memory[6203] <=  8'h00;      memory[6204] <=  8'h00;      memory[6205] <=  8'h00;      memory[6206] <=  8'h00;      memory[6207] <=  8'h00;      memory[6208] <=  8'h00;      memory[6209] <=  8'h00;      memory[6210] <=  8'h00;      memory[6211] <=  8'h00;      memory[6212] <=  8'h00;      memory[6213] <=  8'h00;      memory[6214] <=  8'h00;      memory[6215] <=  8'h00;      memory[6216] <=  8'h00;      memory[6217] <=  8'h00;      memory[6218] <=  8'h00;      memory[6219] <=  8'h00;      memory[6220] <=  8'h00;      memory[6221] <=  8'h00;      memory[6222] <=  8'h00;      memory[6223] <=  8'h00;      memory[6224] <=  8'h00;      memory[6225] <=  8'h00;      memory[6226] <=  8'h00;      memory[6227] <=  8'h00;      memory[6228] <=  8'h00;      memory[6229] <=  8'h00;      memory[6230] <=  8'h00;      memory[6231] <=  8'h00;      memory[6232] <=  8'h00;      memory[6233] <=  8'h00;      memory[6234] <=  8'h00;      memory[6235] <=  8'h00;      memory[6236] <=  8'h00;      memory[6237] <=  8'h00;      memory[6238] <=  8'h00;      memory[6239] <=  8'h00;      memory[6240] <=  8'h00;      memory[6241] <=  8'h00;      memory[6242] <=  8'h00;      memory[6243] <=  8'h00;      memory[6244] <=  8'h00;      memory[6245] <=  8'h00;      memory[6246] <=  8'h00;      memory[6247] <=  8'h00;      memory[6248] <=  8'h00;      memory[6249] <=  8'h00;      memory[6250] <=  8'h00;      memory[6251] <=  8'h00;      memory[6252] <=  8'h00;      memory[6253] <=  8'h00;      memory[6254] <=  8'h00;      memory[6255] <=  8'h00;      memory[6256] <=  8'h00;      memory[6257] <=  8'h00;      memory[6258] <=  8'h00;      memory[6259] <=  8'h00;      memory[6260] <=  8'h00;      memory[6261] <=  8'h00;      memory[6262] <=  8'h00;      memory[6263] <=  8'h00;      memory[6264] <=  8'h00;      memory[6265] <=  8'h00;      memory[6266] <=  8'h00;      memory[6267] <=  8'h00;      memory[6268] <=  8'h00;      memory[6269] <=  8'h00;      memory[6270] <=  8'h00;      memory[6271] <=  8'h00;      memory[6272] <=  8'h00;      memory[6273] <=  8'h00;      memory[6274] <=  8'h00;      memory[6275] <=  8'h00;      memory[6276] <=  8'h00;      memory[6277] <=  8'h00;      memory[6278] <=  8'h00;      memory[6279] <=  8'h00;      memory[6280] <=  8'h00;      memory[6281] <=  8'h00;      memory[6282] <=  8'h00;      memory[6283] <=  8'h00;      memory[6284] <=  8'h00;      memory[6285] <=  8'h00;      memory[6286] <=  8'h00;      memory[6287] <=  8'h00;      memory[6288] <=  8'h00;      memory[6289] <=  8'h00;      memory[6290] <=  8'h00;      memory[6291] <=  8'h00;      memory[6292] <=  8'h00;      memory[6293] <=  8'h00;      memory[6294] <=  8'h00;      memory[6295] <=  8'h00;      memory[6296] <=  8'h00;      memory[6297] <=  8'h00;      memory[6298] <=  8'h00;      memory[6299] <=  8'h00;      memory[6300] <=  8'h00;      memory[6301] <=  8'h00;      memory[6302] <=  8'h00;      memory[6303] <=  8'h00;      memory[6304] <=  8'h00;      memory[6305] <=  8'h00;      memory[6306] <=  8'h00;      memory[6307] <=  8'h00;      memory[6308] <=  8'h00;      memory[6309] <=  8'h00;      memory[6310] <=  8'h00;      memory[6311] <=  8'h00;      memory[6312] <=  8'h00;      memory[6313] <=  8'h00;      memory[6314] <=  8'h00;      memory[6315] <=  8'h00;      memory[6316] <=  8'h00;      memory[6317] <=  8'h00;      memory[6318] <=  8'h00;      memory[6319] <=  8'h00;      memory[6320] <=  8'h00;      memory[6321] <=  8'h00;      memory[6322] <=  8'h00;      memory[6323] <=  8'h00;      memory[6324] <=  8'h00;      memory[6325] <=  8'h00;      memory[6326] <=  8'h00;      memory[6327] <=  8'h00;      memory[6328] <=  8'h00;      memory[6329] <=  8'h00;      memory[6330] <=  8'h00;      memory[6331] <=  8'h00;      memory[6332] <=  8'h00;      memory[6333] <=  8'h00;      memory[6334] <=  8'h00;      memory[6335] <=  8'h00;      memory[6336] <=  8'h00;      memory[6337] <=  8'h00;      memory[6338] <=  8'h00;      memory[6339] <=  8'h00;      memory[6340] <=  8'h00;      memory[6341] <=  8'h00;      memory[6342] <=  8'h00;      memory[6343] <=  8'h00;      memory[6344] <=  8'h00;      memory[6345] <=  8'h00;      memory[6346] <=  8'h00;      memory[6347] <=  8'h00;      memory[6348] <=  8'h00;      memory[6349] <=  8'h00;      memory[6350] <=  8'h00;      memory[6351] <=  8'h00;      memory[6352] <=  8'h00;      memory[6353] <=  8'h00;      memory[6354] <=  8'h00;      memory[6355] <=  8'h00;      memory[6356] <=  8'h00;      memory[6357] <=  8'h00;      memory[6358] <=  8'h00;      memory[6359] <=  8'h00;      memory[6360] <=  8'h00;      memory[6361] <=  8'h00;      memory[6362] <=  8'h00;      memory[6363] <=  8'h00;      memory[6364] <=  8'h00;      memory[6365] <=  8'h00;      memory[6366] <=  8'h00;      memory[6367] <=  8'h00;      memory[6368] <=  8'h00;      memory[6369] <=  8'h00;      memory[6370] <=  8'h00;      memory[6371] <=  8'h00;      memory[6372] <=  8'h00;      memory[6373] <=  8'h00;      memory[6374] <=  8'h00;      memory[6375] <=  8'h00;      memory[6376] <=  8'h00;      memory[6377] <=  8'h00;      memory[6378] <=  8'h00;      memory[6379] <=  8'h00;      memory[6380] <=  8'h00;      memory[6381] <=  8'h00;      memory[6382] <=  8'h00;      memory[6383] <=  8'h00;      memory[6384] <=  8'h00;      memory[6385] <=  8'h00;      memory[6386] <=  8'h00;      memory[6387] <=  8'h00;      memory[6388] <=  8'h00;      memory[6389] <=  8'h00;      memory[6390] <=  8'h00;      memory[6391] <=  8'h00;      memory[6392] <=  8'h00;      memory[6393] <=  8'h00;      memory[6394] <=  8'h00;      memory[6395] <=  8'h00;      memory[6396] <=  8'h00;      memory[6397] <=  8'h00;      memory[6398] <=  8'h00;      memory[6399] <=  8'h00;      memory[6400] <=  8'h00;      memory[6401] <=  8'h00;      memory[6402] <=  8'h00;      memory[6403] <=  8'h00;      memory[6404] <=  8'h00;      memory[6405] <=  8'h00;      memory[6406] <=  8'h00;      memory[6407] <=  8'h00;      memory[6408] <=  8'h00;      memory[6409] <=  8'h00;      memory[6410] <=  8'h00;      memory[6411] <=  8'h00;      memory[6412] <=  8'h00;      memory[6413] <=  8'h00;      memory[6414] <=  8'h00;      memory[6415] <=  8'h00;      memory[6416] <=  8'h00;      memory[6417] <=  8'h00;      memory[6418] <=  8'h00;      memory[6419] <=  8'h00;      memory[6420] <=  8'h00;      memory[6421] <=  8'h00;      memory[6422] <=  8'h00;      memory[6423] <=  8'h00;      memory[6424] <=  8'h00;      memory[6425] <=  8'h00;      memory[6426] <=  8'h00;      memory[6427] <=  8'h00;      memory[6428] <=  8'h00;      memory[6429] <=  8'h00;      memory[6430] <=  8'h00;      memory[6431] <=  8'h00;      memory[6432] <=  8'h00;      memory[6433] <=  8'h00;      memory[6434] <=  8'h00;      memory[6435] <=  8'h00;      memory[6436] <=  8'h00;      memory[6437] <=  8'h00;      memory[6438] <=  8'h00;      memory[6439] <=  8'h00;      memory[6440] <=  8'h00;      memory[6441] <=  8'h00;      memory[6442] <=  8'h00;      memory[6443] <=  8'h00;      memory[6444] <=  8'h00;      memory[6445] <=  8'h00;      memory[6446] <=  8'h00;      memory[6447] <=  8'h00;      memory[6448] <=  8'h00;      memory[6449] <=  8'h00;      memory[6450] <=  8'h00;      memory[6451] <=  8'h00;      memory[6452] <=  8'h00;      memory[6453] <=  8'h00;      memory[6454] <=  8'h00;      memory[6455] <=  8'h00;      memory[6456] <=  8'h00;      memory[6457] <=  8'h00;      memory[6458] <=  8'h00;      memory[6459] <=  8'h00;      memory[6460] <=  8'h00;      memory[6461] <=  8'h00;      memory[6462] <=  8'h00;      memory[6463] <=  8'h00;      memory[6464] <=  8'h00;      memory[6465] <=  8'h00;      memory[6466] <=  8'h00;      memory[6467] <=  8'h00;      memory[6468] <=  8'h00;      memory[6469] <=  8'h00;      memory[6470] <=  8'h00;      memory[6471] <=  8'h00;      memory[6472] <=  8'h00;      memory[6473] <=  8'h00;      memory[6474] <=  8'h00;      memory[6475] <=  8'h00;      memory[6476] <=  8'h00;      memory[6477] <=  8'h00;      memory[6478] <=  8'h00;      memory[6479] <=  8'h00;      memory[6480] <=  8'h00;      memory[6481] <=  8'h00;      memory[6482] <=  8'h00;      memory[6483] <=  8'h00;      memory[6484] <=  8'h00;      memory[6485] <=  8'h00;      memory[6486] <=  8'h00;      memory[6487] <=  8'h00;      memory[6488] <=  8'h00;      memory[6489] <=  8'h00;      memory[6490] <=  8'h00;      memory[6491] <=  8'h00;      memory[6492] <=  8'h00;      memory[6493] <=  8'h00;      memory[6494] <=  8'h00;      memory[6495] <=  8'h00;      memory[6496] <=  8'h00;      memory[6497] <=  8'h00;      memory[6498] <=  8'h00;      memory[6499] <=  8'h00;      memory[6500] <=  8'h00;      memory[6501] <=  8'h00;      memory[6502] <=  8'h00;      memory[6503] <=  8'h00;      memory[6504] <=  8'h00;      memory[6505] <=  8'h00;      memory[6506] <=  8'h00;      memory[6507] <=  8'h00;      memory[6508] <=  8'h00;      memory[6509] <=  8'h00;      memory[6510] <=  8'h00;      memory[6511] <=  8'h00;      memory[6512] <=  8'h00;      memory[6513] <=  8'h00;      memory[6514] <=  8'h00;      memory[6515] <=  8'h00;      memory[6516] <=  8'h00;      memory[6517] <=  8'h00;      memory[6518] <=  8'h00;      memory[6519] <=  8'h00;      memory[6520] <=  8'h00;      memory[6521] <=  8'h00;      memory[6522] <=  8'h00;      memory[6523] <=  8'h00;      memory[6524] <=  8'h00;      memory[6525] <=  8'h00;      memory[6526] <=  8'h00;      memory[6527] <=  8'h00;      memory[6528] <=  8'h00;      memory[6529] <=  8'h00;      memory[6530] <=  8'h00;      memory[6531] <=  8'h00;      memory[6532] <=  8'h00;      memory[6533] <=  8'h00;      memory[6534] <=  8'h00;      memory[6535] <=  8'h00;      memory[6536] <=  8'h00;      memory[6537] <=  8'h00;      memory[6538] <=  8'h00;      memory[6539] <=  8'h00;      memory[6540] <=  8'h00;      memory[6541] <=  8'h00;      memory[6542] <=  8'h00;      memory[6543] <=  8'h00;      memory[6544] <=  8'h00;      memory[6545] <=  8'h00;      memory[6546] <=  8'h00;      memory[6547] <=  8'h00;      memory[6548] <=  8'h00;      memory[6549] <=  8'h00;      memory[6550] <=  8'h00;      memory[6551] <=  8'h00;      memory[6552] <=  8'h00;      memory[6553] <=  8'h00;      memory[6554] <=  8'h00;      memory[6555] <=  8'h00;      memory[6556] <=  8'h00;      memory[6557] <=  8'h00;      memory[6558] <=  8'h00;      memory[6559] <=  8'h00;      memory[6560] <=  8'h00;      memory[6561] <=  8'h00;      memory[6562] <=  8'h00;      memory[6563] <=  8'h00;      memory[6564] <=  8'h00;      memory[6565] <=  8'h00;      memory[6566] <=  8'h00;      memory[6567] <=  8'h00;      memory[6568] <=  8'h00;      memory[6569] <=  8'h00;      memory[6570] <=  8'h00;      memory[6571] <=  8'h00;      memory[6572] <=  8'h00;      memory[6573] <=  8'h00;      memory[6574] <=  8'h00;      memory[6575] <=  8'h00;      memory[6576] <=  8'h00;      memory[6577] <=  8'h00;      memory[6578] <=  8'h00;      memory[6579] <=  8'h00;      memory[6580] <=  8'h00;      memory[6581] <=  8'h00;      memory[6582] <=  8'h00;      memory[6583] <=  8'h00;      memory[6584] <=  8'h00;      memory[6585] <=  8'h00;      memory[6586] <=  8'h00;      memory[6587] <=  8'h00;      memory[6588] <=  8'h00;      memory[6589] <=  8'h00;      memory[6590] <=  8'h00;      memory[6591] <=  8'h00;      memory[6592] <=  8'h00;      memory[6593] <=  8'h00;      memory[6594] <=  8'h00;      memory[6595] <=  8'h00;      memory[6596] <=  8'h00;      memory[6597] <=  8'h00;      memory[6598] <=  8'h00;      memory[6599] <=  8'h00;      memory[6600] <=  8'h00;      memory[6601] <=  8'h00;      memory[6602] <=  8'h00;      memory[6603] <=  8'h00;      memory[6604] <=  8'h00;      memory[6605] <=  8'h00;      memory[6606] <=  8'h00;      memory[6607] <=  8'h00;      memory[6608] <=  8'h00;      memory[6609] <=  8'h00;      memory[6610] <=  8'h00;      memory[6611] <=  8'h00;      memory[6612] <=  8'h00;      memory[6613] <=  8'h00;      memory[6614] <=  8'h00;      memory[6615] <=  8'h00;      memory[6616] <=  8'h00;      memory[6617] <=  8'h00;      memory[6618] <=  8'h00;      memory[6619] <=  8'h00;      memory[6620] <=  8'h00;      memory[6621] <=  8'h00;      memory[6622] <=  8'h00;      memory[6623] <=  8'h00;      memory[6624] <=  8'h00;      memory[6625] <=  8'h00;      memory[6626] <=  8'h00;      memory[6627] <=  8'h00;      memory[6628] <=  8'h00;      memory[6629] <=  8'h00;      memory[6630] <=  8'h00;      memory[6631] <=  8'h00;      memory[6632] <=  8'h00;      memory[6633] <=  8'h00;      memory[6634] <=  8'h00;      memory[6635] <=  8'h00;      memory[6636] <=  8'h00;      memory[6637] <=  8'h00;      memory[6638] <=  8'h00;      memory[6639] <=  8'h00;      memory[6640] <=  8'h00;      memory[6641] <=  8'h00;      memory[6642] <=  8'h00;      memory[6643] <=  8'h00;      memory[6644] <=  8'h00;      memory[6645] <=  8'h00;      memory[6646] <=  8'h00;      memory[6647] <=  8'h00;      memory[6648] <=  8'h00;      memory[6649] <=  8'h00;      memory[6650] <=  8'h00;      memory[6651] <=  8'h00;      memory[6652] <=  8'h00;      memory[6653] <=  8'h00;      memory[6654] <=  8'h00;      memory[6655] <=  8'h00;      memory[6656] <=  8'h00;      memory[6657] <=  8'h00;      memory[6658] <=  8'h00;      memory[6659] <=  8'h00;      memory[6660] <=  8'h00;      memory[6661] <=  8'h00;      memory[6662] <=  8'h00;      memory[6663] <=  8'h00;      memory[6664] <=  8'h00;      memory[6665] <=  8'h00;      memory[6666] <=  8'h00;      memory[6667] <=  8'h00;      memory[6668] <=  8'h00;      memory[6669] <=  8'h00;      memory[6670] <=  8'h00;      memory[6671] <=  8'h00;      memory[6672] <=  8'h00;      memory[6673] <=  8'h00;      memory[6674] <=  8'h00;      memory[6675] <=  8'h00;      memory[6676] <=  8'h00;      memory[6677] <=  8'h00;      memory[6678] <=  8'h00;      memory[6679] <=  8'h00;      memory[6680] <=  8'h00;      memory[6681] <=  8'h00;      memory[6682] <=  8'h00;      memory[6683] <=  8'h00;      memory[6684] <=  8'h00;      memory[6685] <=  8'h00;      memory[6686] <=  8'h00;      memory[6687] <=  8'h00;      memory[6688] <=  8'h00;      memory[6689] <=  8'h00;      memory[6690] <=  8'h00;      memory[6691] <=  8'h00;      memory[6692] <=  8'h00;      memory[6693] <=  8'h00;      memory[6694] <=  8'h00;      memory[6695] <=  8'h00;      memory[6696] <=  8'h00;      memory[6697] <=  8'h00;      memory[6698] <=  8'h00;      memory[6699] <=  8'h00;      memory[6700] <=  8'h00;      memory[6701] <=  8'h00;      memory[6702] <=  8'h00;      memory[6703] <=  8'h00;      memory[6704] <=  8'h00;      memory[6705] <=  8'h00;      memory[6706] <=  8'h00;      memory[6707] <=  8'h00;      memory[6708] <=  8'h00;      memory[6709] <=  8'h00;      memory[6710] <=  8'h00;      memory[6711] <=  8'h00;      memory[6712] <=  8'h00;      memory[6713] <=  8'h00;      memory[6714] <=  8'h00;      memory[6715] <=  8'h00;      memory[6716] <=  8'h00;      memory[6717] <=  8'h00;      memory[6718] <=  8'h00;      memory[6719] <=  8'h00;      memory[6720] <=  8'h00;      memory[6721] <=  8'h00;      memory[6722] <=  8'h00;      memory[6723] <=  8'h00;      memory[6724] <=  8'h00;      memory[6725] <=  8'h00;      memory[6726] <=  8'h00;      memory[6727] <=  8'h00;      memory[6728] <=  8'h00;      memory[6729] <=  8'h00;      memory[6730] <=  8'h00;      memory[6731] <=  8'h00;      memory[6732] <=  8'h00;      memory[6733] <=  8'h00;      memory[6734] <=  8'h00;      memory[6735] <=  8'h00;      memory[6736] <=  8'h00;      memory[6737] <=  8'h00;      memory[6738] <=  8'h00;      memory[6739] <=  8'h00;      memory[6740] <=  8'h00;      memory[6741] <=  8'h00;      memory[6742] <=  8'h00;      memory[6743] <=  8'h00;      memory[6744] <=  8'h00;      memory[6745] <=  8'h00;      memory[6746] <=  8'h00;      memory[6747] <=  8'h00;      memory[6748] <=  8'h00;      memory[6749] <=  8'h00;      memory[6750] <=  8'h00;      memory[6751] <=  8'h00;      memory[6752] <=  8'h00;      memory[6753] <=  8'h00;      memory[6754] <=  8'h00;      memory[6755] <=  8'h00;      memory[6756] <=  8'h00;      memory[6757] <=  8'h00;      memory[6758] <=  8'h00;      memory[6759] <=  8'h00;      memory[6760] <=  8'h00;      memory[6761] <=  8'h00;      memory[6762] <=  8'h00;      memory[6763] <=  8'h00;      memory[6764] <=  8'h00;      memory[6765] <=  8'h00;      memory[6766] <=  8'h00;      memory[6767] <=  8'h00;      memory[6768] <=  8'h00;      memory[6769] <=  8'h00;      memory[6770] <=  8'h00;      memory[6771] <=  8'h00;      memory[6772] <=  8'h00;      memory[6773] <=  8'h00;      memory[6774] <=  8'h00;      memory[6775] <=  8'h00;      memory[6776] <=  8'h00;      memory[6777] <=  8'h00;      memory[6778] <=  8'h00;      memory[6779] <=  8'h00;      memory[6780] <=  8'h00;      memory[6781] <=  8'h00;      memory[6782] <=  8'h00;      memory[6783] <=  8'h00;      memory[6784] <=  8'h00;      memory[6785] <=  8'h00;      memory[6786] <=  8'h00;      memory[6787] <=  8'h00;      memory[6788] <=  8'h00;      memory[6789] <=  8'h00;      memory[6790] <=  8'h00;      memory[6791] <=  8'h00;      memory[6792] <=  8'h00;      memory[6793] <=  8'h00;      memory[6794] <=  8'h00;      memory[6795] <=  8'h00;      memory[6796] <=  8'h00;      memory[6797] <=  8'h00;      memory[6798] <=  8'h00;      memory[6799] <=  8'h00;      memory[6800] <=  8'h00;      memory[6801] <=  8'h00;      memory[6802] <=  8'h00;      memory[6803] <=  8'h00;      memory[6804] <=  8'h00;      memory[6805] <=  8'h00;      memory[6806] <=  8'h00;      memory[6807] <=  8'h00;      memory[6808] <=  8'h00;      memory[6809] <=  8'h00;      memory[6810] <=  8'h00;      memory[6811] <=  8'h00;      memory[6812] <=  8'h00;      memory[6813] <=  8'h00;      memory[6814] <=  8'h00;      memory[6815] <=  8'h00;      memory[6816] <=  8'h00;      memory[6817] <=  8'h00;      memory[6818] <=  8'h00;      memory[6819] <=  8'h00;      memory[6820] <=  8'h00;      memory[6821] <=  8'h00;      memory[6822] <=  8'h00;      memory[6823] <=  8'h00;      memory[6824] <=  8'h00;      memory[6825] <=  8'h00;      memory[6826] <=  8'h00;      memory[6827] <=  8'h00;      memory[6828] <=  8'h00;      memory[6829] <=  8'h00;      memory[6830] <=  8'h00;      memory[6831] <=  8'h00;      memory[6832] <=  8'h00;      memory[6833] <=  8'h00;      memory[6834] <=  8'h00;      memory[6835] <=  8'h00;      memory[6836] <=  8'h00;      memory[6837] <=  8'h00;      memory[6838] <=  8'h00;      memory[6839] <=  8'h00;      memory[6840] <=  8'h00;      memory[6841] <=  8'h00;      memory[6842] <=  8'h00;      memory[6843] <=  8'h00;      memory[6844] <=  8'h00;      memory[6845] <=  8'h00;      memory[6846] <=  8'h00;      memory[6847] <=  8'h00;      memory[6848] <=  8'h00;      memory[6849] <=  8'h00;      memory[6850] <=  8'h00;      memory[6851] <=  8'h00;      memory[6852] <=  8'h00;      memory[6853] <=  8'h00;      memory[6854] <=  8'h00;      memory[6855] <=  8'h00;      memory[6856] <=  8'h00;      memory[6857] <=  8'h00;      memory[6858] <=  8'h00;      memory[6859] <=  8'h00;      memory[6860] <=  8'h00;      memory[6861] <=  8'h00;      memory[6862] <=  8'h00;      memory[6863] <=  8'h00;      memory[6864] <=  8'h00;      memory[6865] <=  8'h00;      memory[6866] <=  8'h00;      memory[6867] <=  8'h00;      memory[6868] <=  8'h00;      memory[6869] <=  8'h00;      memory[6870] <=  8'h00;      memory[6871] <=  8'h00;      memory[6872] <=  8'h00;      memory[6873] <=  8'h00;      memory[6874] <=  8'h00;      memory[6875] <=  8'h00;      memory[6876] <=  8'h00;      memory[6877] <=  8'h00;      memory[6878] <=  8'h00;      memory[6879] <=  8'h00;      memory[6880] <=  8'h00;      memory[6881] <=  8'h00;      memory[6882] <=  8'h00;      memory[6883] <=  8'h00;      memory[6884] <=  8'h00;      memory[6885] <=  8'h00;      memory[6886] <=  8'h00;      memory[6887] <=  8'h00;      memory[6888] <=  8'h00;      memory[6889] <=  8'h00;      memory[6890] <=  8'h00;      memory[6891] <=  8'h00;      memory[6892] <=  8'h00;      memory[6893] <=  8'h00;      memory[6894] <=  8'h00;      memory[6895] <=  8'h00;      memory[6896] <=  8'h00;      memory[6897] <=  8'h00;      memory[6898] <=  8'h00;      memory[6899] <=  8'h00;      memory[6900] <=  8'h00;      memory[6901] <=  8'h00;      memory[6902] <=  8'h00;      memory[6903] <=  8'h00;      memory[6904] <=  8'h00;      memory[6905] <=  8'h00;      memory[6906] <=  8'h00;      memory[6907] <=  8'h00;      memory[6908] <=  8'h00;      memory[6909] <=  8'h00;      memory[6910] <=  8'h00;      memory[6911] <=  8'h00;      memory[6912] <=  8'h00;      memory[6913] <=  8'h00;      memory[6914] <=  8'h00;      memory[6915] <=  8'h00;      memory[6916] <=  8'h00;      memory[6917] <=  8'h00;      memory[6918] <=  8'h00;      memory[6919] <=  8'h00;      memory[6920] <=  8'h00;      memory[6921] <=  8'h00;      memory[6922] <=  8'h00;      memory[6923] <=  8'h00;      memory[6924] <=  8'h00;      memory[6925] <=  8'h00;      memory[6926] <=  8'h00;      memory[6927] <=  8'h00;      memory[6928] <=  8'h00;      memory[6929] <=  8'h00;      memory[6930] <=  8'h00;      memory[6931] <=  8'h00;      memory[6932] <=  8'h00;      memory[6933] <=  8'h00;      memory[6934] <=  8'h00;      memory[6935] <=  8'h00;      memory[6936] <=  8'h00;      memory[6937] <=  8'h00;      memory[6938] <=  8'h00;      memory[6939] <=  8'h00;      memory[6940] <=  8'h00;      memory[6941] <=  8'h00;      memory[6942] <=  8'h00;      memory[6943] <=  8'h00;      memory[6944] <=  8'h00;      memory[6945] <=  8'h00;      memory[6946] <=  8'h00;      memory[6947] <=  8'h00;      memory[6948] <=  8'h00;      memory[6949] <=  8'h00;      memory[6950] <=  8'h00;      memory[6951] <=  8'h00;      memory[6952] <=  8'h00;      memory[6953] <=  8'h00;      memory[6954] <=  8'h00;      memory[6955] <=  8'h00;      memory[6956] <=  8'h00;      memory[6957] <=  8'h00;      memory[6958] <=  8'h00;      memory[6959] <=  8'h00;      memory[6960] <=  8'h00;      memory[6961] <=  8'h00;      memory[6962] <=  8'h00;      memory[6963] <=  8'h00;      memory[6964] <=  8'h00;      memory[6965] <=  8'h00;      memory[6966] <=  8'h00;      memory[6967] <=  8'h00;      memory[6968] <=  8'h00;      memory[6969] <=  8'h00;      memory[6970] <=  8'h00;      memory[6971] <=  8'h00;      memory[6972] <=  8'h00;      memory[6973] <=  8'h00;      memory[6974] <=  8'h00;      memory[6975] <=  8'h00;      memory[6976] <=  8'h00;      memory[6977] <=  8'h00;      memory[6978] <=  8'h00;      memory[6979] <=  8'h00;      memory[6980] <=  8'h00;      memory[6981] <=  8'h00;      memory[6982] <=  8'h00;      memory[6983] <=  8'h00;      memory[6984] <=  8'h00;      memory[6985] <=  8'h00;      memory[6986] <=  8'h00;      memory[6987] <=  8'h00;      memory[6988] <=  8'h00;      memory[6989] <=  8'h00;      memory[6990] <=  8'h00;      memory[6991] <=  8'h00;      memory[6992] <=  8'h00;      memory[6993] <=  8'h00;      memory[6994] <=  8'h00;      memory[6995] <=  8'h00;      memory[6996] <=  8'h00;      memory[6997] <=  8'h00;      memory[6998] <=  8'h00;      memory[6999] <=  8'h00;      memory[7000] <=  8'h00;      memory[7001] <=  8'h00;      memory[7002] <=  8'h00;      memory[7003] <=  8'h00;      memory[7004] <=  8'h00;      memory[7005] <=  8'h00;      memory[7006] <=  8'h00;      memory[7007] <=  8'h00;      memory[7008] <=  8'h00;      memory[7009] <=  8'h00;      memory[7010] <=  8'h00;      memory[7011] <=  8'h00;      memory[7012] <=  8'h00;      memory[7013] <=  8'h00;      memory[7014] <=  8'h00;      memory[7015] <=  8'h00;      memory[7016] <=  8'h00;      memory[7017] <=  8'h00;      memory[7018] <=  8'h00;      memory[7019] <=  8'h00;      memory[7020] <=  8'h00;      memory[7021] <=  8'h00;      memory[7022] <=  8'h00;      memory[7023] <=  8'h00;      memory[7024] <=  8'h00;      memory[7025] <=  8'h00;      memory[7026] <=  8'h00;      memory[7027] <=  8'h00;      memory[7028] <=  8'h00;      memory[7029] <=  8'h00;      memory[7030] <=  8'h00;      memory[7031] <=  8'h00;      memory[7032] <=  8'h00;      memory[7033] <=  8'h00;      memory[7034] <=  8'h00;      memory[7035] <=  8'h00;      memory[7036] <=  8'h00;      memory[7037] <=  8'h00;      memory[7038] <=  8'h00;      memory[7039] <=  8'h00;      memory[7040] <=  8'h00;      memory[7041] <=  8'h00;      memory[7042] <=  8'h00;      memory[7043] <=  8'h00;      memory[7044] <=  8'h00;      memory[7045] <=  8'h00;      memory[7046] <=  8'h00;      memory[7047] <=  8'h00;      memory[7048] <=  8'h00;      memory[7049] <=  8'h00;      memory[7050] <=  8'h00;      memory[7051] <=  8'h00;      memory[7052] <=  8'h00;      memory[7053] <=  8'h00;      memory[7054] <=  8'h00;      memory[7055] <=  8'h00;      memory[7056] <=  8'h00;      memory[7057] <=  8'h00;      memory[7058] <=  8'h00;      memory[7059] <=  8'h00;      memory[7060] <=  8'h00;      memory[7061] <=  8'h00;      memory[7062] <=  8'h00;      memory[7063] <=  8'h00;      memory[7064] <=  8'h00;      memory[7065] <=  8'h00;      memory[7066] <=  8'h00;      memory[7067] <=  8'h00;      memory[7068] <=  8'h00;      memory[7069] <=  8'h00;      memory[7070] <=  8'h00;      memory[7071] <=  8'h00;      memory[7072] <=  8'h00;      memory[7073] <=  8'h00;      memory[7074] <=  8'h00;      memory[7075] <=  8'h00;      memory[7076] <=  8'h00;      memory[7077] <=  8'h00;      memory[7078] <=  8'h00;      memory[7079] <=  8'h00;      memory[7080] <=  8'h00;      memory[7081] <=  8'h00;      memory[7082] <=  8'h00;      memory[7083] <=  8'h00;      memory[7084] <=  8'h00;      memory[7085] <=  8'h00;      memory[7086] <=  8'h00;      memory[7087] <=  8'h00;      memory[7088] <=  8'h00;      memory[7089] <=  8'h00;      memory[7090] <=  8'h00;      memory[7091] <=  8'h00;      memory[7092] <=  8'h00;      memory[7093] <=  8'h00;      memory[7094] <=  8'h00;      memory[7095] <=  8'h00;      memory[7096] <=  8'h00;      memory[7097] <=  8'h00;      memory[7098] <=  8'h00;      memory[7099] <=  8'h00;      memory[7100] <=  8'h00;      memory[7101] <=  8'h00;      memory[7102] <=  8'h00;      memory[7103] <=  8'h00;      memory[7104] <=  8'h00;      memory[7105] <=  8'h00;      memory[7106] <=  8'h00;      memory[7107] <=  8'h00;      memory[7108] <=  8'h00;      memory[7109] <=  8'h00;      memory[7110] <=  8'h00;      memory[7111] <=  8'h00;      memory[7112] <=  8'h00;      memory[7113] <=  8'h00;      memory[7114] <=  8'h00;      memory[7115] <=  8'h00;      memory[7116] <=  8'h00;      memory[7117] <=  8'h00;      memory[7118] <=  8'h00;      memory[7119] <=  8'h00;      memory[7120] <=  8'h00;      memory[7121] <=  8'h00;      memory[7122] <=  8'h00;      memory[7123] <=  8'h00;      memory[7124] <=  8'h00;      memory[7125] <=  8'h00;      memory[7126] <=  8'h00;      memory[7127] <=  8'h00;      memory[7128] <=  8'h00;      memory[7129] <=  8'h00;      memory[7130] <=  8'h00;      memory[7131] <=  8'h00;      memory[7132] <=  8'h00;      memory[7133] <=  8'h00;      memory[7134] <=  8'h00;      memory[7135] <=  8'h00;      memory[7136] <=  8'h00;      memory[7137] <=  8'h00;      memory[7138] <=  8'h00;      memory[7139] <=  8'h00;      memory[7140] <=  8'h00;      memory[7141] <=  8'h00;      memory[7142] <=  8'h00;      memory[7143] <=  8'h00;      memory[7144] <=  8'h00;      memory[7145] <=  8'h00;      memory[7146] <=  8'h00;      memory[7147] <=  8'h00;      memory[7148] <=  8'h00;      memory[7149] <=  8'h00;      memory[7150] <=  8'h00;      memory[7151] <=  8'h00;      memory[7152] <=  8'h00;      memory[7153] <=  8'h00;      memory[7154] <=  8'h00;      memory[7155] <=  8'h00;      memory[7156] <=  8'h00;      memory[7157] <=  8'h00;      memory[7158] <=  8'h00;      memory[7159] <=  8'h00;      memory[7160] <=  8'h00;      memory[7161] <=  8'h00;      memory[7162] <=  8'h00;      memory[7163] <=  8'h00;      memory[7164] <=  8'h00;      memory[7165] <=  8'h00;      memory[7166] <=  8'h00;      memory[7167] <=  8'h00;      memory[7168] <=  8'h00;      memory[7169] <=  8'h00;      memory[7170] <=  8'h00;      memory[7171] <=  8'h00;      memory[7172] <=  8'h00;      memory[7173] <=  8'h00;      memory[7174] <=  8'h00;      memory[7175] <=  8'h00;      memory[7176] <=  8'h00;      memory[7177] <=  8'h00;      memory[7178] <=  8'h00;      memory[7179] <=  8'h00;      memory[7180] <=  8'h00;      memory[7181] <=  8'h00;      memory[7182] <=  8'h00;      memory[7183] <=  8'h00;      memory[7184] <=  8'h00;      memory[7185] <=  8'h00;      memory[7186] <=  8'h00;      memory[7187] <=  8'h00;      memory[7188] <=  8'h00;      memory[7189] <=  8'h00;      memory[7190] <=  8'h00;      memory[7191] <=  8'h00;      memory[7192] <=  8'h00;      memory[7193] <=  8'h00;      memory[7194] <=  8'h00;      memory[7195] <=  8'h00;      memory[7196] <=  8'h00;      memory[7197] <=  8'h00;      memory[7198] <=  8'h00;      memory[7199] <=  8'h00;      memory[7200] <=  8'h00;      memory[7201] <=  8'h00;      memory[7202] <=  8'h00;      memory[7203] <=  8'h00;      memory[7204] <=  8'h00;      memory[7205] <=  8'h00;      memory[7206] <=  8'h00;      memory[7207] <=  8'h00;      memory[7208] <=  8'h00;      memory[7209] <=  8'h00;      memory[7210] <=  8'h00;      memory[7211] <=  8'h00;      memory[7212] <=  8'h00;      memory[7213] <=  8'h00;      memory[7214] <=  8'h00;      memory[7215] <=  8'h00;      memory[7216] <=  8'h00;      memory[7217] <=  8'h00;      memory[7218] <=  8'h00;      memory[7219] <=  8'h00;      memory[7220] <=  8'h00;      memory[7221] <=  8'h00;      memory[7222] <=  8'h00;      memory[7223] <=  8'h00;      memory[7224] <=  8'h00;      memory[7225] <=  8'h00;      memory[7226] <=  8'h00;      memory[7227] <=  8'h00;      memory[7228] <=  8'h00;      memory[7229] <=  8'h00;      memory[7230] <=  8'h00;      memory[7231] <=  8'h00;      memory[7232] <=  8'h00;      memory[7233] <=  8'h00;      memory[7234] <=  8'h00;      memory[7235] <=  8'h00;      memory[7236] <=  8'h00;      memory[7237] <=  8'h00;      memory[7238] <=  8'h00;      memory[7239] <=  8'h00;      memory[7240] <=  8'h00;      memory[7241] <=  8'h00;      memory[7242] <=  8'h00;      memory[7243] <=  8'h00;      memory[7244] <=  8'h00;      memory[7245] <=  8'h00;      memory[7246] <=  8'h00;      memory[7247] <=  8'h00;      memory[7248] <=  8'h00;      memory[7249] <=  8'h00;      memory[7250] <=  8'h00;      memory[7251] <=  8'h00;      memory[7252] <=  8'h00;      memory[7253] <=  8'h00;      memory[7254] <=  8'h00;      memory[7255] <=  8'h00;      memory[7256] <=  8'h00;      memory[7257] <=  8'h00;      memory[7258] <=  8'h00;      memory[7259] <=  8'h00;      memory[7260] <=  8'h00;      memory[7261] <=  8'h00;      memory[7262] <=  8'h00;      memory[7263] <=  8'h00;      memory[7264] <=  8'h00;      memory[7265] <=  8'h00;      memory[7266] <=  8'h00;      memory[7267] <=  8'h00;      memory[7268] <=  8'h00;      memory[7269] <=  8'h00;      memory[7270] <=  8'h00;      memory[7271] <=  8'h00;      memory[7272] <=  8'h00;      memory[7273] <=  8'h00;      memory[7274] <=  8'h00;      memory[7275] <=  8'h00;      memory[7276] <=  8'h00;      memory[7277] <=  8'h00;      memory[7278] <=  8'h00;      memory[7279] <=  8'h00;      memory[7280] <=  8'h00;      memory[7281] <=  8'h00;      memory[7282] <=  8'h00;      memory[7283] <=  8'h00;      memory[7284] <=  8'h00;      memory[7285] <=  8'h00;      memory[7286] <=  8'h00;      memory[7287] <=  8'h00;      memory[7288] <=  8'h00;      memory[7289] <=  8'h00;      memory[7290] <=  8'h00;      memory[7291] <=  8'h00;      memory[7292] <=  8'h00;      memory[7293] <=  8'h00;      memory[7294] <=  8'h00;      memory[7295] <=  8'h00;      memory[7296] <=  8'h00;      memory[7297] <=  8'h00;      memory[7298] <=  8'h00;      memory[7299] <=  8'h00;      memory[7300] <=  8'h00;      memory[7301] <=  8'h00;      memory[7302] <=  8'h00;      memory[7303] <=  8'h00;      memory[7304] <=  8'h00;      memory[7305] <=  8'h00;      memory[7306] <=  8'h00;      memory[7307] <=  8'h00;      memory[7308] <=  8'h00;      memory[7309] <=  8'h00;      memory[7310] <=  8'h00;      memory[7311] <=  8'h00;      memory[7312] <=  8'h00;      memory[7313] <=  8'h00;      memory[7314] <=  8'h00;      memory[7315] <=  8'h00;      memory[7316] <=  8'h00;      memory[7317] <=  8'h00;      memory[7318] <=  8'h00;      memory[7319] <=  8'h00;      memory[7320] <=  8'h00;      memory[7321] <=  8'h00;      memory[7322] <=  8'h00;      memory[7323] <=  8'h00;      memory[7324] <=  8'h00;      memory[7325] <=  8'h00;      memory[7326] <=  8'h00;      memory[7327] <=  8'h00;      memory[7328] <=  8'h00;      memory[7329] <=  8'h00;      memory[7330] <=  8'h00;      memory[7331] <=  8'h00;      memory[7332] <=  8'h00;      memory[7333] <=  8'h00;      memory[7334] <=  8'h00;      memory[7335] <=  8'h00;      memory[7336] <=  8'h00;      memory[7337] <=  8'h00;      memory[7338] <=  8'h00;      memory[7339] <=  8'h00;      memory[7340] <=  8'h00;      memory[7341] <=  8'h00;      memory[7342] <=  8'h00;      memory[7343] <=  8'h00;      memory[7344] <=  8'h00;      memory[7345] <=  8'h00;      memory[7346] <=  8'h00;      memory[7347] <=  8'h00;      memory[7348] <=  8'h00;      memory[7349] <=  8'h00;      memory[7350] <=  8'h00;      memory[7351] <=  8'h00;      memory[7352] <=  8'h00;      memory[7353] <=  8'h00;      memory[7354] <=  8'h00;      memory[7355] <=  8'h00;      memory[7356] <=  8'h00;      memory[7357] <=  8'h00;      memory[7358] <=  8'h00;      memory[7359] <=  8'h00;      memory[7360] <=  8'h00;      memory[7361] <=  8'h00;      memory[7362] <=  8'h00;      memory[7363] <=  8'h00;      memory[7364] <=  8'h00;      memory[7365] <=  8'h00;      memory[7366] <=  8'h00;      memory[7367] <=  8'h00;      memory[7368] <=  8'h00;      memory[7369] <=  8'h00;      memory[7370] <=  8'h00;      memory[7371] <=  8'h00;      memory[7372] <=  8'h00;      memory[7373] <=  8'h00;      memory[7374] <=  8'h00;      memory[7375] <=  8'h00;      memory[7376] <=  8'h00;      memory[7377] <=  8'h00;      memory[7378] <=  8'h00;      memory[7379] <=  8'h00;      memory[7380] <=  8'h00;      memory[7381] <=  8'h00;      memory[7382] <=  8'h00;      memory[7383] <=  8'h00;      memory[7384] <=  8'h00;      memory[7385] <=  8'h00;      memory[7386] <=  8'h00;      memory[7387] <=  8'h00;      memory[7388] <=  8'h00;      memory[7389] <=  8'h00;      memory[7390] <=  8'h00;      memory[7391] <=  8'h00;      memory[7392] <=  8'h00;      memory[7393] <=  8'h00;      memory[7394] <=  8'h00;      memory[7395] <=  8'h00;      memory[7396] <=  8'h00;      memory[7397] <=  8'h00;      memory[7398] <=  8'h00;      memory[7399] <=  8'h00;      memory[7400] <=  8'h00;      memory[7401] <=  8'h00;      memory[7402] <=  8'h00;      memory[7403] <=  8'h00;      memory[7404] <=  8'h00;      memory[7405] <=  8'h00;      memory[7406] <=  8'h00;      memory[7407] <=  8'h00;      memory[7408] <=  8'h00;      memory[7409] <=  8'h00;      memory[7410] <=  8'h00;      memory[7411] <=  8'h00;      memory[7412] <=  8'h00;      memory[7413] <=  8'h00;      memory[7414] <=  8'h00;      memory[7415] <=  8'h00;      memory[7416] <=  8'h00;      memory[7417] <=  8'h00;      memory[7418] <=  8'h00;      memory[7419] <=  8'h00;      memory[7420] <=  8'h00;      memory[7421] <=  8'h00;      memory[7422] <=  8'h00;      memory[7423] <=  8'h00;      memory[7424] <=  8'h00;      memory[7425] <=  8'h00;      memory[7426] <=  8'h00;      memory[7427] <=  8'h00;      memory[7428] <=  8'h00;      memory[7429] <=  8'h00;      memory[7430] <=  8'h00;      memory[7431] <=  8'h00;      memory[7432] <=  8'h00;      memory[7433] <=  8'h00;      memory[7434] <=  8'h00;      memory[7435] <=  8'h00;      memory[7436] <=  8'h00;      memory[7437] <=  8'h00;      memory[7438] <=  8'h00;      memory[7439] <=  8'h00;      memory[7440] <=  8'h00;      memory[7441] <=  8'h00;      memory[7442] <=  8'h00;      memory[7443] <=  8'h00;      memory[7444] <=  8'h00;      memory[7445] <=  8'h00;      memory[7446] <=  8'h00;      memory[7447] <=  8'h00;      memory[7448] <=  8'h00;      memory[7449] <=  8'h00;      memory[7450] <=  8'h00;      memory[7451] <=  8'h00;      memory[7452] <=  8'h00;      memory[7453] <=  8'h00;      memory[7454] <=  8'h00;      memory[7455] <=  8'h00;      memory[7456] <=  8'h00;      memory[7457] <=  8'h00;      memory[7458] <=  8'h00;      memory[7459] <=  8'h00;      memory[7460] <=  8'h00;      memory[7461] <=  8'h00;      memory[7462] <=  8'h00;      memory[7463] <=  8'h00;      memory[7464] <=  8'h00;      memory[7465] <=  8'h00;      memory[7466] <=  8'h00;      memory[7467] <=  8'h00;      memory[7468] <=  8'h00;      memory[7469] <=  8'h00;      memory[7470] <=  8'h00;      memory[7471] <=  8'h00;      memory[7472] <=  8'h00;      memory[7473] <=  8'h00;      memory[7474] <=  8'h00;      memory[7475] <=  8'h00;      memory[7476] <=  8'h00;      memory[7477] <=  8'h00;      memory[7478] <=  8'h00;      memory[7479] <=  8'h00;      memory[7480] <=  8'h00;      memory[7481] <=  8'h00;      memory[7482] <=  8'h00;      memory[7483] <=  8'h00;      memory[7484] <=  8'h00;      memory[7485] <=  8'h00;      memory[7486] <=  8'h00;      memory[7487] <=  8'h00;      memory[7488] <=  8'h00;      memory[7489] <=  8'h00;      memory[7490] <=  8'h00;      memory[7491] <=  8'h00;      memory[7492] <=  8'h00;      memory[7493] <=  8'h00;      memory[7494] <=  8'h00;      memory[7495] <=  8'h00;      memory[7496] <=  8'h00;      memory[7497] <=  8'h00;      memory[7498] <=  8'h00;      memory[7499] <=  8'h00;      memory[7500] <=  8'h00;      memory[7501] <=  8'h00;      memory[7502] <=  8'h00;      memory[7503] <=  8'h00;      memory[7504] <=  8'h00;      memory[7505] <=  8'h00;      memory[7506] <=  8'h00;      memory[7507] <=  8'h00;      memory[7508] <=  8'h00;      memory[7509] <=  8'h00;      memory[7510] <=  8'h00;      memory[7511] <=  8'h00;      memory[7512] <=  8'h00;      memory[7513] <=  8'h00;      memory[7514] <=  8'h00;      memory[7515] <=  8'h00;      memory[7516] <=  8'h00;      memory[7517] <=  8'h00;      memory[7518] <=  8'h00;      memory[7519] <=  8'h00;      memory[7520] <=  8'h00;      memory[7521] <=  8'h00;      memory[7522] <=  8'h00;      memory[7523] <=  8'h00;      memory[7524] <=  8'h00;      memory[7525] <=  8'h00;      memory[7526] <=  8'h00;      memory[7527] <=  8'h00;      memory[7528] <=  8'h00;      memory[7529] <=  8'h00;      memory[7530] <=  8'h00;      memory[7531] <=  8'h00;      memory[7532] <=  8'h00;      memory[7533] <=  8'h00;      memory[7534] <=  8'h00;      memory[7535] <=  8'h00;      memory[7536] <=  8'h00;      memory[7537] <=  8'h00;      memory[7538] <=  8'h00;      memory[7539] <=  8'h00;      memory[7540] <=  8'h00;      memory[7541] <=  8'h00;      memory[7542] <=  8'h00;      memory[7543] <=  8'h00;      memory[7544] <=  8'h00;      memory[7545] <=  8'h00;      memory[7546] <=  8'h00;      memory[7547] <=  8'h00;      memory[7548] <=  8'h00;      memory[7549] <=  8'h00;      memory[7550] <=  8'h00;      memory[7551] <=  8'h00;      memory[7552] <=  8'h00;      memory[7553] <=  8'h00;      memory[7554] <=  8'h00;      memory[7555] <=  8'h00;      memory[7556] <=  8'h00;      memory[7557] <=  8'h00;      memory[7558] <=  8'h00;      memory[7559] <=  8'h00;      memory[7560] <=  8'h00;      memory[7561] <=  8'h00;      memory[7562] <=  8'h00;      memory[7563] <=  8'h00;      memory[7564] <=  8'h00;      memory[7565] <=  8'h00;      memory[7566] <=  8'h00;      memory[7567] <=  8'h00;      memory[7568] <=  8'h00;      memory[7569] <=  8'h00;      memory[7570] <=  8'h00;      memory[7571] <=  8'h00;      memory[7572] <=  8'h00;      memory[7573] <=  8'h00;      memory[7574] <=  8'h00;      memory[7575] <=  8'h00;      memory[7576] <=  8'h00;      memory[7577] <=  8'h00;      memory[7578] <=  8'h00;      memory[7579] <=  8'h00;      memory[7580] <=  8'h00;      memory[7581] <=  8'h00;      memory[7582] <=  8'h00;      memory[7583] <=  8'h00;      memory[7584] <=  8'h00;      memory[7585] <=  8'h00;      memory[7586] <=  8'h00;      memory[7587] <=  8'h00;      memory[7588] <=  8'h00;      memory[7589] <=  8'h00;      memory[7590] <=  8'h00;      memory[7591] <=  8'h00;      memory[7592] <=  8'h00;      memory[7593] <=  8'h00;      memory[7594] <=  8'h00;      memory[7595] <=  8'h00;      memory[7596] <=  8'h00;      memory[7597] <=  8'h00;      memory[7598] <=  8'h00;      memory[7599] <=  8'h00;      memory[7600] <=  8'h00;      memory[7601] <=  8'h00;      memory[7602] <=  8'h00;      memory[7603] <=  8'h00;      memory[7604] <=  8'h00;      memory[7605] <=  8'h00;      memory[7606] <=  8'h00;      memory[7607] <=  8'h00;      memory[7608] <=  8'h00;      memory[7609] <=  8'h00;      memory[7610] <=  8'h00;      memory[7611] <=  8'h00;      memory[7612] <=  8'h00;      memory[7613] <=  8'h00;      memory[7614] <=  8'h00;      memory[7615] <=  8'h00;      memory[7616] <=  8'h00;      memory[7617] <=  8'h00;      memory[7618] <=  8'h00;      memory[7619] <=  8'h00;      memory[7620] <=  8'h00;      memory[7621] <=  8'h00;      memory[7622] <=  8'h00;      memory[7623] <=  8'h00;      memory[7624] <=  8'h00;      memory[7625] <=  8'h00;      memory[7626] <=  8'h00;      memory[7627] <=  8'h00;      memory[7628] <=  8'h00;      memory[7629] <=  8'h00;      memory[7630] <=  8'h00;      memory[7631] <=  8'h00;      memory[7632] <=  8'h00;      memory[7633] <=  8'h00;      memory[7634] <=  8'h00;      memory[7635] <=  8'h00;      memory[7636] <=  8'h00;      memory[7637] <=  8'h00;      memory[7638] <=  8'h00;      memory[7639] <=  8'h00;      memory[7640] <=  8'h00;      memory[7641] <=  8'h00;      memory[7642] <=  8'h00;      memory[7643] <=  8'h00;      memory[7644] <=  8'h00;      memory[7645] <=  8'h00;      memory[7646] <=  8'h00;      memory[7647] <=  8'h00;      memory[7648] <=  8'h00;      memory[7649] <=  8'h00;      memory[7650] <=  8'h00;      memory[7651] <=  8'h00;      memory[7652] <=  8'h00;      memory[7653] <=  8'h00;      memory[7654] <=  8'h00;      memory[7655] <=  8'h00;      memory[7656] <=  8'h00;      memory[7657] <=  8'h00;      memory[7658] <=  8'h00;      memory[7659] <=  8'h00;      memory[7660] <=  8'h00;      memory[7661] <=  8'h00;      memory[7662] <=  8'h00;      memory[7663] <=  8'h00;      memory[7664] <=  8'h00;      memory[7665] <=  8'h00;      memory[7666] <=  8'h00;      memory[7667] <=  8'h00;      memory[7668] <=  8'h00;      memory[7669] <=  8'h00;      memory[7670] <=  8'h00;      memory[7671] <=  8'h00;      memory[7672] <=  8'h00;      memory[7673] <=  8'h00;      memory[7674] <=  8'h00;      memory[7675] <=  8'h00;      memory[7676] <=  8'h00;      memory[7677] <=  8'h00;      memory[7678] <=  8'h00;      memory[7679] <=  8'h00;      memory[7680] <=  8'h00;      memory[7681] <=  8'h00;      memory[7682] <=  8'h00;      memory[7683] <=  8'h00;      memory[7684] <=  8'h00;      memory[7685] <=  8'h00;      memory[7686] <=  8'h00;      memory[7687] <=  8'h00;      memory[7688] <=  8'h00;      memory[7689] <=  8'h00;      memory[7690] <=  8'h00;      memory[7691] <=  8'h00;      memory[7692] <=  8'h00;      memory[7693] <=  8'h00;      memory[7694] <=  8'h00;      memory[7695] <=  8'h00;      memory[7696] <=  8'h00;      memory[7697] <=  8'h00;      memory[7698] <=  8'h00;      memory[7699] <=  8'h00;      memory[7700] <=  8'h00;      memory[7701] <=  8'h00;      memory[7702] <=  8'h00;      memory[7703] <=  8'h00;      memory[7704] <=  8'h00;      memory[7705] <=  8'h00;      memory[7706] <=  8'h00;      memory[7707] <=  8'h00;      memory[7708] <=  8'h00;      memory[7709] <=  8'h00;      memory[7710] <=  8'h00;      memory[7711] <=  8'h00;      memory[7712] <=  8'h00;      memory[7713] <=  8'h00;      memory[7714] <=  8'h00;      memory[7715] <=  8'h00;      memory[7716] <=  8'h00;      memory[7717] <=  8'h00;      memory[7718] <=  8'h00;      memory[7719] <=  8'h00;      memory[7720] <=  8'h00;      memory[7721] <=  8'h00;      memory[7722] <=  8'h00;      memory[7723] <=  8'h00;      memory[7724] <=  8'h00;      memory[7725] <=  8'h00;      memory[7726] <=  8'h00;      memory[7727] <=  8'h00;      memory[7728] <=  8'h00;      memory[7729] <=  8'h00;      memory[7730] <=  8'h00;      memory[7731] <=  8'h00;      memory[7732] <=  8'h00;      memory[7733] <=  8'h00;      memory[7734] <=  8'h00;      memory[7735] <=  8'h00;      memory[7736] <=  8'h00;      memory[7737] <=  8'h00;      memory[7738] <=  8'h00;      memory[7739] <=  8'h00;      memory[7740] <=  8'h00;      memory[7741] <=  8'h00;      memory[7742] <=  8'h00;      memory[7743] <=  8'h00;      memory[7744] <=  8'h00;      memory[7745] <=  8'h00;      memory[7746] <=  8'h00;      memory[7747] <=  8'h00;      memory[7748] <=  8'h00;      memory[7749] <=  8'h00;      memory[7750] <=  8'h00;      memory[7751] <=  8'h00;      memory[7752] <=  8'h00;      memory[7753] <=  8'h00;      memory[7754] <=  8'h00;      memory[7755] <=  8'h00;      memory[7756] <=  8'h00;      memory[7757] <=  8'h00;      memory[7758] <=  8'h00;      memory[7759] <=  8'h00;      memory[7760] <=  8'h00;      memory[7761] <=  8'h00;      memory[7762] <=  8'h00;      memory[7763] <=  8'h00;      memory[7764] <=  8'h00;      memory[7765] <=  8'h00;      memory[7766] <=  8'h00;      memory[7767] <=  8'h00;      memory[7768] <=  8'h00;      memory[7769] <=  8'h00;      memory[7770] <=  8'h00;      memory[7771] <=  8'h00;      memory[7772] <=  8'h00;      memory[7773] <=  8'h00;      memory[7774] <=  8'h00;      memory[7775] <=  8'h00;      memory[7776] <=  8'h00;      memory[7777] <=  8'h00;      memory[7778] <=  8'h00;      memory[7779] <=  8'h00;      memory[7780] <=  8'h00;      memory[7781] <=  8'h00;      memory[7782] <=  8'h00;      memory[7783] <=  8'h00;      memory[7784] <=  8'h00;      memory[7785] <=  8'h00;      memory[7786] <=  8'h00;      memory[7787] <=  8'h00;      memory[7788] <=  8'h00;      memory[7789] <=  8'h00;      memory[7790] <=  8'h00;      memory[7791] <=  8'h00;      memory[7792] <=  8'h00;      memory[7793] <=  8'h00;      memory[7794] <=  8'h00;      memory[7795] <=  8'h00;      memory[7796] <=  8'h00;      memory[7797] <=  8'h00;      memory[7798] <=  8'h00;      memory[7799] <=  8'h00;      memory[7800] <=  8'h00;      memory[7801] <=  8'h00;      memory[7802] <=  8'h00;      memory[7803] <=  8'h00;      memory[7804] <=  8'h00;      memory[7805] <=  8'h00;      memory[7806] <=  8'h00;      memory[7807] <=  8'h00;      memory[7808] <=  8'h00;      memory[7809] <=  8'h00;      memory[7810] <=  8'h00;      memory[7811] <=  8'h00;      memory[7812] <=  8'h00;      memory[7813] <=  8'h00;      memory[7814] <=  8'h00;      memory[7815] <=  8'h00;      memory[7816] <=  8'h00;      memory[7817] <=  8'h00;      memory[7818] <=  8'h00;      memory[7819] <=  8'h00;      memory[7820] <=  8'h00;      memory[7821] <=  8'h00;      memory[7822] <=  8'h00;      memory[7823] <=  8'h00;      memory[7824] <=  8'h00;      memory[7825] <=  8'h00;      memory[7826] <=  8'h00;      memory[7827] <=  8'h00;      memory[7828] <=  8'h00;      memory[7829] <=  8'h00;      memory[7830] <=  8'h00;      memory[7831] <=  8'h00;      memory[7832] <=  8'h00;      memory[7833] <=  8'h00;      memory[7834] <=  8'h00;      memory[7835] <=  8'h00;      memory[7836] <=  8'h00;      memory[7837] <=  8'h00;      memory[7838] <=  8'h00;      memory[7839] <=  8'h00;      memory[7840] <=  8'h00;      memory[7841] <=  8'h00;      memory[7842] <=  8'h00;      memory[7843] <=  8'h00;      memory[7844] <=  8'h00;      memory[7845] <=  8'h00;      memory[7846] <=  8'h00;      memory[7847] <=  8'h00;      memory[7848] <=  8'h00;      memory[7849] <=  8'h00;      memory[7850] <=  8'h00;      memory[7851] <=  8'h00;      memory[7852] <=  8'h00;      memory[7853] <=  8'h00;      memory[7854] <=  8'h00;      memory[7855] <=  8'h00;      memory[7856] <=  8'h00;      memory[7857] <=  8'h00;      memory[7858] <=  8'h00;      memory[7859] <=  8'h00;      memory[7860] <=  8'h00;      memory[7861] <=  8'h00;      memory[7862] <=  8'h00;      memory[7863] <=  8'h00;      memory[7864] <=  8'h00;      memory[7865] <=  8'h00;      memory[7866] <=  8'h00;      memory[7867] <=  8'h00;      memory[7868] <=  8'h00;      memory[7869] <=  8'h00;      memory[7870] <=  8'h00;      memory[7871] <=  8'h00;      memory[7872] <=  8'h00;      memory[7873] <=  8'h00;      memory[7874] <=  8'h00;      memory[7875] <=  8'h00;      memory[7876] <=  8'h00;      memory[7877] <=  8'h00;      memory[7878] <=  8'h00;      memory[7879] <=  8'h00;      memory[7880] <=  8'h00;      memory[7881] <=  8'h00;      memory[7882] <=  8'h00;      memory[7883] <=  8'h00;      memory[7884] <=  8'h00;      memory[7885] <=  8'h00;      memory[7886] <=  8'h00;      memory[7887] <=  8'h00;      memory[7888] <=  8'h00;      memory[7889] <=  8'h00;      memory[7890] <=  8'h00;      memory[7891] <=  8'h00;      memory[7892] <=  8'h00;      memory[7893] <=  8'h00;      memory[7894] <=  8'h00;      memory[7895] <=  8'h00;      memory[7896] <=  8'h00;      memory[7897] <=  8'h00;      memory[7898] <=  8'h00;      memory[7899] <=  8'h00;      memory[7900] <=  8'h00;      memory[7901] <=  8'h00;      memory[7902] <=  8'h00;      memory[7903] <=  8'h00;      memory[7904] <=  8'h00;      memory[7905] <=  8'h00;      memory[7906] <=  8'h00;      memory[7907] <=  8'h00;      memory[7908] <=  8'h00;      memory[7909] <=  8'h00;      memory[7910] <=  8'h00;      memory[7911] <=  8'h00;      memory[7912] <=  8'h00;      memory[7913] <=  8'h00;      memory[7914] <=  8'h00;      memory[7915] <=  8'h00;      memory[7916] <=  8'h00;      memory[7917] <=  8'h00;      memory[7918] <=  8'h00;      memory[7919] <=  8'h00;      memory[7920] <=  8'h00;      memory[7921] <=  8'h00;      memory[7922] <=  8'h00;      memory[7923] <=  8'h00;      memory[7924] <=  8'h00;      memory[7925] <=  8'h00;      memory[7926] <=  8'h00;      memory[7927] <=  8'h00;      memory[7928] <=  8'h00;      memory[7929] <=  8'h00;      memory[7930] <=  8'h00;      memory[7931] <=  8'h00;      memory[7932] <=  8'h00;      memory[7933] <=  8'h00;      memory[7934] <=  8'h00;      memory[7935] <=  8'h00;      memory[7936] <=  8'h00;      memory[7937] <=  8'h00;      memory[7938] <=  8'h00;      memory[7939] <=  8'h00;      memory[7940] <=  8'h00;      memory[7941] <=  8'h00;      memory[7942] <=  8'h00;      memory[7943] <=  8'h00;      memory[7944] <=  8'h00;      memory[7945] <=  8'h00;      memory[7946] <=  8'h00;      memory[7947] <=  8'h00;      memory[7948] <=  8'h00;      memory[7949] <=  8'h00;      memory[7950] <=  8'h00;      memory[7951] <=  8'h00;      memory[7952] <=  8'h00;      memory[7953] <=  8'h00;      memory[7954] <=  8'h00;      memory[7955] <=  8'h00;      memory[7956] <=  8'h00;      memory[7957] <=  8'h00;      memory[7958] <=  8'h00;      memory[7959] <=  8'h00;      memory[7960] <=  8'h00;      memory[7961] <=  8'h00;      memory[7962] <=  8'h00;      memory[7963] <=  8'h00;      memory[7964] <=  8'h00;      memory[7965] <=  8'h00;      memory[7966] <=  8'h00;      memory[7967] <=  8'h00;      memory[7968] <=  8'h00;      memory[7969] <=  8'h00;      memory[7970] <=  8'h00;      memory[7971] <=  8'h00;      memory[7972] <=  8'h00;      memory[7973] <=  8'h00;      memory[7974] <=  8'h00;      memory[7975] <=  8'h00;      memory[7976] <=  8'h00;      memory[7977] <=  8'h00;      memory[7978] <=  8'h00;      memory[7979] <=  8'h00;      memory[7980] <=  8'h00;      memory[7981] <=  8'h00;      memory[7982] <=  8'h00;      memory[7983] <=  8'h00;      memory[7984] <=  8'h00;      memory[7985] <=  8'h00;      memory[7986] <=  8'h00;      memory[7987] <=  8'h00;      memory[7988] <=  8'h00;      memory[7989] <=  8'h00;      memory[7990] <=  8'h00;      memory[7991] <=  8'h00;      memory[7992] <=  8'h00;      memory[7993] <=  8'h00;      memory[7994] <=  8'h00;      memory[7995] <=  8'h00;      memory[7996] <=  8'h00;      memory[7997] <=  8'h00;      memory[7998] <=  8'h00;      memory[7999] <=  8'h00;      memory[8000] <=  8'h00;      memory[8001] <=  8'h00;      memory[8002] <=  8'h00;      memory[8003] <=  8'h00;      memory[8004] <=  8'h00;      memory[8005] <=  8'h00;      memory[8006] <=  8'h00;      memory[8007] <=  8'h00;      memory[8008] <=  8'h00;      memory[8009] <=  8'h00;      memory[8010] <=  8'h00;      memory[8011] <=  8'h00;      memory[8012] <=  8'h00;      memory[8013] <=  8'h00;      memory[8014] <=  8'h00;      memory[8015] <=  8'h00;      memory[8016] <=  8'h00;      memory[8017] <=  8'h00;      memory[8018] <=  8'h00;      memory[8019] <=  8'h00;      memory[8020] <=  8'h00;      memory[8021] <=  8'h00;      memory[8022] <=  8'h00;      memory[8023] <=  8'h00;      memory[8024] <=  8'h00;      memory[8025] <=  8'h00;      memory[8026] <=  8'h00;      memory[8027] <=  8'h00;      memory[8028] <=  8'h00;      memory[8029] <=  8'h00;      memory[8030] <=  8'h00;      memory[8031] <=  8'h00;      memory[8032] <=  8'h00;      memory[8033] <=  8'h00;      memory[8034] <=  8'h00;      memory[8035] <=  8'h00;      memory[8036] <=  8'h00;      memory[8037] <=  8'h00;      memory[8038] <=  8'h00;      memory[8039] <=  8'h00;      memory[8040] <=  8'h00;      memory[8041] <=  8'h00;      memory[8042] <=  8'h00;      memory[8043] <=  8'h00;      memory[8044] <=  8'h00;      memory[8045] <=  8'h00;      memory[8046] <=  8'h00;      memory[8047] <=  8'h00;      memory[8048] <=  8'h00;      memory[8049] <=  8'h00;      memory[8050] <=  8'h00;      memory[8051] <=  8'h00;      memory[8052] <=  8'h00;      memory[8053] <=  8'h00;      memory[8054] <=  8'h00;      memory[8055] <=  8'h00;      memory[8056] <=  8'h00;      memory[8057] <=  8'h00;      memory[8058] <=  8'h00;      memory[8059] <=  8'h00;      memory[8060] <=  8'h00;      memory[8061] <=  8'h00;      memory[8062] <=  8'h00;      memory[8063] <=  8'h00;      memory[8064] <=  8'h00;      memory[8065] <=  8'h00;      memory[8066] <=  8'h00;      memory[8067] <=  8'h00;      memory[8068] <=  8'h00;      memory[8069] <=  8'h00;      memory[8070] <=  8'h00;      memory[8071] <=  8'h00;      memory[8072] <=  8'h00;      memory[8073] <=  8'h00;      memory[8074] <=  8'h00;      memory[8075] <=  8'h00;      memory[8076] <=  8'h00;      memory[8077] <=  8'h00;      memory[8078] <=  8'h00;      memory[8079] <=  8'h00;      memory[8080] <=  8'h00;      memory[8081] <=  8'h00;      memory[8082] <=  8'h00;      memory[8083] <=  8'h00;      memory[8084] <=  8'h00;      memory[8085] <=  8'h00;      memory[8086] <=  8'h00;      memory[8087] <=  8'h00;      memory[8088] <=  8'h00;      memory[8089] <=  8'h00;      memory[8090] <=  8'h00;      memory[8091] <=  8'h00;      memory[8092] <=  8'h00;      memory[8093] <=  8'h00;      memory[8094] <=  8'h00;      memory[8095] <=  8'h00;      memory[8096] <=  8'h00;      memory[8097] <=  8'h00;      memory[8098] <=  8'h00;      memory[8099] <=  8'h00;      memory[8100] <=  8'h00;      memory[8101] <=  8'h00;      memory[8102] <=  8'h00;      memory[8103] <=  8'h00;      memory[8104] <=  8'h00;      memory[8105] <=  8'h00;      memory[8106] <=  8'h00;      memory[8107] <=  8'h00;      memory[8108] <=  8'h00;      memory[8109] <=  8'h00;      memory[8110] <=  8'h00;      memory[8111] <=  8'h00;      memory[8112] <=  8'h00;      memory[8113] <=  8'h00;      memory[8114] <=  8'h00;      memory[8115] <=  8'h00;      memory[8116] <=  8'h00;      memory[8117] <=  8'h00;      memory[8118] <=  8'h00;      memory[8119] <=  8'h00;      memory[8120] <=  8'h00;      memory[8121] <=  8'h00;      memory[8122] <=  8'h00;      memory[8123] <=  8'h00;      memory[8124] <=  8'h00;      memory[8125] <=  8'h00;      memory[8126] <=  8'h00;      memory[8127] <=  8'h00;      memory[8128] <=  8'h00;      memory[8129] <=  8'h00;      memory[8130] <=  8'h00;      memory[8131] <=  8'h00;      memory[8132] <=  8'h00;      memory[8133] <=  8'h00;      memory[8134] <=  8'h00;      memory[8135] <=  8'h00;      memory[8136] <=  8'h00;      memory[8137] <=  8'h00;      memory[8138] <=  8'h00;      memory[8139] <=  8'h00;      memory[8140] <=  8'h00;      memory[8141] <=  8'h00;      memory[8142] <=  8'h00;      memory[8143] <=  8'h00;      memory[8144] <=  8'h00;      memory[8145] <=  8'h00;      memory[8146] <=  8'h00;      memory[8147] <=  8'h00;      memory[8148] <=  8'h00;      memory[8149] <=  8'h00;      memory[8150] <=  8'h00;      memory[8151] <=  8'h00;      memory[8152] <=  8'h00;      memory[8153] <=  8'h00;      memory[8154] <=  8'h00;      memory[8155] <=  8'h00;      memory[8156] <=  8'h00;      memory[8157] <=  8'h00;      memory[8158] <=  8'h00;      memory[8159] <=  8'h00;      memory[8160] <=  8'h00;      memory[8161] <=  8'h00;      memory[8162] <=  8'h00;      memory[8163] <=  8'h00;      memory[8164] <=  8'h00;      memory[8165] <=  8'h00;      memory[8166] <=  8'h00;      memory[8167] <=  8'h00;      memory[8168] <=  8'h00;      memory[8169] <=  8'h00;      memory[8170] <=  8'h00;      memory[8171] <=  8'h00;      memory[8172] <=  8'h00;      memory[8173] <=  8'h00;      memory[8174] <=  8'h00;      memory[8175] <=  8'h00;      memory[8176] <=  8'h00;      memory[8177] <=  8'h00;      memory[8178] <=  8'h00;      memory[8179] <=  8'h00;      memory[8180] <=  8'h00;      memory[8181] <=  8'h00;      memory[8182] <=  8'h00;      memory[8183] <=  8'h00;      memory[8184] <=  8'h00;      memory[8185] <=  8'h00;      memory[8186] <=  8'h00;      memory[8187] <=  8'h00;      memory[8188] <=  8'h00;      memory[8189] <=  8'h00;      memory[8190] <=  8'h00;      memory[8191] <=  8'h00;      memory[8192] <=  8'h00;      memory[8193] <=  8'h00;      memory[8194] <=  8'h00;      memory[8195] <=  8'h00;      memory[8196] <=  8'h00;      memory[8197] <=  8'h00;      memory[8198] <=  8'h00;      memory[8199] <=  8'h00;      memory[8200] <=  8'h00;      memory[8201] <=  8'h00;      memory[8202] <=  8'h00;      memory[8203] <=  8'h00;      memory[8204] <=  8'h00;      memory[8205] <=  8'h00;      memory[8206] <=  8'h00;      memory[8207] <=  8'h00;      memory[8208] <=  8'h00;      memory[8209] <=  8'h00;      memory[8210] <=  8'h00;      memory[8211] <=  8'h00;      memory[8212] <=  8'h00;      memory[8213] <=  8'h00;      memory[8214] <=  8'h00;      memory[8215] <=  8'h00;      memory[8216] <=  8'h00;      memory[8217] <=  8'h00;      memory[8218] <=  8'h00;      memory[8219] <=  8'h00;      memory[8220] <=  8'h00;      memory[8221] <=  8'h00;      memory[8222] <=  8'h00;      memory[8223] <=  8'h00;      memory[8224] <=  8'h00;      memory[8225] <=  8'h00;      memory[8226] <=  8'h00;      memory[8227] <=  8'h00;      memory[8228] <=  8'h00;      memory[8229] <=  8'h00;      memory[8230] <=  8'h00;      memory[8231] <=  8'h00;      memory[8232] <=  8'h00;      memory[8233] <=  8'h00;      memory[8234] <=  8'h00;      memory[8235] <=  8'h00;      memory[8236] <=  8'h00;      memory[8237] <=  8'h00;      memory[8238] <=  8'h00;      memory[8239] <=  8'h00;      memory[8240] <=  8'h00;      memory[8241] <=  8'h00;      memory[8242] <=  8'h00;      memory[8243] <=  8'h00;      memory[8244] <=  8'h00;      memory[8245] <=  8'h00;      memory[8246] <=  8'h00;      memory[8247] <=  8'h00;      memory[8248] <=  8'h00;      memory[8249] <=  8'h00;      memory[8250] <=  8'h00;      memory[8251] <=  8'h00;      memory[8252] <=  8'h00;      memory[8253] <=  8'h00;      memory[8254] <=  8'h00;      memory[8255] <=  8'h00;      memory[8256] <=  8'h00;      memory[8257] <=  8'h00;      memory[8258] <=  8'h00;      memory[8259] <=  8'h00;      memory[8260] <=  8'h00;      memory[8261] <=  8'h00;      memory[8262] <=  8'h00;      memory[8263] <=  8'h00;      memory[8264] <=  8'h00;      memory[8265] <=  8'h00;      memory[8266] <=  8'h00;      memory[8267] <=  8'h00;      memory[8268] <=  8'h00;      memory[8269] <=  8'h00;      memory[8270] <=  8'h00;      memory[8271] <=  8'h00;      memory[8272] <=  8'h00;      memory[8273] <=  8'h00;      memory[8274] <=  8'h00;      memory[8275] <=  8'h00;      memory[8276] <=  8'h00;      memory[8277] <=  8'h00;      memory[8278] <=  8'h00;      memory[8279] <=  8'h00;      memory[8280] <=  8'h00;      memory[8281] <=  8'h00;      memory[8282] <=  8'h00;      memory[8283] <=  8'h00;      memory[8284] <=  8'h00;      memory[8285] <=  8'h00;      memory[8286] <=  8'h00;      memory[8287] <=  8'h00;      memory[8288] <=  8'h00;      memory[8289] <=  8'h00;      memory[8290] <=  8'h00;      memory[8291] <=  8'h00;      memory[8292] <=  8'h00;      memory[8293] <=  8'h00;      memory[8294] <=  8'h00;      memory[8295] <=  8'h00;      memory[8296] <=  8'h00;      memory[8297] <=  8'h00;      memory[8298] <=  8'h00;      memory[8299] <=  8'h00;      memory[8300] <=  8'h00;      memory[8301] <=  8'h00;      memory[8302] <=  8'h00;      memory[8303] <=  8'h00;      memory[8304] <=  8'h00;      memory[8305] <=  8'h00;      memory[8306] <=  8'h00;      memory[8307] <=  8'h00;      memory[8308] <=  8'h00;      memory[8309] <=  8'h00;      memory[8310] <=  8'h00;      memory[8311] <=  8'h00;      memory[8312] <=  8'h00;      memory[8313] <=  8'h00;      memory[8314] <=  8'h00;      memory[8315] <=  8'h00;      memory[8316] <=  8'h00;      memory[8317] <=  8'h00;      memory[8318] <=  8'h00;      memory[8319] <=  8'h00;      memory[8320] <=  8'h00;      memory[8321] <=  8'h00;      memory[8322] <=  8'h00;      memory[8323] <=  8'h00;      memory[8324] <=  8'h00;      memory[8325] <=  8'h00;      memory[8326] <=  8'h00;      memory[8327] <=  8'h00;      memory[8328] <=  8'h00;      memory[8329] <=  8'h00;      memory[8330] <=  8'h00;      memory[8331] <=  8'h00;      memory[8332] <=  8'h00;      memory[8333] <=  8'h00;      memory[8334] <=  8'h00;      memory[8335] <=  8'h00;      memory[8336] <=  8'h00;      memory[8337] <=  8'h00;      memory[8338] <=  8'h00;      memory[8339] <=  8'h00;      memory[8340] <=  8'h00;      memory[8341] <=  8'h00;      memory[8342] <=  8'h00;      memory[8343] <=  8'h00;      memory[8344] <=  8'h00;      memory[8345] <=  8'h00;      memory[8346] <=  8'h00;      memory[8347] <=  8'h00;      memory[8348] <=  8'h00;      memory[8349] <=  8'h00;      memory[8350] <=  8'h00;      memory[8351] <=  8'h00;      memory[8352] <=  8'h00;      memory[8353] <=  8'h00;      memory[8354] <=  8'h00;      memory[8355] <=  8'h00;      memory[8356] <=  8'h00;      memory[8357] <=  8'h00;      memory[8358] <=  8'h00;      memory[8359] <=  8'h00;      memory[8360] <=  8'h00;      memory[8361] <=  8'h00;      memory[8362] <=  8'h00;      memory[8363] <=  8'h00;      memory[8364] <=  8'h00;      memory[8365] <=  8'h00;      memory[8366] <=  8'h00;      memory[8367] <=  8'h00;      memory[8368] <=  8'h00;      memory[8369] <=  8'h00;      memory[8370] <=  8'h00;      memory[8371] <=  8'h00;      memory[8372] <=  8'h00;      memory[8373] <=  8'h00;      memory[8374] <=  8'h00;      memory[8375] <=  8'h00;      memory[8376] <=  8'h00;      memory[8377] <=  8'h00;      memory[8378] <=  8'h00;      memory[8379] <=  8'h00;      memory[8380] <=  8'h00;      memory[8381] <=  8'h00;      memory[8382] <=  8'h00;      memory[8383] <=  8'h00;      memory[8384] <=  8'h00;      memory[8385] <=  8'h00;      memory[8386] <=  8'h00;      memory[8387] <=  8'h00;      memory[8388] <=  8'h00;      memory[8389] <=  8'h00;      memory[8390] <=  8'h00;      memory[8391] <=  8'h00;      memory[8392] <=  8'h00;      memory[8393] <=  8'h00;      memory[8394] <=  8'h00;      memory[8395] <=  8'h00;      memory[8396] <=  8'h00;      memory[8397] <=  8'h00;      memory[8398] <=  8'h00;      memory[8399] <=  8'h00;      memory[8400] <=  8'h00;      memory[8401] <=  8'h00;      memory[8402] <=  8'h00;      memory[8403] <=  8'h00;      memory[8404] <=  8'h00;      memory[8405] <=  8'h00;      memory[8406] <=  8'h00;      memory[8407] <=  8'h00;      memory[8408] <=  8'h00;      memory[8409] <=  8'h00;      memory[8410] <=  8'h00;      memory[8411] <=  8'h00;      memory[8412] <=  8'h00;      memory[8413] <=  8'h00;      memory[8414] <=  8'h00;      memory[8415] <=  8'h00;      memory[8416] <=  8'h00;      memory[8417] <=  8'h00;      memory[8418] <=  8'h00;      memory[8419] <=  8'h00;      memory[8420] <=  8'h00;      memory[8421] <=  8'h00;      memory[8422] <=  8'h00;      memory[8423] <=  8'h00;      memory[8424] <=  8'h00;      memory[8425] <=  8'h00;      memory[8426] <=  8'h00;      memory[8427] <=  8'h00;      memory[8428] <=  8'h00;      memory[8429] <=  8'h00;      memory[8430] <=  8'h00;      memory[8431] <=  8'h00;      memory[8432] <=  8'h00;      memory[8433] <=  8'h00;      memory[8434] <=  8'h00;      memory[8435] <=  8'h00;      memory[8436] <=  8'h00;      memory[8437] <=  8'h00;      memory[8438] <=  8'h00;      memory[8439] <=  8'h00;      memory[8440] <=  8'h00;      memory[8441] <=  8'h00;      memory[8442] <=  8'h00;      memory[8443] <=  8'h00;      memory[8444] <=  8'h00;      memory[8445] <=  8'h00;      memory[8446] <=  8'h00;      memory[8447] <=  8'h00;      memory[8448] <=  8'h00;      memory[8449] <=  8'h00;      memory[8450] <=  8'h00;      memory[8451] <=  8'h00;      memory[8452] <=  8'h00;      memory[8453] <=  8'h00;      memory[8454] <=  8'h00;      memory[8455] <=  8'h00;      memory[8456] <=  8'h00;      memory[8457] <=  8'h00;      memory[8458] <=  8'h00;      memory[8459] <=  8'h00;      memory[8460] <=  8'h00;      memory[8461] <=  8'h00;      memory[8462] <=  8'h00;      memory[8463] <=  8'h00;      memory[8464] <=  8'h00;      memory[8465] <=  8'h00;      memory[8466] <=  8'h00;      memory[8467] <=  8'h00;      memory[8468] <=  8'h00;      memory[8469] <=  8'h00;      memory[8470] <=  8'h00;      memory[8471] <=  8'h00;      memory[8472] <=  8'h00;      memory[8473] <=  8'h00;      memory[8474] <=  8'h00;      memory[8475] <=  8'h00;      memory[8476] <=  8'h00;      memory[8477] <=  8'h00;      memory[8478] <=  8'h00;      memory[8479] <=  8'h00;      memory[8480] <=  8'h00;      memory[8481] <=  8'h00;      memory[8482] <=  8'h00;      memory[8483] <=  8'h00;      memory[8484] <=  8'h00;      memory[8485] <=  8'h00;      memory[8486] <=  8'h00;      memory[8487] <=  8'h00;      memory[8488] <=  8'h00;      memory[8489] <=  8'h00;      memory[8490] <=  8'h00;      memory[8491] <=  8'h00;      memory[8492] <=  8'h00;      memory[8493] <=  8'h00;      memory[8494] <=  8'h00;      memory[8495] <=  8'h00;      memory[8496] <=  8'h00;      memory[8497] <=  8'h00;      memory[8498] <=  8'h00;      memory[8499] <=  8'h00;      memory[8500] <=  8'h00;      memory[8501] <=  8'h00;      memory[8502] <=  8'h00;      memory[8503] <=  8'h00;      memory[8504] <=  8'h00;      memory[8505] <=  8'h00;      memory[8506] <=  8'h00;      memory[8507] <=  8'h00;      memory[8508] <=  8'h00;      memory[8509] <=  8'h00;      memory[8510] <=  8'h00;      memory[8511] <=  8'h00;      memory[8512] <=  8'h00;      memory[8513] <=  8'h00;      memory[8514] <=  8'h00;      memory[8515] <=  8'h00;      memory[8516] <=  8'h00;      memory[8517] <=  8'h00;      memory[8518] <=  8'h00;      memory[8519] <=  8'h00;      memory[8520] <=  8'h00;      memory[8521] <=  8'h00;      memory[8522] <=  8'h00;      memory[8523] <=  8'h00;      memory[8524] <=  8'h00;      memory[8525] <=  8'h00;      memory[8526] <=  8'h00;      memory[8527] <=  8'h00;      memory[8528] <=  8'h00;      memory[8529] <=  8'h00;      memory[8530] <=  8'h00;      memory[8531] <=  8'h00;      memory[8532] <=  8'h00;      memory[8533] <=  8'h00;      memory[8534] <=  8'h00;      memory[8535] <=  8'h00;      memory[8536] <=  8'h00;      memory[8537] <=  8'h00;      memory[8538] <=  8'h00;      memory[8539] <=  8'h00;      memory[8540] <=  8'h00;      memory[8541] <=  8'h00;      memory[8542] <=  8'h00;      memory[8543] <=  8'h00;      memory[8544] <=  8'h00;      memory[8545] <=  8'h00;      memory[8546] <=  8'h00;      memory[8547] <=  8'h00;      memory[8548] <=  8'h00;      memory[8549] <=  8'h00;      memory[8550] <=  8'h00;      memory[8551] <=  8'h00;      memory[8552] <=  8'h00;      memory[8553] <=  8'h00;      memory[8554] <=  8'h00;      memory[8555] <=  8'h00;      memory[8556] <=  8'h00;      memory[8557] <=  8'h00;      memory[8558] <=  8'h00;      memory[8559] <=  8'h00;      memory[8560] <=  8'h00;      memory[8561] <=  8'h00;      memory[8562] <=  8'h00;      memory[8563] <=  8'h00;      memory[8564] <=  8'h00;      memory[8565] <=  8'h00;      memory[8566] <=  8'h00;      memory[8567] <=  8'h00;      memory[8568] <=  8'h00;      memory[8569] <=  8'h00;      memory[8570] <=  8'h00;      memory[8571] <=  8'h00;      memory[8572] <=  8'h00;      memory[8573] <=  8'h00;      memory[8574] <=  8'h00;      memory[8575] <=  8'h00;      memory[8576] <=  8'h00;      memory[8577] <=  8'h00;      memory[8578] <=  8'h00;      memory[8579] <=  8'h00;      memory[8580] <=  8'h00;      memory[8581] <=  8'h00;      memory[8582] <=  8'h00;      memory[8583] <=  8'h00;      memory[8584] <=  8'h00;      memory[8585] <=  8'h00;      memory[8586] <=  8'h00;      memory[8587] <=  8'h00;      memory[8588] <=  8'h00;      memory[8589] <=  8'h00;      memory[8590] <=  8'h00;      memory[8591] <=  8'h00;      memory[8592] <=  8'h00;      memory[8593] <=  8'h00;      memory[8594] <=  8'h00;      memory[8595] <=  8'h00;      memory[8596] <=  8'h00;      memory[8597] <=  8'h00;      memory[8598] <=  8'h00;      memory[8599] <=  8'h00;      memory[8600] <=  8'h00;      memory[8601] <=  8'h00;      memory[8602] <=  8'h00;      memory[8603] <=  8'h00;      memory[8604] <=  8'h00;      memory[8605] <=  8'h00;      memory[8606] <=  8'h00;      memory[8607] <=  8'h00;      memory[8608] <=  8'h00;      memory[8609] <=  8'h00;      memory[8610] <=  8'h00;      memory[8611] <=  8'h00;      memory[8612] <=  8'h00;      memory[8613] <=  8'h00;      memory[8614] <=  8'h00;      memory[8615] <=  8'h00;      memory[8616] <=  8'h00;      memory[8617] <=  8'h00;      memory[8618] <=  8'h00;      memory[8619] <=  8'h00;      memory[8620] <=  8'h00;      memory[8621] <=  8'h00;      memory[8622] <=  8'h00;      memory[8623] <=  8'h00;      memory[8624] <=  8'h00;      memory[8625] <=  8'h00;      memory[8626] <=  8'h00;      memory[8627] <=  8'h00;      memory[8628] <=  8'h00;      memory[8629] <=  8'h00;      memory[8630] <=  8'h00;      memory[8631] <=  8'h00;      memory[8632] <=  8'h00;      memory[8633] <=  8'h00;      memory[8634] <=  8'h00;      memory[8635] <=  8'h00;      memory[8636] <=  8'h00;      memory[8637] <=  8'h00;      memory[8638] <=  8'h00;      memory[8639] <=  8'h00;      memory[8640] <=  8'h00;      memory[8641] <=  8'h00;      memory[8642] <=  8'h00;      memory[8643] <=  8'h00;      memory[8644] <=  8'h00;      memory[8645] <=  8'h00;      memory[8646] <=  8'h00;      memory[8647] <=  8'h00;      memory[8648] <=  8'h00;      memory[8649] <=  8'h00;      memory[8650] <=  8'h00;      memory[8651] <=  8'h00;      memory[8652] <=  8'h00;      memory[8653] <=  8'h00;      memory[8654] <=  8'h00;      memory[8655] <=  8'h00;      memory[8656] <=  8'h00;      memory[8657] <=  8'h00;      memory[8658] <=  8'h00;      memory[8659] <=  8'h00;      memory[8660] <=  8'h00;      memory[8661] <=  8'h00;      memory[8662] <=  8'h00;      memory[8663] <=  8'h00;      memory[8664] <=  8'h00;      memory[8665] <=  8'h00;      memory[8666] <=  8'h00;      memory[8667] <=  8'h00;      memory[8668] <=  8'h00;      memory[8669] <=  8'h00;      memory[8670] <=  8'h00;      memory[8671] <=  8'h00;      memory[8672] <=  8'h00;      memory[8673] <=  8'h00;      memory[8674] <=  8'h00;      memory[8675] <=  8'h00;      memory[8676] <=  8'h00;      memory[8677] <=  8'h00;      memory[8678] <=  8'h00;      memory[8679] <=  8'h00;      memory[8680] <=  8'h00;      memory[8681] <=  8'h00;      memory[8682] <=  8'h00;      memory[8683] <=  8'h00;      memory[8684] <=  8'h00;      memory[8685] <=  8'h00;      memory[8686] <=  8'h00;      memory[8687] <=  8'h00;      memory[8688] <=  8'h00;      memory[8689] <=  8'h00;      memory[8690] <=  8'h00;      memory[8691] <=  8'h00;      memory[8692] <=  8'h00;      memory[8693] <=  8'h00;      memory[8694] <=  8'h00;      memory[8695] <=  8'h00;      memory[8696] <=  8'h00;      memory[8697] <=  8'h00;      memory[8698] <=  8'h00;      memory[8699] <=  8'h00;      memory[8700] <=  8'h00;      memory[8701] <=  8'h00;      memory[8702] <=  8'h00;      memory[8703] <=  8'h00;      memory[8704] <=  8'h00;      memory[8705] <=  8'h00;      memory[8706] <=  8'h00;      memory[8707] <=  8'h00;      memory[8708] <=  8'h00;      memory[8709] <=  8'h00;      memory[8710] <=  8'h00;      memory[8711] <=  8'h00;      memory[8712] <=  8'h00;      memory[8713] <=  8'h00;      memory[8714] <=  8'h00;      memory[8715] <=  8'h00;      memory[8716] <=  8'h00;      memory[8717] <=  8'h00;      memory[8718] <=  8'h00;      memory[8719] <=  8'h00;      memory[8720] <=  8'h00;      memory[8721] <=  8'h00;      memory[8722] <=  8'h00;      memory[8723] <=  8'h00;      memory[8724] <=  8'h00;      memory[8725] <=  8'h00;      memory[8726] <=  8'h00;      memory[8727] <=  8'h00;      memory[8728] <=  8'h00;      memory[8729] <=  8'h00;      memory[8730] <=  8'h00;      memory[8731] <=  8'h00;      memory[8732] <=  8'h00;      memory[8733] <=  8'h00;      memory[8734] <=  8'h00;      memory[8735] <=  8'h00;      memory[8736] <=  8'h00;      memory[8737] <=  8'h00;      memory[8738] <=  8'h00;      memory[8739] <=  8'h00;      memory[8740] <=  8'h00;      memory[8741] <=  8'h00;      memory[8742] <=  8'h00;      memory[8743] <=  8'h00;      memory[8744] <=  8'h00;      memory[8745] <=  8'h00;      memory[8746] <=  8'h00;      memory[8747] <=  8'h00;      memory[8748] <=  8'h00;      memory[8749] <=  8'h00;      memory[8750] <=  8'h00;      memory[8751] <=  8'h00;      memory[8752] <=  8'h00;      memory[8753] <=  8'h00;      memory[8754] <=  8'h00;      memory[8755] <=  8'h00;      memory[8756] <=  8'h00;      memory[8757] <=  8'h00;      memory[8758] <=  8'h00;      memory[8759] <=  8'h00;      memory[8760] <=  8'h00;      memory[8761] <=  8'h00;      memory[8762] <=  8'h00;      memory[8763] <=  8'h00;      memory[8764] <=  8'h00;      memory[8765] <=  8'h00;      memory[8766] <=  8'h00;      memory[8767] <=  8'h00;      memory[8768] <=  8'h00;      memory[8769] <=  8'h00;      memory[8770] <=  8'h00;      memory[8771] <=  8'h00;      memory[8772] <=  8'h00;      memory[8773] <=  8'h00;      memory[8774] <=  8'h00;      memory[8775] <=  8'h00;      memory[8776] <=  8'h00;      memory[8777] <=  8'h00;      memory[8778] <=  8'h00;      memory[8779] <=  8'h00;      memory[8780] <=  8'h00;      memory[8781] <=  8'h00;      memory[8782] <=  8'h00;      memory[8783] <=  8'h00;      memory[8784] <=  8'h00;      memory[8785] <=  8'h00;      memory[8786] <=  8'h00;      memory[8787] <=  8'h00;      memory[8788] <=  8'h00;      memory[8789] <=  8'h00;      memory[8790] <=  8'h00;      memory[8791] <=  8'h00;      memory[8792] <=  8'h00;      memory[8793] <=  8'h00;      memory[8794] <=  8'h00;      memory[8795] <=  8'h00;      memory[8796] <=  8'h00;      memory[8797] <=  8'h00;      memory[8798] <=  8'h00;      memory[8799] <=  8'h00;      memory[8800] <=  8'h00;      memory[8801] <=  8'h00;      memory[8802] <=  8'h00;      memory[8803] <=  8'h00;      memory[8804] <=  8'h00;      memory[8805] <=  8'h00;      memory[8806] <=  8'h00;      memory[8807] <=  8'h00;      memory[8808] <=  8'h00;      memory[8809] <=  8'h00;      memory[8810] <=  8'h00;      memory[8811] <=  8'h00;      memory[8812] <=  8'h00;      memory[8813] <=  8'h00;      memory[8814] <=  8'h00;      memory[8815] <=  8'h00;      memory[8816] <=  8'h00;      memory[8817] <=  8'h00;      memory[8818] <=  8'h00;      memory[8819] <=  8'h00;      memory[8820] <=  8'h00;      memory[8821] <=  8'h00;      memory[8822] <=  8'h00;      memory[8823] <=  8'h00;      memory[8824] <=  8'h00;      memory[8825] <=  8'h00;      memory[8826] <=  8'h00;      memory[8827] <=  8'h00;      memory[8828] <=  8'h00;      memory[8829] <=  8'h00;      memory[8830] <=  8'h00;      memory[8831] <=  8'h00;      memory[8832] <=  8'h00;      memory[8833] <=  8'h00;      memory[8834] <=  8'h00;      memory[8835] <=  8'h00;      memory[8836] <=  8'h00;      memory[8837] <=  8'h00;      memory[8838] <=  8'h00;      memory[8839] <=  8'h00;      memory[8840] <=  8'h00;      memory[8841] <=  8'h00;      memory[8842] <=  8'h00;      memory[8843] <=  8'h00;      memory[8844] <=  8'h00;      memory[8845] <=  8'h00;      memory[8846] <=  8'h00;      memory[8847] <=  8'h00;      memory[8848] <=  8'h00;      memory[8849] <=  8'h00;      memory[8850] <=  8'h00;      memory[8851] <=  8'h00;      memory[8852] <=  8'h00;      memory[8853] <=  8'h00;      memory[8854] <=  8'h00;      memory[8855] <=  8'h00;      memory[8856] <=  8'h00;      memory[8857] <=  8'h00;      memory[8858] <=  8'h00;      memory[8859] <=  8'h00;      memory[8860] <=  8'h00;      memory[8861] <=  8'h00;      memory[8862] <=  8'h00;      memory[8863] <=  8'h00;      memory[8864] <=  8'h00;      memory[8865] <=  8'h00;      memory[8866] <=  8'h00;      memory[8867] <=  8'h00;      memory[8868] <=  8'h00;      memory[8869] <=  8'h00;      memory[8870] <=  8'h00;      memory[8871] <=  8'h00;      memory[8872] <=  8'h00;      memory[8873] <=  8'h00;      memory[8874] <=  8'h00;      memory[8875] <=  8'h00;      memory[8876] <=  8'h00;      memory[8877] <=  8'h00;      memory[8878] <=  8'h00;      memory[8879] <=  8'h00;      memory[8880] <=  8'h00;      memory[8881] <=  8'h00;      memory[8882] <=  8'h00;      memory[8883] <=  8'h00;      memory[8884] <=  8'h00;      memory[8885] <=  8'h00;      memory[8886] <=  8'h00;      memory[8887] <=  8'h00;      memory[8888] <=  8'h00;      memory[8889] <=  8'h00;      memory[8890] <=  8'h00;      memory[8891] <=  8'h00;      memory[8892] <=  8'h00;      memory[8893] <=  8'h00;      memory[8894] <=  8'h00;      memory[8895] <=  8'h00;      memory[8896] <=  8'h00;      memory[8897] <=  8'h00;      memory[8898] <=  8'h00;      memory[8899] <=  8'h00;      memory[8900] <=  8'h00;      memory[8901] <=  8'h00;      memory[8902] <=  8'h00;      memory[8903] <=  8'h00;      memory[8904] <=  8'h00;      memory[8905] <=  8'h00;      memory[8906] <=  8'h00;      memory[8907] <=  8'h00;      memory[8908] <=  8'h00;      memory[8909] <=  8'h00;      memory[8910] <=  8'h00;      memory[8911] <=  8'h00;      memory[8912] <=  8'h00;      memory[8913] <=  8'h00;      memory[8914] <=  8'h00;      memory[8915] <=  8'h00;      memory[8916] <=  8'h00;      memory[8917] <=  8'h00;      memory[8918] <=  8'h00;      memory[8919] <=  8'h00;      memory[8920] <=  8'h00;      memory[8921] <=  8'h00;      memory[8922] <=  8'h00;      memory[8923] <=  8'h00;      memory[8924] <=  8'h00;      memory[8925] <=  8'h00;      memory[8926] <=  8'h00;      memory[8927] <=  8'h00;      memory[8928] <=  8'h00;      memory[8929] <=  8'h00;      memory[8930] <=  8'h00;      memory[8931] <=  8'h00;      memory[8932] <=  8'h00;      memory[8933] <=  8'h00;      memory[8934] <=  8'h00;      memory[8935] <=  8'h00;      memory[8936] <=  8'h00;      memory[8937] <=  8'h00;      memory[8938] <=  8'h00;      memory[8939] <=  8'h00;      memory[8940] <=  8'h00;      memory[8941] <=  8'h00;      memory[8942] <=  8'h00;      memory[8943] <=  8'h00;      memory[8944] <=  8'h00;      memory[8945] <=  8'h00;      memory[8946] <=  8'h00;      memory[8947] <=  8'h00;      memory[8948] <=  8'h00;      memory[8949] <=  8'h00;      memory[8950] <=  8'h00;      memory[8951] <=  8'h00;      memory[8952] <=  8'h00;      memory[8953] <=  8'h00;      memory[8954] <=  8'h00;      memory[8955] <=  8'h00;      memory[8956] <=  8'h00;      memory[8957] <=  8'h00;      memory[8958] <=  8'h00;      memory[8959] <=  8'h00;      memory[8960] <=  8'h00;      memory[8961] <=  8'h00;      memory[8962] <=  8'h00;      memory[8963] <=  8'h00;      memory[8964] <=  8'h00;      memory[8965] <=  8'h00;      memory[8966] <=  8'h00;      memory[8967] <=  8'h00;      memory[8968] <=  8'h00;      memory[8969] <=  8'h00;      memory[8970] <=  8'h00;      memory[8971] <=  8'h00;      memory[8972] <=  8'h00;      memory[8973] <=  8'h00;      memory[8974] <=  8'h00;      memory[8975] <=  8'h00;      memory[8976] <=  8'h00;      memory[8977] <=  8'h00;      memory[8978] <=  8'h00;      memory[8979] <=  8'h00;      memory[8980] <=  8'h00;      memory[8981] <=  8'h00;      memory[8982] <=  8'h00;      memory[8983] <=  8'h00;      memory[8984] <=  8'h00;      memory[8985] <=  8'h00;      memory[8986] <=  8'h00;      memory[8987] <=  8'h00;      memory[8988] <=  8'h00;      memory[8989] <=  8'h00;      memory[8990] <=  8'h00;      memory[8991] <=  8'h00;      memory[8992] <=  8'h00;      memory[8993] <=  8'h00;      memory[8994] <=  8'h00;      memory[8995] <=  8'h00;      memory[8996] <=  8'h00;      memory[8997] <=  8'h00;      memory[8998] <=  8'h00;      memory[8999] <=  8'h00;      memory[9000] <=  8'h00;      memory[9001] <=  8'h00;      memory[9002] <=  8'h00;      memory[9003] <=  8'h00;      memory[9004] <=  8'h00;      memory[9005] <=  8'h00;      memory[9006] <=  8'h00;      memory[9007] <=  8'h00;      memory[9008] <=  8'h00;      memory[9009] <=  8'h00;      memory[9010] <=  8'h00;      memory[9011] <=  8'h00;      memory[9012] <=  8'h00;      memory[9013] <=  8'h00;      memory[9014] <=  8'h00;      memory[9015] <=  8'h00;      memory[9016] <=  8'h00;      memory[9017] <=  8'h00;      memory[9018] <=  8'h00;      memory[9019] <=  8'h00;      memory[9020] <=  8'h00;      memory[9021] <=  8'h00;      memory[9022] <=  8'h00;      memory[9023] <=  8'h00;      memory[9024] <=  8'h00;      memory[9025] <=  8'h00;      memory[9026] <=  8'h00;      memory[9027] <=  8'h00;      memory[9028] <=  8'h00;      memory[9029] <=  8'h00;      memory[9030] <=  8'h00;      memory[9031] <=  8'h00;      memory[9032] <=  8'h00;      memory[9033] <=  8'h00;      memory[9034] <=  8'h00;      memory[9035] <=  8'h00;      memory[9036] <=  8'h00;      memory[9037] <=  8'h00;      memory[9038] <=  8'h00;      memory[9039] <=  8'h00;      memory[9040] <=  8'h00;      memory[9041] <=  8'h00;      memory[9042] <=  8'h00;      memory[9043] <=  8'h00;      memory[9044] <=  8'h00;      memory[9045] <=  8'h00;      memory[9046] <=  8'h00;      memory[9047] <=  8'h00;      memory[9048] <=  8'h00;      memory[9049] <=  8'h00;      memory[9050] <=  8'h00;      memory[9051] <=  8'h00;      memory[9052] <=  8'h00;      memory[9053] <=  8'h00;      memory[9054] <=  8'h00;      memory[9055] <=  8'h00;      memory[9056] <=  8'h00;      memory[9057] <=  8'h00;      memory[9058] <=  8'h00;      memory[9059] <=  8'h00;      memory[9060] <=  8'h00;      memory[9061] <=  8'h00;      memory[9062] <=  8'h00;      memory[9063] <=  8'h00;      memory[9064] <=  8'h00;      memory[9065] <=  8'h00;      memory[9066] <=  8'h00;      memory[9067] <=  8'h00;      memory[9068] <=  8'h00;      memory[9069] <=  8'h00;      memory[9070] <=  8'h00;      memory[9071] <=  8'h00;      memory[9072] <=  8'h00;      memory[9073] <=  8'h00;      memory[9074] <=  8'h00;      memory[9075] <=  8'h00;      memory[9076] <=  8'h00;      memory[9077] <=  8'h00;      memory[9078] <=  8'h00;      memory[9079] <=  8'h00;      memory[9080] <=  8'h00;      memory[9081] <=  8'h00;      memory[9082] <=  8'h00;      memory[9083] <=  8'h00;      memory[9084] <=  8'h00;      memory[9085] <=  8'h00;      memory[9086] <=  8'h00;      memory[9087] <=  8'h00;      memory[9088] <=  8'h00;      memory[9089] <=  8'h00;      memory[9090] <=  8'h00;      memory[9091] <=  8'h00;      memory[9092] <=  8'h00;      memory[9093] <=  8'h00;      memory[9094] <=  8'h00;      memory[9095] <=  8'h00;      memory[9096] <=  8'h00;      memory[9097] <=  8'h00;      memory[9098] <=  8'h00;      memory[9099] <=  8'h00;      memory[9100] <=  8'h00;      memory[9101] <=  8'h00;      memory[9102] <=  8'h00;      memory[9103] <=  8'h00;      memory[9104] <=  8'h00;      memory[9105] <=  8'h00;      memory[9106] <=  8'h00;      memory[9107] <=  8'h00;      memory[9108] <=  8'h00;      memory[9109] <=  8'h00;      memory[9110] <=  8'h00;      memory[9111] <=  8'h00;      memory[9112] <=  8'h00;      memory[9113] <=  8'h00;      memory[9114] <=  8'h00;      memory[9115] <=  8'h00;      memory[9116] <=  8'h00;      memory[9117] <=  8'h00;      memory[9118] <=  8'h00;      memory[9119] <=  8'h00;      memory[9120] <=  8'h00;      memory[9121] <=  8'h00;      memory[9122] <=  8'h00;      memory[9123] <=  8'h00;      memory[9124] <=  8'h00;      memory[9125] <=  8'h00;      memory[9126] <=  8'h00;      memory[9127] <=  8'h00;      memory[9128] <=  8'h00;      memory[9129] <=  8'h00;      memory[9130] <=  8'h00;      memory[9131] <=  8'h00;      memory[9132] <=  8'h00;      memory[9133] <=  8'h00;      memory[9134] <=  8'h00;      memory[9135] <=  8'h00;      memory[9136] <=  8'h00;      memory[9137] <=  8'h00;      memory[9138] <=  8'h00;      memory[9139] <=  8'h00;      memory[9140] <=  8'h00;      memory[9141] <=  8'h00;      memory[9142] <=  8'h00;      memory[9143] <=  8'h00;      memory[9144] <=  8'h00;      memory[9145] <=  8'h00;      memory[9146] <=  8'h00;      memory[9147] <=  8'h00;      memory[9148] <=  8'h00;      memory[9149] <=  8'h00;      memory[9150] <=  8'h00;      memory[9151] <=  8'h00;      memory[9152] <=  8'h00;      memory[9153] <=  8'h00;      memory[9154] <=  8'h00;      memory[9155] <=  8'h00;      memory[9156] <=  8'h00;      memory[9157] <=  8'h00;      memory[9158] <=  8'h00;      memory[9159] <=  8'h00;      memory[9160] <=  8'h00;      memory[9161] <=  8'h00;      memory[9162] <=  8'h00;      memory[9163] <=  8'h00;      memory[9164] <=  8'h00;      memory[9165] <=  8'h00;      memory[9166] <=  8'h00;      memory[9167] <=  8'h00;      memory[9168] <=  8'h00;      memory[9169] <=  8'h00;      memory[9170] <=  8'h00;      memory[9171] <=  8'h00;      memory[9172] <=  8'h00;      memory[9173] <=  8'h00;      memory[9174] <=  8'h00;      memory[9175] <=  8'h00;      memory[9176] <=  8'h00;      memory[9177] <=  8'h00;      memory[9178] <=  8'h00;      memory[9179] <=  8'h00;      memory[9180] <=  8'h00;      memory[9181] <=  8'h00;      memory[9182] <=  8'h00;      memory[9183] <=  8'h00;      memory[9184] <=  8'h00;      memory[9185] <=  8'h00;      memory[9186] <=  8'h00;      memory[9187] <=  8'h00;      memory[9188] <=  8'h00;      memory[9189] <=  8'h00;      memory[9190] <=  8'h00;      memory[9191] <=  8'h00;      memory[9192] <=  8'h00;      memory[9193] <=  8'h00;      memory[9194] <=  8'h00;      memory[9195] <=  8'h00;      memory[9196] <=  8'h00;      memory[9197] <=  8'h00;      memory[9198] <=  8'h00;      memory[9199] <=  8'h00;      memory[9200] <=  8'h00;      memory[9201] <=  8'h00;      memory[9202] <=  8'h00;      memory[9203] <=  8'h00;      memory[9204] <=  8'h00;      memory[9205] <=  8'h00;      memory[9206] <=  8'h00;      memory[9207] <=  8'h00;      memory[9208] <=  8'h00;      memory[9209] <=  8'h00;      memory[9210] <=  8'h00;      memory[9211] <=  8'h00;      memory[9212] <=  8'h00;      memory[9213] <=  8'h00;      memory[9214] <=  8'h00;      memory[9215] <=  8'h00;      memory[9216] <=  8'h00;      memory[9217] <=  8'h00;      memory[9218] <=  8'h00;      memory[9219] <=  8'h00;      memory[9220] <=  8'h00;      memory[9221] <=  8'h00;      memory[9222] <=  8'h00;      memory[9223] <=  8'h00;      memory[9224] <=  8'h00;      memory[9225] <=  8'h00;      memory[9226] <=  8'h00;      memory[9227] <=  8'h00;      memory[9228] <=  8'h00;      memory[9229] <=  8'h00;      memory[9230] <=  8'h00;      memory[9231] <=  8'h00;      memory[9232] <=  8'h00;      memory[9233] <=  8'h00;      memory[9234] <=  8'h00;      memory[9235] <=  8'h00;      memory[9236] <=  8'h00;      memory[9237] <=  8'h00;      memory[9238] <=  8'h00;      memory[9239] <=  8'h00;      memory[9240] <=  8'h00;      memory[9241] <=  8'h00;      memory[9242] <=  8'h00;      memory[9243] <=  8'h00;      memory[9244] <=  8'h00;      memory[9245] <=  8'h00;      memory[9246] <=  8'h00;      memory[9247] <=  8'h00;      memory[9248] <=  8'h00;      memory[9249] <=  8'h00;      memory[9250] <=  8'h00;      memory[9251] <=  8'h00;      memory[9252] <=  8'h00;      memory[9253] <=  8'h00;      memory[9254] <=  8'h00;      memory[9255] <=  8'h00;      memory[9256] <=  8'h00;      memory[9257] <=  8'h00;      memory[9258] <=  8'h00;      memory[9259] <=  8'h00;      memory[9260] <=  8'h00;      memory[9261] <=  8'h00;      memory[9262] <=  8'h00;      memory[9263] <=  8'h00;      memory[9264] <=  8'h00;      memory[9265] <=  8'h00;      memory[9266] <=  8'h00;      memory[9267] <=  8'h00;      memory[9268] <=  8'h00;      memory[9269] <=  8'h00;      memory[9270] <=  8'h00;      memory[9271] <=  8'h00;      memory[9272] <=  8'h00;      memory[9273] <=  8'h00;      memory[9274] <=  8'h00;      memory[9275] <=  8'h00;      memory[9276] <=  8'h00;      memory[9277] <=  8'h00;      memory[9278] <=  8'h00;      memory[9279] <=  8'h00;      memory[9280] <=  8'h00;      memory[9281] <=  8'h00;      memory[9282] <=  8'h00;      memory[9283] <=  8'h00;      memory[9284] <=  8'h00;      memory[9285] <=  8'h00;      memory[9286] <=  8'h00;      memory[9287] <=  8'h00;      memory[9288] <=  8'h00;      memory[9289] <=  8'h00;      memory[9290] <=  8'h00;      memory[9291] <=  8'h00;      memory[9292] <=  8'h00;      memory[9293] <=  8'h00;      memory[9294] <=  8'h00;      memory[9295] <=  8'h00;      memory[9296] <=  8'h00;      memory[9297] <=  8'h00;      memory[9298] <=  8'h00;      memory[9299] <=  8'h00;      memory[9300] <=  8'h00;      memory[9301] <=  8'h00;      memory[9302] <=  8'h00;      memory[9303] <=  8'h00;      memory[9304] <=  8'h00;      memory[9305] <=  8'h00;      memory[9306] <=  8'h00;      memory[9307] <=  8'h00;      memory[9308] <=  8'h00;      memory[9309] <=  8'h00;      memory[9310] <=  8'h00;      memory[9311] <=  8'h00;      memory[9312] <=  8'h00;      memory[9313] <=  8'h00;      memory[9314] <=  8'h00;      memory[9315] <=  8'h00;      memory[9316] <=  8'h00;      memory[9317] <=  8'h00;      memory[9318] <=  8'h00;      memory[9319] <=  8'h00;      memory[9320] <=  8'h00;      memory[9321] <=  8'h00;      memory[9322] <=  8'h00;      memory[9323] <=  8'h00;      memory[9324] <=  8'h00;      memory[9325] <=  8'h00;      memory[9326] <=  8'h00;      memory[9327] <=  8'h00;      memory[9328] <=  8'h00;      memory[9329] <=  8'h00;      memory[9330] <=  8'h00;      memory[9331] <=  8'h00;      memory[9332] <=  8'h00;      memory[9333] <=  8'h00;      memory[9334] <=  8'h00;      memory[9335] <=  8'h00;      memory[9336] <=  8'h00;      memory[9337] <=  8'h00;      memory[9338] <=  8'h00;      memory[9339] <=  8'h00;      memory[9340] <=  8'h00;      memory[9341] <=  8'h00;      memory[9342] <=  8'h00;      memory[9343] <=  8'h00;      memory[9344] <=  8'h00;      memory[9345] <=  8'h00;      memory[9346] <=  8'h00;      memory[9347] <=  8'h00;      memory[9348] <=  8'h00;      memory[9349] <=  8'h00;      memory[9350] <=  8'h00;      memory[9351] <=  8'h00;      memory[9352] <=  8'h00;      memory[9353] <=  8'h00;      memory[9354] <=  8'h00;      memory[9355] <=  8'h00;      memory[9356] <=  8'h00;      memory[9357] <=  8'h00;      memory[9358] <=  8'h00;      memory[9359] <=  8'h00;      memory[9360] <=  8'h00;      memory[9361] <=  8'h00;      memory[9362] <=  8'h00;      memory[9363] <=  8'h00;      memory[9364] <=  8'h00;      memory[9365] <=  8'h00;      memory[9366] <=  8'h00;      memory[9367] <=  8'h00;      memory[9368] <=  8'h00;      memory[9369] <=  8'h00;      memory[9370] <=  8'h00;      memory[9371] <=  8'h00;      memory[9372] <=  8'h00;      memory[9373] <=  8'h00;      memory[9374] <=  8'h00;      memory[9375] <=  8'h00;      memory[9376] <=  8'h00;      memory[9377] <=  8'h00;      memory[9378] <=  8'h00;      memory[9379] <=  8'h00;      memory[9380] <=  8'h00;      memory[9381] <=  8'h00;      memory[9382] <=  8'h00;      memory[9383] <=  8'h00;      memory[9384] <=  8'h00;      memory[9385] <=  8'h00;      memory[9386] <=  8'h00;      memory[9387] <=  8'h00;      memory[9388] <=  8'h00;      memory[9389] <=  8'h00;      memory[9390] <=  8'h00;      memory[9391] <=  8'h00;      memory[9392] <=  8'h00;      memory[9393] <=  8'h00;      memory[9394] <=  8'h00;      memory[9395] <=  8'h00;      memory[9396] <=  8'h00;      memory[9397] <=  8'h00;      memory[9398] <=  8'h00;      memory[9399] <=  8'h00;      memory[9400] <=  8'h00;      memory[9401] <=  8'h00;      memory[9402] <=  8'h00;      memory[9403] <=  8'h00;      memory[9404] <=  8'h00;      memory[9405] <=  8'h00;      memory[9406] <=  8'h00;      memory[9407] <=  8'h00;      memory[9408] <=  8'h00;      memory[9409] <=  8'h00;      memory[9410] <=  8'h00;      memory[9411] <=  8'h00;      memory[9412] <=  8'h00;      memory[9413] <=  8'h00;      memory[9414] <=  8'h00;      memory[9415] <=  8'h00;      memory[9416] <=  8'h00;      memory[9417] <=  8'h00;      memory[9418] <=  8'h00;      memory[9419] <=  8'h00;      memory[9420] <=  8'h00;      memory[9421] <=  8'h00;      memory[9422] <=  8'h00;      memory[9423] <=  8'h00;      memory[9424] <=  8'h00;      memory[9425] <=  8'h00;      memory[9426] <=  8'h00;      memory[9427] <=  8'h00;      memory[9428] <=  8'h00;      memory[9429] <=  8'h00;      memory[9430] <=  8'h00;      memory[9431] <=  8'h00;      memory[9432] <=  8'h00;      memory[9433] <=  8'h00;      memory[9434] <=  8'h00;      memory[9435] <=  8'h00;      memory[9436] <=  8'h00;      memory[9437] <=  8'h00;      memory[9438] <=  8'h00;      memory[9439] <=  8'h00;      memory[9440] <=  8'h00;      memory[9441] <=  8'h00;      memory[9442] <=  8'h00;      memory[9443] <=  8'h00;      memory[9444] <=  8'h00;      memory[9445] <=  8'h00;      memory[9446] <=  8'h00;      memory[9447] <=  8'h00;      memory[9448] <=  8'h00;      memory[9449] <=  8'h00;      memory[9450] <=  8'h00;      memory[9451] <=  8'h00;      memory[9452] <=  8'h00;      memory[9453] <=  8'h00;      memory[9454] <=  8'h00;      memory[9455] <=  8'h00;      memory[9456] <=  8'h00;      memory[9457] <=  8'h00;      memory[9458] <=  8'h00;      memory[9459] <=  8'h00;      memory[9460] <=  8'h00;      memory[9461] <=  8'h00;      memory[9462] <=  8'h00;      memory[9463] <=  8'h00;      memory[9464] <=  8'h00;      memory[9465] <=  8'h00;      memory[9466] <=  8'h00;      memory[9467] <=  8'h00;      memory[9468] <=  8'h00;      memory[9469] <=  8'h00;      memory[9470] <=  8'h00;      memory[9471] <=  8'h00;      memory[9472] <=  8'h00;      memory[9473] <=  8'h00;      memory[9474] <=  8'h00;      memory[9475] <=  8'h00;      memory[9476] <=  8'h00;      memory[9477] <=  8'h00;      memory[9478] <=  8'h00;      memory[9479] <=  8'h00;      memory[9480] <=  8'h00;      memory[9481] <=  8'h00;      memory[9482] <=  8'h00;      memory[9483] <=  8'h00;      memory[9484] <=  8'h00;      memory[9485] <=  8'h00;      memory[9486] <=  8'h00;      memory[9487] <=  8'h00;      memory[9488] <=  8'h00;      memory[9489] <=  8'h00;      memory[9490] <=  8'h00;      memory[9491] <=  8'h00;      memory[9492] <=  8'h00;      memory[9493] <=  8'h00;      memory[9494] <=  8'h00;      memory[9495] <=  8'h00;      memory[9496] <=  8'h00;      memory[9497] <=  8'h00;      memory[9498] <=  8'h00;      memory[9499] <=  8'h00;      memory[9500] <=  8'h00;      memory[9501] <=  8'h00;      memory[9502] <=  8'h00;      memory[9503] <=  8'h00;      memory[9504] <=  8'h00;      memory[9505] <=  8'h00;      memory[9506] <=  8'h00;      memory[9507] <=  8'h00;      memory[9508] <=  8'h00;      memory[9509] <=  8'h00;      memory[9510] <=  8'h00;      memory[9511] <=  8'h00;      memory[9512] <=  8'h00;      memory[9513] <=  8'h00;      memory[9514] <=  8'h00;      memory[9515] <=  8'h00;      memory[9516] <=  8'h00;      memory[9517] <=  8'h00;      memory[9518] <=  8'h00;      memory[9519] <=  8'h00;      memory[9520] <=  8'h00;      memory[9521] <=  8'h00;      memory[9522] <=  8'h00;      memory[9523] <=  8'h00;      memory[9524] <=  8'h00;      memory[9525] <=  8'h00;      memory[9526] <=  8'h00;      memory[9527] <=  8'h00;      memory[9528] <=  8'h00;      memory[9529] <=  8'h00;      memory[9530] <=  8'h00;      memory[9531] <=  8'h00;      memory[9532] <=  8'h00;      memory[9533] <=  8'h00;      memory[9534] <=  8'h00;      memory[9535] <=  8'h00;      memory[9536] <=  8'h00;      memory[9537] <=  8'h00;      memory[9538] <=  8'h00;      memory[9539] <=  8'h00;      memory[9540] <=  8'h00;      memory[9541] <=  8'h00;      memory[9542] <=  8'h00;      memory[9543] <=  8'h00;      memory[9544] <=  8'h00;      memory[9545] <=  8'h00;      memory[9546] <=  8'h00;      memory[9547] <=  8'h00;      memory[9548] <=  8'h00;      memory[9549] <=  8'h00;      memory[9550] <=  8'h00;      memory[9551] <=  8'h00;      memory[9552] <=  8'h00;      memory[9553] <=  8'h00;      memory[9554] <=  8'h00;      memory[9555] <=  8'h00;      memory[9556] <=  8'h00;      memory[9557] <=  8'h00;      memory[9558] <=  8'h00;      memory[9559] <=  8'h00;      memory[9560] <=  8'h00;      memory[9561] <=  8'h00;      memory[9562] <=  8'h00;      memory[9563] <=  8'h00;      memory[9564] <=  8'h00;      memory[9565] <=  8'h00;      memory[9566] <=  8'h00;      memory[9567] <=  8'h00;      memory[9568] <=  8'h00;      memory[9569] <=  8'h00;      memory[9570] <=  8'h00;      memory[9571] <=  8'h00;      memory[9572] <=  8'h00;      memory[9573] <=  8'h00;      memory[9574] <=  8'h00;      memory[9575] <=  8'h00;      memory[9576] <=  8'h00;      memory[9577] <=  8'h00;      memory[9578] <=  8'h00;      memory[9579] <=  8'h00;      memory[9580] <=  8'h00;      memory[9581] <=  8'h00;      memory[9582] <=  8'h00;      memory[9583] <=  8'h00;      memory[9584] <=  8'h00;      memory[9585] <=  8'h00;      memory[9586] <=  8'h00;      memory[9587] <=  8'h00;      memory[9588] <=  8'h00;      memory[9589] <=  8'h00;      memory[9590] <=  8'h00;      memory[9591] <=  8'h00;      memory[9592] <=  8'h00;      memory[9593] <=  8'h00;      memory[9594] <=  8'h00;      memory[9595] <=  8'h00;      memory[9596] <=  8'h00;      memory[9597] <=  8'h00;      memory[9598] <=  8'h00;      memory[9599] <=  8'h00;      memory[9600] <=  8'h00;      memory[9601] <=  8'h00;      memory[9602] <=  8'h00;      memory[9603] <=  8'h00;      memory[9604] <=  8'h00;      memory[9605] <=  8'h00;      memory[9606] <=  8'h00;      memory[9607] <=  8'h00;      memory[9608] <=  8'h00;      memory[9609] <=  8'h00;      memory[9610] <=  8'h00;      memory[9611] <=  8'h00;      memory[9612] <=  8'h00;      memory[9613] <=  8'h00;      memory[9614] <=  8'h00;      memory[9615] <=  8'h00;      memory[9616] <=  8'h00;      memory[9617] <=  8'h00;      memory[9618] <=  8'h00;      memory[9619] <=  8'h00;      memory[9620] <=  8'h00;      memory[9621] <=  8'h00;      memory[9622] <=  8'h00;      memory[9623] <=  8'h00;      memory[9624] <=  8'h00;      memory[9625] <=  8'h00;      memory[9626] <=  8'h00;      memory[9627] <=  8'h00;      memory[9628] <=  8'h00;      memory[9629] <=  8'h00;      memory[9630] <=  8'h00;      memory[9631] <=  8'h00;      memory[9632] <=  8'h00;      memory[9633] <=  8'h00;      memory[9634] <=  8'h00;      memory[9635] <=  8'h00;      memory[9636] <=  8'h00;      memory[9637] <=  8'h00;      memory[9638] <=  8'h00;      memory[9639] <=  8'h00;      memory[9640] <=  8'h00;      memory[9641] <=  8'h00;      memory[9642] <=  8'h00;      memory[9643] <=  8'h00;      memory[9644] <=  8'h00;      memory[9645] <=  8'h00;      memory[9646] <=  8'h00;      memory[9647] <=  8'h00;      memory[9648] <=  8'h00;      memory[9649] <=  8'h00;      memory[9650] <=  8'h00;      memory[9651] <=  8'h00;      memory[9652] <=  8'h00;      memory[9653] <=  8'h00;      memory[9654] <=  8'h00;      memory[9655] <=  8'h00;      memory[9656] <=  8'h00;      memory[9657] <=  8'h00;      memory[9658] <=  8'h00;      memory[9659] <=  8'h00;      memory[9660] <=  8'h00;      memory[9661] <=  8'h00;      memory[9662] <=  8'h00;      memory[9663] <=  8'h00;      memory[9664] <=  8'h00;      memory[9665] <=  8'h00;      memory[9666] <=  8'h00;      memory[9667] <=  8'h00;      memory[9668] <=  8'h00;      memory[9669] <=  8'h00;      memory[9670] <=  8'h00;      memory[9671] <=  8'h00;      memory[9672] <=  8'h00;      memory[9673] <=  8'h00;      memory[9674] <=  8'h00;      memory[9675] <=  8'h00;      memory[9676] <=  8'h00;      memory[9677] <=  8'h00;      memory[9678] <=  8'h00;      memory[9679] <=  8'h00;      memory[9680] <=  8'h00;      memory[9681] <=  8'h00;      memory[9682] <=  8'h00;      memory[9683] <=  8'h00;      memory[9684] <=  8'h00;      memory[9685] <=  8'h00;      memory[9686] <=  8'h00;      memory[9687] <=  8'h00;      memory[9688] <=  8'h00;      memory[9689] <=  8'h00;      memory[9690] <=  8'h00;      memory[9691] <=  8'h00;      memory[9692] <=  8'h00;      memory[9693] <=  8'h00;      memory[9694] <=  8'h00;      memory[9695] <=  8'h00;      memory[9696] <=  8'h00;      memory[9697] <=  8'h00;      memory[9698] <=  8'h00;      memory[9699] <=  8'h00;      memory[9700] <=  8'h00;      memory[9701] <=  8'h00;      memory[9702] <=  8'h00;      memory[9703] <=  8'h00;      memory[9704] <=  8'h00;      memory[9705] <=  8'h00;      memory[9706] <=  8'h00;      memory[9707] <=  8'h00;      memory[9708] <=  8'h00;      memory[9709] <=  8'h00;      memory[9710] <=  8'h00;      memory[9711] <=  8'h00;      memory[9712] <=  8'h00;      memory[9713] <=  8'h00;      memory[9714] <=  8'h00;      memory[9715] <=  8'h00;      memory[9716] <=  8'h00;      memory[9717] <=  8'h00;      memory[9718] <=  8'h00;      memory[9719] <=  8'h00;      memory[9720] <=  8'h00;      memory[9721] <=  8'h00;      memory[9722] <=  8'h00;      memory[9723] <=  8'h00;      memory[9724] <=  8'h00;      memory[9725] <=  8'h00;      memory[9726] <=  8'h00;      memory[9727] <=  8'h00;      memory[9728] <=  8'h00;      memory[9729] <=  8'h00;      memory[9730] <=  8'h00;      memory[9731] <=  8'h00;      memory[9732] <=  8'h00;      memory[9733] <=  8'h00;      memory[9734] <=  8'h00;      memory[9735] <=  8'h00;      memory[9736] <=  8'h00;      memory[9737] <=  8'h00;      memory[9738] <=  8'h00;      memory[9739] <=  8'h00;      memory[9740] <=  8'h00;      memory[9741] <=  8'h00;      memory[9742] <=  8'h00;      memory[9743] <=  8'h00;      memory[9744] <=  8'h00;      memory[9745] <=  8'h00;      memory[9746] <=  8'h00;      memory[9747] <=  8'h00;      memory[9748] <=  8'h00;      memory[9749] <=  8'h00;      memory[9750] <=  8'h00;      memory[9751] <=  8'h00;      memory[9752] <=  8'h00;      memory[9753] <=  8'h00;      memory[9754] <=  8'h00;      memory[9755] <=  8'h00;      memory[9756] <=  8'h00;      memory[9757] <=  8'h00;      memory[9758] <=  8'h00;      memory[9759] <=  8'h00;      memory[9760] <=  8'h00;      memory[9761] <=  8'h00;      memory[9762] <=  8'h00;      memory[9763] <=  8'h00;      memory[9764] <=  8'h00;      memory[9765] <=  8'h00;      memory[9766] <=  8'h00;      memory[9767] <=  8'h00;      memory[9768] <=  8'h00;      memory[9769] <=  8'h00;      memory[9770] <=  8'h00;      memory[9771] <=  8'h00;      memory[9772] <=  8'h00;      memory[9773] <=  8'h00;      memory[9774] <=  8'h00;      memory[9775] <=  8'h00;      memory[9776] <=  8'h00;      memory[9777] <=  8'h00;      memory[9778] <=  8'h00;      memory[9779] <=  8'h00;      memory[9780] <=  8'h00;      memory[9781] <=  8'h00;      memory[9782] <=  8'h00;      memory[9783] <=  8'h00;      memory[9784] <=  8'h00;      memory[9785] <=  8'h00;      memory[9786] <=  8'h00;      memory[9787] <=  8'h00;      memory[9788] <=  8'h00;      memory[9789] <=  8'h00;      memory[9790] <=  8'h00;      memory[9791] <=  8'h00;      memory[9792] <=  8'h00;      memory[9793] <=  8'h00;      memory[9794] <=  8'h00;      memory[9795] <=  8'h00;      memory[9796] <=  8'h00;      memory[9797] <=  8'h00;      memory[9798] <=  8'h00;      memory[9799] <=  8'h00;      memory[9800] <=  8'h00;      memory[9801] <=  8'h00;      memory[9802] <=  8'h00;      memory[9803] <=  8'h00;      memory[9804] <=  8'h00;      memory[9805] <=  8'h00;      memory[9806] <=  8'h00;      memory[9807] <=  8'h00;      memory[9808] <=  8'h00;      memory[9809] <=  8'h00;      memory[9810] <=  8'h00;      memory[9811] <=  8'h00;      memory[9812] <=  8'h00;      memory[9813] <=  8'h00;      memory[9814] <=  8'h00;      memory[9815] <=  8'h00;      memory[9816] <=  8'h00;      memory[9817] <=  8'h00;      memory[9818] <=  8'h00;      memory[9819] <=  8'h00;      memory[9820] <=  8'h00;      memory[9821] <=  8'h00;      memory[9822] <=  8'h00;      memory[9823] <=  8'h00;      memory[9824] <=  8'h00;      memory[9825] <=  8'h00;      memory[9826] <=  8'h00;      memory[9827] <=  8'h00;      memory[9828] <=  8'h00;      memory[9829] <=  8'h00;      memory[9830] <=  8'h00;      memory[9831] <=  8'h00;      memory[9832] <=  8'h00;      memory[9833] <=  8'h00;      memory[9834] <=  8'h00;      memory[9835] <=  8'h00;      memory[9836] <=  8'h00;      memory[9837] <=  8'h00;      memory[9838] <=  8'h00;      memory[9839] <=  8'h00;      memory[9840] <=  8'h00;      memory[9841] <=  8'h00;      memory[9842] <=  8'h00;      memory[9843] <=  8'h00;      memory[9844] <=  8'h00;      memory[9845] <=  8'h00;      memory[9846] <=  8'h00;      memory[9847] <=  8'h00;      memory[9848] <=  8'h00;      memory[9849] <=  8'h00;      memory[9850] <=  8'h00;      memory[9851] <=  8'h00;      memory[9852] <=  8'h00;      memory[9853] <=  8'h00;      memory[9854] <=  8'h00;      memory[9855] <=  8'h00;      memory[9856] <=  8'h00;      memory[9857] <=  8'h00;      memory[9858] <=  8'h00;      memory[9859] <=  8'h00;      memory[9860] <=  8'h00;      memory[9861] <=  8'h00;      memory[9862] <=  8'h00;      memory[9863] <=  8'h00;      memory[9864] <=  8'h00;      memory[9865] <=  8'h00;      memory[9866] <=  8'h00;      memory[9867] <=  8'h00;      memory[9868] <=  8'h00;      memory[9869] <=  8'h00;      memory[9870] <=  8'h00;      memory[9871] <=  8'h00;      memory[9872] <=  8'h00;      memory[9873] <=  8'h00;      memory[9874] <=  8'h00;      memory[9875] <=  8'h00;      memory[9876] <=  8'h00;      memory[9877] <=  8'h00;      memory[9878] <=  8'h00;      memory[9879] <=  8'h00;      memory[9880] <=  8'h00;      memory[9881] <=  8'h00;      memory[9882] <=  8'h00;      memory[9883] <=  8'h00;      memory[9884] <=  8'h00;      memory[9885] <=  8'h00;      memory[9886] <=  8'h00;      memory[9887] <=  8'h00;      memory[9888] <=  8'h00;      memory[9889] <=  8'h00;      memory[9890] <=  8'h00;      memory[9891] <=  8'h00;      memory[9892] <=  8'h00;      memory[9893] <=  8'h00;      memory[9894] <=  8'h00;      memory[9895] <=  8'h00;      memory[9896] <=  8'h00;      memory[9897] <=  8'h00;      memory[9898] <=  8'h00;      memory[9899] <=  8'h00;      memory[9900] <=  8'h00;      memory[9901] <=  8'h00;      memory[9902] <=  8'h00;      memory[9903] <=  8'h00;      memory[9904] <=  8'h00;      memory[9905] <=  8'h00;      memory[9906] <=  8'h00;      memory[9907] <=  8'h00;      memory[9908] <=  8'h00;      memory[9909] <=  8'h00;      memory[9910] <=  8'h00;      memory[9911] <=  8'h00;      memory[9912] <=  8'h00;      memory[9913] <=  8'h00;      memory[9914] <=  8'h00;      memory[9915] <=  8'h00;      memory[9916] <=  8'h00;      memory[9917] <=  8'h00;      memory[9918] <=  8'h00;      memory[9919] <=  8'h00;      memory[9920] <=  8'h00;      memory[9921] <=  8'h00;      memory[9922] <=  8'h00;      memory[9923] <=  8'h00;      memory[9924] <=  8'h00;      memory[9925] <=  8'h00;      memory[9926] <=  8'h00;      memory[9927] <=  8'h00;      memory[9928] <=  8'h00;      memory[9929] <=  8'h00;      memory[9930] <=  8'h00;      memory[9931] <=  8'h00;      memory[9932] <=  8'h00;      memory[9933] <=  8'h00;      memory[9934] <=  8'h00;      memory[9935] <=  8'h00;      memory[9936] <=  8'h00;      memory[9937] <=  8'h00;      memory[9938] <=  8'h00;      memory[9939] <=  8'h00;      memory[9940] <=  8'h00;      memory[9941] <=  8'h00;      memory[9942] <=  8'h00;      memory[9943] <=  8'h00;      memory[9944] <=  8'h00;      memory[9945] <=  8'h00;      memory[9946] <=  8'h00;      memory[9947] <=  8'h00;      memory[9948] <=  8'h00;      memory[9949] <=  8'h00;      memory[9950] <=  8'h00;      memory[9951] <=  8'h00;      memory[9952] <=  8'h00;      memory[9953] <=  8'h00;      memory[9954] <=  8'h00;      memory[9955] <=  8'h00;      memory[9956] <=  8'h00;      memory[9957] <=  8'h00;      memory[9958] <=  8'h00;      memory[9959] <=  8'h00;      memory[9960] <=  8'h00;      memory[9961] <=  8'h00;      memory[9962] <=  8'h00;      memory[9963] <=  8'h00;      memory[9964] <=  8'h00;      memory[9965] <=  8'h00;      memory[9966] <=  8'h00;      memory[9967] <=  8'h00;      memory[9968] <=  8'h00;      memory[9969] <=  8'h00;      memory[9970] <=  8'h00;      memory[9971] <=  8'h00;      memory[9972] <=  8'h00;      memory[9973] <=  8'h00;      memory[9974] <=  8'h00;      memory[9975] <=  8'h00;      memory[9976] <=  8'h00;      memory[9977] <=  8'h00;      memory[9978] <=  8'h00;      memory[9979] <=  8'h00;      memory[9980] <=  8'h00;      memory[9981] <=  8'h00;      memory[9982] <=  8'h00;      memory[9983] <=  8'h00;      memory[9984] <=  8'h00;      memory[9985] <=  8'h00;      memory[9986] <=  8'h00;      memory[9987] <=  8'h00;      memory[9988] <=  8'h00;      memory[9989] <=  8'h00;      memory[9990] <=  8'h00;      memory[9991] <=  8'h00;      memory[9992] <=  8'h00;      memory[9993] <=  8'h00;      memory[9994] <=  8'h00;      memory[9995] <=  8'h00;      memory[9996] <=  8'h00;      memory[9997] <=  8'h00;      memory[9998] <=  8'h00;      memory[9999] <=  8'h00;      memory[10000] <=  8'h00;      memory[10001] <=  8'h00;      memory[10002] <=  8'h00;      memory[10003] <=  8'h00;      memory[10004] <=  8'h00;      memory[10005] <=  8'h00;      memory[10006] <=  8'h00;      memory[10007] <=  8'h00;      memory[10008] <=  8'h00;      memory[10009] <=  8'h00;      memory[10010] <=  8'h00;      memory[10011] <=  8'h00;      memory[10012] <=  8'h00;      memory[10013] <=  8'h00;      memory[10014] <=  8'h00;      memory[10015] <=  8'h00;      memory[10016] <=  8'h00;      memory[10017] <=  8'h00;      memory[10018] <=  8'h00;      memory[10019] <=  8'h00;      memory[10020] <=  8'h00;      memory[10021] <=  8'h00;      memory[10022] <=  8'h00;      memory[10023] <=  8'h00;      memory[10024] <=  8'h00;      memory[10025] <=  8'h00;      memory[10026] <=  8'h00;      memory[10027] <=  8'h00;      memory[10028] <=  8'h00;      memory[10029] <=  8'h00;      memory[10030] <=  8'h00;      memory[10031] <=  8'h00;      memory[10032] <=  8'h00;      memory[10033] <=  8'h00;      memory[10034] <=  8'h00;      memory[10035] <=  8'h00;      memory[10036] <=  8'h00;      memory[10037] <=  8'h00;      memory[10038] <=  8'h00;      memory[10039] <=  8'h00;      memory[10040] <=  8'h00;      memory[10041] <=  8'h00;      memory[10042] <=  8'h00;      memory[10043] <=  8'h00;      memory[10044] <=  8'h00;      memory[10045] <=  8'h00;      memory[10046] <=  8'h00;      memory[10047] <=  8'h00;      memory[10048] <=  8'h00;      memory[10049] <=  8'h00;      memory[10050] <=  8'h00;      memory[10051] <=  8'h00;      memory[10052] <=  8'h00;      memory[10053] <=  8'h00;      memory[10054] <=  8'h00;      memory[10055] <=  8'h00;      memory[10056] <=  8'h00;      memory[10057] <=  8'h00;      memory[10058] <=  8'h00;      memory[10059] <=  8'h00;      memory[10060] <=  8'h00;      memory[10061] <=  8'h00;      memory[10062] <=  8'h00;      memory[10063] <=  8'h00;      memory[10064] <=  8'h00;      memory[10065] <=  8'h00;      memory[10066] <=  8'h00;      memory[10067] <=  8'h00;      memory[10068] <=  8'h00;      memory[10069] <=  8'h00;      memory[10070] <=  8'h00;      memory[10071] <=  8'h00;      memory[10072] <=  8'h00;      memory[10073] <=  8'h00;      memory[10074] <=  8'h00;      memory[10075] <=  8'h00;      memory[10076] <=  8'h00;      memory[10077] <=  8'h00;      memory[10078] <=  8'h00;      memory[10079] <=  8'h00;      memory[10080] <=  8'h00;      memory[10081] <=  8'h00;      memory[10082] <=  8'h00;      memory[10083] <=  8'h00;      memory[10084] <=  8'h00;      memory[10085] <=  8'h00;      memory[10086] <=  8'h00;      memory[10087] <=  8'h00;      memory[10088] <=  8'h00;      memory[10089] <=  8'h00;      memory[10090] <=  8'h00;      memory[10091] <=  8'h00;      memory[10092] <=  8'h00;      memory[10093] <=  8'h00;      memory[10094] <=  8'h00;      memory[10095] <=  8'h00;      memory[10096] <=  8'h00;      memory[10097] <=  8'h00;      memory[10098] <=  8'h00;      memory[10099] <=  8'h00;      memory[10100] <=  8'h00;      memory[10101] <=  8'h00;      memory[10102] <=  8'h00;      memory[10103] <=  8'h00;      memory[10104] <=  8'h00;      memory[10105] <=  8'h00;      memory[10106] <=  8'h00;      memory[10107] <=  8'h00;      memory[10108] <=  8'h00;      memory[10109] <=  8'h00;      memory[10110] <=  8'h00;      memory[10111] <=  8'h00;      memory[10112] <=  8'h00;      memory[10113] <=  8'h00;      memory[10114] <=  8'h00;      memory[10115] <=  8'h00;      memory[10116] <=  8'h00;      memory[10117] <=  8'h00;      memory[10118] <=  8'h00;      memory[10119] <=  8'h00;      memory[10120] <=  8'h00;      memory[10121] <=  8'h00;      memory[10122] <=  8'h00;      memory[10123] <=  8'h00;      memory[10124] <=  8'h00;      memory[10125] <=  8'h00;      memory[10126] <=  8'h00;      memory[10127] <=  8'h00;      memory[10128] <=  8'h00;      memory[10129] <=  8'h00;      memory[10130] <=  8'h00;      memory[10131] <=  8'h00;      memory[10132] <=  8'h00;      memory[10133] <=  8'h00;      memory[10134] <=  8'h00;      memory[10135] <=  8'h00;      memory[10136] <=  8'h00;      memory[10137] <=  8'h00;      memory[10138] <=  8'h00;      memory[10139] <=  8'h00;      memory[10140] <=  8'h00;      memory[10141] <=  8'h00;      memory[10142] <=  8'h00;      memory[10143] <=  8'h00;      memory[10144] <=  8'h00;      memory[10145] <=  8'h00;      memory[10146] <=  8'h00;      memory[10147] <=  8'h00;      memory[10148] <=  8'h00;      memory[10149] <=  8'h00;      memory[10150] <=  8'h00;      memory[10151] <=  8'h00;      memory[10152] <=  8'h00;      memory[10153] <=  8'h00;      memory[10154] <=  8'h00;      memory[10155] <=  8'h00;      memory[10156] <=  8'h00;      memory[10157] <=  8'h00;      memory[10158] <=  8'h00;      memory[10159] <=  8'h00;      memory[10160] <=  8'h00;      memory[10161] <=  8'h00;      memory[10162] <=  8'h00;      memory[10163] <=  8'h00;      memory[10164] <=  8'h00;      memory[10165] <=  8'h00;      memory[10166] <=  8'h00;      memory[10167] <=  8'h00;      memory[10168] <=  8'h00;      memory[10169] <=  8'h00;      memory[10170] <=  8'h00;      memory[10171] <=  8'h00;      memory[10172] <=  8'h00;      memory[10173] <=  8'h00;      memory[10174] <=  8'h00;      memory[10175] <=  8'h00;      memory[10176] <=  8'h00;      memory[10177] <=  8'h00;      memory[10178] <=  8'h00;      memory[10179] <=  8'h00;      memory[10180] <=  8'h00;      memory[10181] <=  8'h00;      memory[10182] <=  8'h00;      memory[10183] <=  8'h00;      memory[10184] <=  8'h00;      memory[10185] <=  8'h00;      memory[10186] <=  8'h00;      memory[10187] <=  8'h00;      memory[10188] <=  8'h00;      memory[10189] <=  8'h00;      memory[10190] <=  8'h00;      memory[10191] <=  8'h00;      memory[10192] <=  8'h00;      memory[10193] <=  8'h00;      memory[10194] <=  8'h00;      memory[10195] <=  8'h00;      memory[10196] <=  8'h00;      memory[10197] <=  8'h00;      memory[10198] <=  8'h00;      memory[10199] <=  8'h00;      memory[10200] <=  8'h00;      memory[10201] <=  8'h00;      memory[10202] <=  8'h00;      memory[10203] <=  8'h00;      memory[10204] <=  8'h00;      memory[10205] <=  8'h00;      memory[10206] <=  8'h00;      memory[10207] <=  8'h00;      memory[10208] <=  8'h00;      memory[10209] <=  8'h00;      memory[10210] <=  8'h00;      memory[10211] <=  8'h00;      memory[10212] <=  8'h00;      memory[10213] <=  8'h00;      memory[10214] <=  8'h00;      memory[10215] <=  8'h00;      memory[10216] <=  8'h00;      memory[10217] <=  8'h00;      memory[10218] <=  8'h00;      memory[10219] <=  8'h00;      memory[10220] <=  8'h00;      memory[10221] <=  8'h00;      memory[10222] <=  8'h00;      memory[10223] <=  8'h00;      memory[10224] <=  8'h00;      memory[10225] <=  8'h00;      memory[10226] <=  8'h00;      memory[10227] <=  8'h00;      memory[10228] <=  8'h00;      memory[10229] <=  8'h00;      memory[10230] <=  8'h00;      memory[10231] <=  8'h00;      memory[10232] <=  8'h00;      memory[10233] <=  8'h00;      memory[10234] <=  8'h00;      memory[10235] <=  8'h00;      memory[10236] <=  8'h00;      memory[10237] <=  8'h00;      memory[10238] <=  8'h00;      memory[10239] <=  8'h00;      memory[10240] <=  8'h00;      memory[10241] <=  8'h00;      memory[10242] <=  8'h00;      memory[10243] <=  8'h00;      memory[10244] <=  8'h00;      memory[10245] <=  8'h00;      memory[10246] <=  8'h00;      memory[10247] <=  8'h00;      memory[10248] <=  8'h00;      memory[10249] <=  8'h00;      memory[10250] <=  8'h00;      memory[10251] <=  8'h00;      memory[10252] <=  8'h00;      memory[10253] <=  8'h00;      memory[10254] <=  8'h00;      memory[10255] <=  8'h00;      memory[10256] <=  8'h00;      memory[10257] <=  8'h00;      memory[10258] <=  8'h00;      memory[10259] <=  8'h00;      memory[10260] <=  8'h00;      memory[10261] <=  8'h00;      memory[10262] <=  8'h00;      memory[10263] <=  8'h00;      memory[10264] <=  8'h00;      memory[10265] <=  8'h00;      memory[10266] <=  8'h00;      memory[10267] <=  8'h00;      memory[10268] <=  8'h00;      memory[10269] <=  8'h00;      memory[10270] <=  8'h00;      memory[10271] <=  8'h00;      memory[10272] <=  8'h00;      memory[10273] <=  8'h00;      memory[10274] <=  8'h00;      memory[10275] <=  8'h00;      memory[10276] <=  8'h00;      memory[10277] <=  8'h00;      memory[10278] <=  8'h00;      memory[10279] <=  8'h00;      memory[10280] <=  8'h00;      memory[10281] <=  8'h00;      memory[10282] <=  8'h00;      memory[10283] <=  8'h00;      memory[10284] <=  8'h00;      memory[10285] <=  8'h00;      memory[10286] <=  8'h00;      memory[10287] <=  8'h00;      memory[10288] <=  8'h00;      memory[10289] <=  8'h00;      memory[10290] <=  8'h00;      memory[10291] <=  8'h00;      memory[10292] <=  8'h00;      memory[10293] <=  8'h00;      memory[10294] <=  8'h00;      memory[10295] <=  8'h00;      memory[10296] <=  8'h00;      memory[10297] <=  8'h00;      memory[10298] <=  8'h00;      memory[10299] <=  8'h00;      memory[10300] <=  8'h00;      memory[10301] <=  8'h00;      memory[10302] <=  8'h00;      memory[10303] <=  8'h00;      memory[10304] <=  8'h00;      memory[10305] <=  8'h00;      memory[10306] <=  8'h00;      memory[10307] <=  8'h00;      memory[10308] <=  8'h00;      memory[10309] <=  8'h00;      memory[10310] <=  8'h00;      memory[10311] <=  8'h00;      memory[10312] <=  8'h00;      memory[10313] <=  8'h00;      memory[10314] <=  8'h00;      memory[10315] <=  8'h00;      memory[10316] <=  8'h00;      memory[10317] <=  8'h00;      memory[10318] <=  8'h00;      memory[10319] <=  8'h00;      memory[10320] <=  8'h00;      memory[10321] <=  8'h00;      memory[10322] <=  8'h00;      memory[10323] <=  8'h00;      memory[10324] <=  8'h00;      memory[10325] <=  8'h00;      memory[10326] <=  8'h00;      memory[10327] <=  8'h00;      memory[10328] <=  8'h00;      memory[10329] <=  8'h00;      memory[10330] <=  8'h00;      memory[10331] <=  8'h00;      memory[10332] <=  8'h00;      memory[10333] <=  8'h00;      memory[10334] <=  8'h00;      memory[10335] <=  8'h00;      memory[10336] <=  8'h00;      memory[10337] <=  8'h00;      memory[10338] <=  8'h00;      memory[10339] <=  8'h00;      memory[10340] <=  8'h00;      memory[10341] <=  8'h00;      memory[10342] <=  8'h00;      memory[10343] <=  8'h00;      memory[10344] <=  8'h00;      memory[10345] <=  8'h00;      memory[10346] <=  8'h00;      memory[10347] <=  8'h00;      memory[10348] <=  8'h00;      memory[10349] <=  8'h00;      memory[10350] <=  8'h00;      memory[10351] <=  8'h00;      memory[10352] <=  8'h00;      memory[10353] <=  8'h00;      memory[10354] <=  8'h00;      memory[10355] <=  8'h00;      memory[10356] <=  8'h00;      memory[10357] <=  8'h00;      memory[10358] <=  8'h00;      memory[10359] <=  8'h00;      memory[10360] <=  8'h00;      memory[10361] <=  8'h00;      memory[10362] <=  8'h00;      memory[10363] <=  8'h00;      memory[10364] <=  8'h00;      memory[10365] <=  8'h00;      memory[10366] <=  8'h00;      memory[10367] <=  8'h00;      memory[10368] <=  8'h00;      memory[10369] <=  8'h00;      memory[10370] <=  8'h00;      memory[10371] <=  8'h00;      memory[10372] <=  8'h00;      memory[10373] <=  8'h00;      memory[10374] <=  8'h00;      memory[10375] <=  8'h00;      memory[10376] <=  8'h00;      memory[10377] <=  8'h00;      memory[10378] <=  8'h00;      memory[10379] <=  8'h00;      memory[10380] <=  8'h00;      memory[10381] <=  8'h00;      memory[10382] <=  8'h00;      memory[10383] <=  8'h00;      memory[10384] <=  8'h00;      memory[10385] <=  8'h00;      memory[10386] <=  8'h00;      memory[10387] <=  8'h00;      memory[10388] <=  8'h00;      memory[10389] <=  8'h00;      memory[10390] <=  8'h00;      memory[10391] <=  8'h00;      memory[10392] <=  8'h00;      memory[10393] <=  8'h00;      memory[10394] <=  8'h00;      memory[10395] <=  8'h00;      memory[10396] <=  8'h00;      memory[10397] <=  8'h00;      memory[10398] <=  8'h00;      memory[10399] <=  8'h00;      memory[10400] <=  8'h00;      memory[10401] <=  8'h00;      memory[10402] <=  8'h00;      memory[10403] <=  8'h00;      memory[10404] <=  8'h00;      memory[10405] <=  8'h00;      memory[10406] <=  8'h00;      memory[10407] <=  8'h00;      memory[10408] <=  8'h00;      memory[10409] <=  8'h00;      memory[10410] <=  8'h00;      memory[10411] <=  8'h00;      memory[10412] <=  8'h00;      memory[10413] <=  8'h00;      memory[10414] <=  8'h00;      memory[10415] <=  8'h00;      memory[10416] <=  8'h00;      memory[10417] <=  8'h00;      memory[10418] <=  8'h00;      memory[10419] <=  8'h00;      memory[10420] <=  8'h00;      memory[10421] <=  8'h00;      memory[10422] <=  8'h00;      memory[10423] <=  8'h00;      memory[10424] <=  8'h00;      memory[10425] <=  8'h00;      memory[10426] <=  8'h00;      memory[10427] <=  8'h00;      memory[10428] <=  8'h00;      memory[10429] <=  8'h00;      memory[10430] <=  8'h00;      memory[10431] <=  8'h00;      memory[10432] <=  8'h00;      memory[10433] <=  8'h00;      memory[10434] <=  8'h00;      memory[10435] <=  8'h00;      memory[10436] <=  8'h00;      memory[10437] <=  8'h00;      memory[10438] <=  8'h00;      memory[10439] <=  8'h00;      memory[10440] <=  8'h00;      memory[10441] <=  8'h00;      memory[10442] <=  8'h00;      memory[10443] <=  8'h00;      memory[10444] <=  8'h00;      memory[10445] <=  8'h00;      memory[10446] <=  8'h00;      memory[10447] <=  8'h00;      memory[10448] <=  8'h00;      memory[10449] <=  8'h00;      memory[10450] <=  8'h00;      memory[10451] <=  8'h00;      memory[10452] <=  8'h00;      memory[10453] <=  8'h00;      memory[10454] <=  8'h00;      memory[10455] <=  8'h00;      memory[10456] <=  8'h00;      memory[10457] <=  8'h00;      memory[10458] <=  8'h00;      memory[10459] <=  8'h00;      memory[10460] <=  8'h00;      memory[10461] <=  8'h00;      memory[10462] <=  8'h00;      memory[10463] <=  8'h00;      memory[10464] <=  8'h00;      memory[10465] <=  8'h00;      memory[10466] <=  8'h00;      memory[10467] <=  8'h00;      memory[10468] <=  8'h00;      memory[10469] <=  8'h00;      memory[10470] <=  8'h00;      memory[10471] <=  8'h00;      memory[10472] <=  8'h00;      memory[10473] <=  8'h00;      memory[10474] <=  8'h00;      memory[10475] <=  8'h00;      memory[10476] <=  8'h00;      memory[10477] <=  8'h00;      memory[10478] <=  8'h00;      memory[10479] <=  8'h00;      memory[10480] <=  8'h00;      memory[10481] <=  8'h00;      memory[10482] <=  8'h00;      memory[10483] <=  8'h00;      memory[10484] <=  8'h00;      memory[10485] <=  8'h00;      memory[10486] <=  8'h00;      memory[10487] <=  8'h00;      memory[10488] <=  8'h00;      memory[10489] <=  8'h00;      memory[10490] <=  8'h00;      memory[10491] <=  8'h00;      memory[10492] <=  8'h00;      memory[10493] <=  8'h00;      memory[10494] <=  8'h00;      memory[10495] <=  8'h00;      memory[10496] <=  8'h00;      memory[10497] <=  8'h00;      memory[10498] <=  8'h00;      memory[10499] <=  8'h00;      memory[10500] <=  8'h00;      memory[10501] <=  8'h00;      memory[10502] <=  8'h00;      memory[10503] <=  8'h00;      memory[10504] <=  8'h00;      memory[10505] <=  8'h00;      memory[10506] <=  8'h00;      memory[10507] <=  8'h00;      memory[10508] <=  8'h00;      memory[10509] <=  8'h00;      memory[10510] <=  8'h00;      memory[10511] <=  8'h00;      memory[10512] <=  8'h00;      memory[10513] <=  8'h00;      memory[10514] <=  8'h00;      memory[10515] <=  8'h00;      memory[10516] <=  8'h00;      memory[10517] <=  8'h00;      memory[10518] <=  8'h00;      memory[10519] <=  8'h00;      memory[10520] <=  8'h00;      memory[10521] <=  8'h00;      memory[10522] <=  8'h00;      memory[10523] <=  8'h00;      memory[10524] <=  8'h00;      memory[10525] <=  8'h00;      memory[10526] <=  8'h00;      memory[10527] <=  8'h00;      memory[10528] <=  8'h00;      memory[10529] <=  8'h00;      memory[10530] <=  8'h00;      memory[10531] <=  8'h00;      memory[10532] <=  8'h00;      memory[10533] <=  8'h00;      memory[10534] <=  8'h00;      memory[10535] <=  8'h00;      memory[10536] <=  8'h00;      memory[10537] <=  8'h00;      memory[10538] <=  8'h00;      memory[10539] <=  8'h00;      memory[10540] <=  8'h00;      memory[10541] <=  8'h00;      memory[10542] <=  8'h00;      memory[10543] <=  8'h00;      memory[10544] <=  8'h00;      memory[10545] <=  8'h00;      memory[10546] <=  8'h00;      memory[10547] <=  8'h00;      memory[10548] <=  8'h00;      memory[10549] <=  8'h00;      memory[10550] <=  8'h00;      memory[10551] <=  8'h00;      memory[10552] <=  8'h00;      memory[10553] <=  8'h00;      memory[10554] <=  8'h00;      memory[10555] <=  8'h00;      memory[10556] <=  8'h00;      memory[10557] <=  8'h00;      memory[10558] <=  8'h00;      memory[10559] <=  8'h00;      memory[10560] <=  8'h00;      memory[10561] <=  8'h00;      memory[10562] <=  8'h00;      memory[10563] <=  8'h00;      memory[10564] <=  8'h00;      memory[10565] <=  8'h00;      memory[10566] <=  8'h00;      memory[10567] <=  8'h00;      memory[10568] <=  8'h00;      memory[10569] <=  8'h00;      memory[10570] <=  8'h00;      memory[10571] <=  8'h00;      memory[10572] <=  8'h00;      memory[10573] <=  8'h00;      memory[10574] <=  8'h00;      memory[10575] <=  8'h00;      memory[10576] <=  8'h00;      memory[10577] <=  8'h00;      memory[10578] <=  8'h00;      memory[10579] <=  8'h00;      memory[10580] <=  8'h00;      memory[10581] <=  8'h00;      memory[10582] <=  8'h00;      memory[10583] <=  8'h00;      memory[10584] <=  8'h00;      memory[10585] <=  8'h00;      memory[10586] <=  8'h00;      memory[10587] <=  8'h00;      memory[10588] <=  8'h00;      memory[10589] <=  8'h00;      memory[10590] <=  8'h00;      memory[10591] <=  8'h00;      memory[10592] <=  8'h00;      memory[10593] <=  8'h00;      memory[10594] <=  8'h00;      memory[10595] <=  8'h00;      memory[10596] <=  8'h00;      memory[10597] <=  8'h00;      memory[10598] <=  8'h00;      memory[10599] <=  8'h00;      memory[10600] <=  8'h00;      memory[10601] <=  8'h00;      memory[10602] <=  8'h00;      memory[10603] <=  8'h00;      memory[10604] <=  8'h00;      memory[10605] <=  8'h00;      memory[10606] <=  8'h00;      memory[10607] <=  8'h00;      memory[10608] <=  8'h00;      memory[10609] <=  8'h00;      memory[10610] <=  8'h00;      memory[10611] <=  8'h00;      memory[10612] <=  8'h00;      memory[10613] <=  8'h00;      memory[10614] <=  8'h00;      memory[10615] <=  8'h00;      memory[10616] <=  8'h00;      memory[10617] <=  8'h00;      memory[10618] <=  8'h00;      memory[10619] <=  8'h00;      memory[10620] <=  8'h00;      memory[10621] <=  8'h00;      memory[10622] <=  8'h00;      memory[10623] <=  8'h00;      memory[10624] <=  8'h00;      memory[10625] <=  8'h00;      memory[10626] <=  8'h00;      memory[10627] <=  8'h00;      memory[10628] <=  8'h00;      memory[10629] <=  8'h00;      memory[10630] <=  8'h00;      memory[10631] <=  8'h00;      memory[10632] <=  8'h00;      memory[10633] <=  8'h00;      memory[10634] <=  8'h00;      memory[10635] <=  8'h00;      memory[10636] <=  8'h00;      memory[10637] <=  8'h00;      memory[10638] <=  8'h00;      memory[10639] <=  8'h00;      memory[10640] <=  8'h00;      memory[10641] <=  8'h00;      memory[10642] <=  8'h00;      memory[10643] <=  8'h00;      memory[10644] <=  8'h00;      memory[10645] <=  8'h00;      memory[10646] <=  8'h00;      memory[10647] <=  8'h00;      memory[10648] <=  8'h00;      memory[10649] <=  8'h00;      memory[10650] <=  8'h00;      memory[10651] <=  8'h00;      memory[10652] <=  8'h00;      memory[10653] <=  8'h00;      memory[10654] <=  8'h00;      memory[10655] <=  8'h00;      memory[10656] <=  8'h00;      memory[10657] <=  8'h00;      memory[10658] <=  8'h00;      memory[10659] <=  8'h00;      memory[10660] <=  8'h00;      memory[10661] <=  8'h00;      memory[10662] <=  8'h00;      memory[10663] <=  8'h00;      memory[10664] <=  8'h00;      memory[10665] <=  8'h00;      memory[10666] <=  8'h00;      memory[10667] <=  8'h00;      memory[10668] <=  8'h00;      memory[10669] <=  8'h00;      memory[10670] <=  8'h00;      memory[10671] <=  8'h00;      memory[10672] <=  8'h00;      memory[10673] <=  8'h00;      memory[10674] <=  8'h00;      memory[10675] <=  8'h00;      memory[10676] <=  8'h00;      memory[10677] <=  8'h00;      memory[10678] <=  8'h00;      memory[10679] <=  8'h00;      memory[10680] <=  8'h00;      memory[10681] <=  8'h00;      memory[10682] <=  8'h00;      memory[10683] <=  8'h00;      memory[10684] <=  8'h00;      memory[10685] <=  8'h00;      memory[10686] <=  8'h00;      memory[10687] <=  8'h00;      memory[10688] <=  8'h00;      memory[10689] <=  8'h00;      memory[10690] <=  8'h00;      memory[10691] <=  8'h00;      memory[10692] <=  8'h00;      memory[10693] <=  8'h00;      memory[10694] <=  8'h00;      memory[10695] <=  8'h00;      memory[10696] <=  8'h00;      memory[10697] <=  8'h00;      memory[10698] <=  8'h00;      memory[10699] <=  8'h00;      memory[10700] <=  8'h00;      memory[10701] <=  8'h00;      memory[10702] <=  8'h00;      memory[10703] <=  8'h00;      memory[10704] <=  8'h00;      memory[10705] <=  8'h00;      memory[10706] <=  8'h00;      memory[10707] <=  8'h00;      memory[10708] <=  8'h00;      memory[10709] <=  8'h00;      memory[10710] <=  8'h00;      memory[10711] <=  8'h00;      memory[10712] <=  8'h00;      memory[10713] <=  8'h00;      memory[10714] <=  8'h00;      memory[10715] <=  8'h00;      memory[10716] <=  8'h00;      memory[10717] <=  8'h00;      memory[10718] <=  8'h00;      memory[10719] <=  8'h00;      memory[10720] <=  8'h00;      memory[10721] <=  8'h00;      memory[10722] <=  8'h00;      memory[10723] <=  8'h00;      memory[10724] <=  8'h00;      memory[10725] <=  8'h00;      memory[10726] <=  8'h00;      memory[10727] <=  8'h00;      memory[10728] <=  8'h00;      memory[10729] <=  8'h00;      memory[10730] <=  8'h00;      memory[10731] <=  8'h00;      memory[10732] <=  8'h00;      memory[10733] <=  8'h00;      memory[10734] <=  8'h00;      memory[10735] <=  8'h00;      memory[10736] <=  8'h00;      memory[10737] <=  8'h00;      memory[10738] <=  8'h00;      memory[10739] <=  8'h00;      memory[10740] <=  8'h00;      memory[10741] <=  8'h00;      memory[10742] <=  8'h00;      memory[10743] <=  8'h00;      memory[10744] <=  8'h00;      memory[10745] <=  8'h00;      memory[10746] <=  8'h00;      memory[10747] <=  8'h00;      memory[10748] <=  8'h00;      memory[10749] <=  8'h00;      memory[10750] <=  8'h00;      memory[10751] <=  8'h00;      memory[10752] <=  8'h00;      memory[10753] <=  8'h00;      memory[10754] <=  8'h00;      memory[10755] <=  8'h00;      memory[10756] <=  8'h00;      memory[10757] <=  8'h00;      memory[10758] <=  8'h00;      memory[10759] <=  8'h00;      memory[10760] <=  8'h00;      memory[10761] <=  8'h00;      memory[10762] <=  8'h00;      memory[10763] <=  8'h00;      memory[10764] <=  8'h00;      memory[10765] <=  8'h00;      memory[10766] <=  8'h00;      memory[10767] <=  8'h00;      memory[10768] <=  8'h00;      memory[10769] <=  8'h00;      memory[10770] <=  8'h00;      memory[10771] <=  8'h00;      memory[10772] <=  8'h00;      memory[10773] <=  8'h00;      memory[10774] <=  8'h00;      memory[10775] <=  8'h00;      memory[10776] <=  8'h00;      memory[10777] <=  8'h00;      memory[10778] <=  8'h00;      memory[10779] <=  8'h00;      memory[10780] <=  8'h00;      memory[10781] <=  8'h00;      memory[10782] <=  8'h00;      memory[10783] <=  8'h00;      memory[10784] <=  8'h00;      memory[10785] <=  8'h00;      memory[10786] <=  8'h00;      memory[10787] <=  8'h00;      memory[10788] <=  8'h00;      memory[10789] <=  8'h00;      memory[10790] <=  8'h00;      memory[10791] <=  8'h00;      memory[10792] <=  8'h00;      memory[10793] <=  8'h00;      memory[10794] <=  8'h00;      memory[10795] <=  8'h00;      memory[10796] <=  8'h00;      memory[10797] <=  8'h00;      memory[10798] <=  8'h00;      memory[10799] <=  8'h00;      memory[10800] <=  8'h00;      memory[10801] <=  8'h00;      memory[10802] <=  8'h00;      memory[10803] <=  8'h00;      memory[10804] <=  8'h00;      memory[10805] <=  8'h00;      memory[10806] <=  8'h00;      memory[10807] <=  8'h00;      memory[10808] <=  8'h00;      memory[10809] <=  8'h00;      memory[10810] <=  8'h00;      memory[10811] <=  8'h00;      memory[10812] <=  8'h00;      memory[10813] <=  8'h00;      memory[10814] <=  8'h00;      memory[10815] <=  8'h00;      memory[10816] <=  8'h00;      memory[10817] <=  8'h00;      memory[10818] <=  8'h00;      memory[10819] <=  8'h00;      memory[10820] <=  8'h00;      memory[10821] <=  8'h00;      memory[10822] <=  8'h00;      memory[10823] <=  8'h00;      memory[10824] <=  8'h00;      memory[10825] <=  8'h00;      memory[10826] <=  8'h00;      memory[10827] <=  8'h00;      memory[10828] <=  8'h00;      memory[10829] <=  8'h00;      memory[10830] <=  8'h00;      memory[10831] <=  8'h00;      memory[10832] <=  8'h00;      memory[10833] <=  8'h00;      memory[10834] <=  8'h00;      memory[10835] <=  8'h00;      memory[10836] <=  8'h00;      memory[10837] <=  8'h00;      memory[10838] <=  8'h00;      memory[10839] <=  8'h00;      memory[10840] <=  8'h00;      memory[10841] <=  8'h00;      memory[10842] <=  8'h00;      memory[10843] <=  8'h00;      memory[10844] <=  8'h00;      memory[10845] <=  8'h00;      memory[10846] <=  8'h00;      memory[10847] <=  8'h00;      memory[10848] <=  8'h00;      memory[10849] <=  8'h00;      memory[10850] <=  8'h00;      memory[10851] <=  8'h00;      memory[10852] <=  8'h00;      memory[10853] <=  8'h00;      memory[10854] <=  8'h00;      memory[10855] <=  8'h00;      memory[10856] <=  8'h00;      memory[10857] <=  8'h00;      memory[10858] <=  8'h00;      memory[10859] <=  8'h00;      memory[10860] <=  8'h00;      memory[10861] <=  8'h00;      memory[10862] <=  8'h00;      memory[10863] <=  8'h00;      memory[10864] <=  8'h00;      memory[10865] <=  8'h00;      memory[10866] <=  8'h00;      memory[10867] <=  8'h00;      memory[10868] <=  8'h00;      memory[10869] <=  8'h00;      memory[10870] <=  8'h00;      memory[10871] <=  8'h00;      memory[10872] <=  8'h00;      memory[10873] <=  8'h00;      memory[10874] <=  8'h00;      memory[10875] <=  8'h00;      memory[10876] <=  8'h00;      memory[10877] <=  8'h00;      memory[10878] <=  8'h00;      memory[10879] <=  8'h00;      memory[10880] <=  8'h00;      memory[10881] <=  8'h00;      memory[10882] <=  8'h00;      memory[10883] <=  8'h00;      memory[10884] <=  8'h00;      memory[10885] <=  8'h00;      memory[10886] <=  8'h00;      memory[10887] <=  8'h00;      memory[10888] <=  8'h00;      memory[10889] <=  8'h00;      memory[10890] <=  8'h00;      memory[10891] <=  8'h00;      memory[10892] <=  8'h00;      memory[10893] <=  8'h00;      memory[10894] <=  8'h00;      memory[10895] <=  8'h00;      memory[10896] <=  8'h00;      memory[10897] <=  8'h00;      memory[10898] <=  8'h00;      memory[10899] <=  8'h00;      memory[10900] <=  8'h00;      memory[10901] <=  8'h00;      memory[10902] <=  8'h00;      memory[10903] <=  8'h00;      memory[10904] <=  8'h00;      memory[10905] <=  8'h00;      memory[10906] <=  8'h00;      memory[10907] <=  8'h00;      memory[10908] <=  8'h00;      memory[10909] <=  8'h00;      memory[10910] <=  8'h00;      memory[10911] <=  8'h00;      memory[10912] <=  8'h00;      memory[10913] <=  8'h00;      memory[10914] <=  8'h00;      memory[10915] <=  8'h00;      memory[10916] <=  8'h00;      memory[10917] <=  8'h00;      memory[10918] <=  8'h00;      memory[10919] <=  8'h00;      memory[10920] <=  8'h00;      memory[10921] <=  8'h00;      memory[10922] <=  8'h00;      memory[10923] <=  8'h00;      memory[10924] <=  8'h00;      memory[10925] <=  8'h00;      memory[10926] <=  8'h00;      memory[10927] <=  8'h00;      memory[10928] <=  8'h00;      memory[10929] <=  8'h00;      memory[10930] <=  8'h00;      memory[10931] <=  8'h00;      memory[10932] <=  8'h00;      memory[10933] <=  8'h00;      memory[10934] <=  8'h00;      memory[10935] <=  8'h00;      memory[10936] <=  8'h00;      memory[10937] <=  8'h00;      memory[10938] <=  8'h00;      memory[10939] <=  8'h00;      memory[10940] <=  8'h00;      memory[10941] <=  8'h00;      memory[10942] <=  8'h00;      memory[10943] <=  8'h00;      memory[10944] <=  8'h00;      memory[10945] <=  8'h00;      memory[10946] <=  8'h00;      memory[10947] <=  8'h00;      memory[10948] <=  8'h00;      memory[10949] <=  8'h00;      memory[10950] <=  8'h00;      memory[10951] <=  8'h00;      memory[10952] <=  8'h00;      memory[10953] <=  8'h00;      memory[10954] <=  8'h00;      memory[10955] <=  8'h00;      memory[10956] <=  8'h00;      memory[10957] <=  8'h00;      memory[10958] <=  8'h00;      memory[10959] <=  8'h00;      memory[10960] <=  8'h00;      memory[10961] <=  8'h00;      memory[10962] <=  8'h00;      memory[10963] <=  8'h00;      memory[10964] <=  8'h00;      memory[10965] <=  8'h00;      memory[10966] <=  8'h00;      memory[10967] <=  8'h00;      memory[10968] <=  8'h00;      memory[10969] <=  8'h00;      memory[10970] <=  8'h00;      memory[10971] <=  8'h00;      memory[10972] <=  8'h00;      memory[10973] <=  8'h00;      memory[10974] <=  8'h00;      memory[10975] <=  8'h00;      memory[10976] <=  8'h00;      memory[10977] <=  8'h00;      memory[10978] <=  8'h00;      memory[10979] <=  8'h00;      memory[10980] <=  8'h00;      memory[10981] <=  8'h00;      memory[10982] <=  8'h00;      memory[10983] <=  8'h00;      memory[10984] <=  8'h00;      memory[10985] <=  8'h00;      memory[10986] <=  8'h00;      memory[10987] <=  8'h00;      memory[10988] <=  8'h00;      memory[10989] <=  8'h00;      memory[10990] <=  8'h00;      memory[10991] <=  8'h00;      memory[10992] <=  8'h00;      memory[10993] <=  8'h00;      memory[10994] <=  8'h00;      memory[10995] <=  8'h00;      memory[10996] <=  8'h00;      memory[10997] <=  8'h00;      memory[10998] <=  8'h00;      memory[10999] <=  8'h00;      memory[11000] <=  8'h00;      memory[11001] <=  8'h00;      memory[11002] <=  8'h00;      memory[11003] <=  8'h00;      memory[11004] <=  8'h00;      memory[11005] <=  8'h00;      memory[11006] <=  8'h00;      memory[11007] <=  8'h00;      memory[11008] <=  8'h00;      memory[11009] <=  8'h00;      memory[11010] <=  8'h00;      memory[11011] <=  8'h00;      memory[11012] <=  8'h00;      memory[11013] <=  8'h00;      memory[11014] <=  8'h00;      memory[11015] <=  8'h00;      memory[11016] <=  8'h00;      memory[11017] <=  8'h00;      memory[11018] <=  8'h00;      memory[11019] <=  8'h00;      memory[11020] <=  8'h00;      memory[11021] <=  8'h00;      memory[11022] <=  8'h00;      memory[11023] <=  8'h00;      memory[11024] <=  8'h00;      memory[11025] <=  8'h00;      memory[11026] <=  8'h00;      memory[11027] <=  8'h00;      memory[11028] <=  8'h00;      memory[11029] <=  8'h00;      memory[11030] <=  8'h00;      memory[11031] <=  8'h00;      memory[11032] <=  8'h00;      memory[11033] <=  8'h00;      memory[11034] <=  8'h00;      memory[11035] <=  8'h00;      memory[11036] <=  8'h00;      memory[11037] <=  8'h00;      memory[11038] <=  8'h00;      memory[11039] <=  8'h00;      memory[11040] <=  8'h00;      memory[11041] <=  8'h00;      memory[11042] <=  8'h00;      memory[11043] <=  8'h00;      memory[11044] <=  8'h00;      memory[11045] <=  8'h00;      memory[11046] <=  8'h00;      memory[11047] <=  8'h00;      memory[11048] <=  8'h00;      memory[11049] <=  8'h00;      memory[11050] <=  8'h00;      memory[11051] <=  8'h00;      memory[11052] <=  8'h00;      memory[11053] <=  8'h00;      memory[11054] <=  8'h00;      memory[11055] <=  8'h00;      memory[11056] <=  8'h00;      memory[11057] <=  8'h00;      memory[11058] <=  8'h00;      memory[11059] <=  8'h00;      memory[11060] <=  8'h00;      memory[11061] <=  8'h00;      memory[11062] <=  8'h00;      memory[11063] <=  8'h00;      memory[11064] <=  8'h00;      memory[11065] <=  8'h00;      memory[11066] <=  8'h00;      memory[11067] <=  8'h00;      memory[11068] <=  8'h00;      memory[11069] <=  8'h00;      memory[11070] <=  8'h00;      memory[11071] <=  8'h00;      memory[11072] <=  8'h00;      memory[11073] <=  8'h00;      memory[11074] <=  8'h00;      memory[11075] <=  8'h00;      memory[11076] <=  8'h00;      memory[11077] <=  8'h00;      memory[11078] <=  8'h00;      memory[11079] <=  8'h00;      memory[11080] <=  8'h00;      memory[11081] <=  8'h00;      memory[11082] <=  8'h00;      memory[11083] <=  8'h00;      memory[11084] <=  8'h00;      memory[11085] <=  8'h00;      memory[11086] <=  8'h00;      memory[11087] <=  8'h00;      memory[11088] <=  8'h00;      memory[11089] <=  8'h00;      memory[11090] <=  8'h00;      memory[11091] <=  8'h00;      memory[11092] <=  8'h00;      memory[11093] <=  8'h00;      memory[11094] <=  8'h00;      memory[11095] <=  8'h00;      memory[11096] <=  8'h00;      memory[11097] <=  8'h00;      memory[11098] <=  8'h00;      memory[11099] <=  8'h00;      memory[11100] <=  8'h00;      memory[11101] <=  8'h00;      memory[11102] <=  8'h00;      memory[11103] <=  8'h00;      memory[11104] <=  8'h00;      memory[11105] <=  8'h00;      memory[11106] <=  8'h00;      memory[11107] <=  8'h00;      memory[11108] <=  8'h00;      memory[11109] <=  8'h00;      memory[11110] <=  8'h00;      memory[11111] <=  8'h00;      memory[11112] <=  8'h00;      memory[11113] <=  8'h00;      memory[11114] <=  8'h00;      memory[11115] <=  8'h00;      memory[11116] <=  8'h00;      memory[11117] <=  8'h00;      memory[11118] <=  8'h00;      memory[11119] <=  8'h00;      memory[11120] <=  8'h00;      memory[11121] <=  8'h00;      memory[11122] <=  8'h00;      memory[11123] <=  8'h00;      memory[11124] <=  8'h00;      memory[11125] <=  8'h00;      memory[11126] <=  8'h00;      memory[11127] <=  8'h00;      memory[11128] <=  8'h00;      memory[11129] <=  8'h00;      memory[11130] <=  8'h00;      memory[11131] <=  8'h00;      memory[11132] <=  8'h00;      memory[11133] <=  8'h00;      memory[11134] <=  8'h00;      memory[11135] <=  8'h00;      memory[11136] <=  8'h00;      memory[11137] <=  8'h00;      memory[11138] <=  8'h00;      memory[11139] <=  8'h00;      memory[11140] <=  8'h00;      memory[11141] <=  8'h00;      memory[11142] <=  8'h00;      memory[11143] <=  8'h00;      memory[11144] <=  8'h00;      memory[11145] <=  8'h00;      memory[11146] <=  8'h00;      memory[11147] <=  8'h00;      memory[11148] <=  8'h00;      memory[11149] <=  8'h00;      memory[11150] <=  8'h00;      memory[11151] <=  8'h00;      memory[11152] <=  8'h00;      memory[11153] <=  8'h00;      memory[11154] <=  8'h00;      memory[11155] <=  8'h00;      memory[11156] <=  8'h00;      memory[11157] <=  8'h00;      memory[11158] <=  8'h00;      memory[11159] <=  8'h00;      memory[11160] <=  8'h00;      memory[11161] <=  8'h00;      memory[11162] <=  8'h00;      memory[11163] <=  8'h00;      memory[11164] <=  8'h00;      memory[11165] <=  8'h00;      memory[11166] <=  8'h00;      memory[11167] <=  8'h00;      memory[11168] <=  8'h00;      memory[11169] <=  8'h00;      memory[11170] <=  8'h00;      memory[11171] <=  8'h00;      memory[11172] <=  8'h00;      memory[11173] <=  8'h00;      memory[11174] <=  8'h00;      memory[11175] <=  8'h00;      memory[11176] <=  8'h00;      memory[11177] <=  8'h00;      memory[11178] <=  8'h00;      memory[11179] <=  8'h00;      memory[11180] <=  8'h00;      memory[11181] <=  8'h00;      memory[11182] <=  8'h00;      memory[11183] <=  8'h00;      memory[11184] <=  8'h00;      memory[11185] <=  8'h00;      memory[11186] <=  8'h00;      memory[11187] <=  8'h00;      memory[11188] <=  8'h00;      memory[11189] <=  8'h00;      memory[11190] <=  8'h00;      memory[11191] <=  8'h00;      memory[11192] <=  8'h00;      memory[11193] <=  8'h00;      memory[11194] <=  8'h00;      memory[11195] <=  8'h00;      memory[11196] <=  8'h00;      memory[11197] <=  8'h00;      memory[11198] <=  8'h00;      memory[11199] <=  8'h00;      memory[11200] <=  8'h00;      memory[11201] <=  8'h00;      memory[11202] <=  8'h00;      memory[11203] <=  8'h00;      memory[11204] <=  8'h00;      memory[11205] <=  8'h00;      memory[11206] <=  8'h00;      memory[11207] <=  8'h00;      memory[11208] <=  8'h00;      memory[11209] <=  8'h00;      memory[11210] <=  8'h00;      memory[11211] <=  8'h00;      memory[11212] <=  8'h00;      memory[11213] <=  8'h00;      memory[11214] <=  8'h00;      memory[11215] <=  8'h00;      memory[11216] <=  8'h00;      memory[11217] <=  8'h00;      memory[11218] <=  8'h00;      memory[11219] <=  8'h00;      memory[11220] <=  8'h00;      memory[11221] <=  8'h00;      memory[11222] <=  8'h00;      memory[11223] <=  8'h00;      memory[11224] <=  8'h00;      memory[11225] <=  8'h00;      memory[11226] <=  8'h00;      memory[11227] <=  8'h00;      memory[11228] <=  8'h00;      memory[11229] <=  8'h00;      memory[11230] <=  8'h00;      memory[11231] <=  8'h00;      memory[11232] <=  8'h00;      memory[11233] <=  8'h00;      memory[11234] <=  8'h00;      memory[11235] <=  8'h00;      memory[11236] <=  8'h00;      memory[11237] <=  8'h00;      memory[11238] <=  8'h00;      memory[11239] <=  8'h00;      memory[11240] <=  8'h00;      memory[11241] <=  8'h00;      memory[11242] <=  8'h00;      memory[11243] <=  8'h00;      memory[11244] <=  8'h00;      memory[11245] <=  8'h00;      memory[11246] <=  8'h00;      memory[11247] <=  8'h00;      memory[11248] <=  8'h00;      memory[11249] <=  8'h00;      memory[11250] <=  8'h00;      memory[11251] <=  8'h00;      memory[11252] <=  8'h00;      memory[11253] <=  8'h00;      memory[11254] <=  8'h00;      memory[11255] <=  8'h00;      memory[11256] <=  8'h00;      memory[11257] <=  8'h00;      memory[11258] <=  8'h00;      memory[11259] <=  8'h00;      memory[11260] <=  8'h00;      memory[11261] <=  8'h00;      memory[11262] <=  8'h00;      memory[11263] <=  8'h00;      memory[11264] <=  8'h00;      memory[11265] <=  8'h00;      memory[11266] <=  8'h00;      memory[11267] <=  8'h00;      memory[11268] <=  8'h00;      memory[11269] <=  8'h00;      memory[11270] <=  8'h00;      memory[11271] <=  8'h00;      memory[11272] <=  8'h00;      memory[11273] <=  8'h00;      memory[11274] <=  8'h00;      memory[11275] <=  8'h00;      memory[11276] <=  8'h00;      memory[11277] <=  8'h00;      memory[11278] <=  8'h00;      memory[11279] <=  8'h00;      memory[11280] <=  8'h00;      memory[11281] <=  8'h00;      memory[11282] <=  8'h00;      memory[11283] <=  8'h00;      memory[11284] <=  8'h00;      memory[11285] <=  8'h00;      memory[11286] <=  8'h00;      memory[11287] <=  8'h00;      memory[11288] <=  8'h00;      memory[11289] <=  8'h00;      memory[11290] <=  8'h00;      memory[11291] <=  8'h00;      memory[11292] <=  8'h00;      memory[11293] <=  8'h00;      memory[11294] <=  8'h00;      memory[11295] <=  8'h00;      memory[11296] <=  8'h00;      memory[11297] <=  8'h00;      memory[11298] <=  8'h00;      memory[11299] <=  8'h00;      memory[11300] <=  8'h00;      memory[11301] <=  8'h00;      memory[11302] <=  8'h00;      memory[11303] <=  8'h00;      memory[11304] <=  8'h00;      memory[11305] <=  8'h00;      memory[11306] <=  8'h00;      memory[11307] <=  8'h00;      memory[11308] <=  8'h00;      memory[11309] <=  8'h00;      memory[11310] <=  8'h00;      memory[11311] <=  8'h00;      memory[11312] <=  8'h00;      memory[11313] <=  8'h00;      memory[11314] <=  8'h00;      memory[11315] <=  8'h00;      memory[11316] <=  8'h00;      memory[11317] <=  8'h00;      memory[11318] <=  8'h00;      memory[11319] <=  8'h00;      memory[11320] <=  8'h00;      memory[11321] <=  8'h00;      memory[11322] <=  8'h00;      memory[11323] <=  8'h00;      memory[11324] <=  8'h00;      memory[11325] <=  8'h00;      memory[11326] <=  8'h00;      memory[11327] <=  8'h00;      memory[11328] <=  8'h00;      memory[11329] <=  8'h00;      memory[11330] <=  8'h00;      memory[11331] <=  8'h00;      memory[11332] <=  8'h00;      memory[11333] <=  8'h00;      memory[11334] <=  8'h00;      memory[11335] <=  8'h00;      memory[11336] <=  8'h00;      memory[11337] <=  8'h00;      memory[11338] <=  8'h00;      memory[11339] <=  8'h00;      memory[11340] <=  8'h00;      memory[11341] <=  8'h00;      memory[11342] <=  8'h00;      memory[11343] <=  8'h00;      memory[11344] <=  8'h00;      memory[11345] <=  8'h00;      memory[11346] <=  8'h00;      memory[11347] <=  8'h00;      memory[11348] <=  8'h00;      memory[11349] <=  8'h00;      memory[11350] <=  8'h00;      memory[11351] <=  8'h00;      memory[11352] <=  8'h00;      memory[11353] <=  8'h00;      memory[11354] <=  8'h00;      memory[11355] <=  8'h00;      memory[11356] <=  8'h00;      memory[11357] <=  8'h00;      memory[11358] <=  8'h00;      memory[11359] <=  8'h00;      memory[11360] <=  8'h00;      memory[11361] <=  8'h00;      memory[11362] <=  8'h00;      memory[11363] <=  8'h00;      memory[11364] <=  8'h00;      memory[11365] <=  8'h00;      memory[11366] <=  8'h00;      memory[11367] <=  8'h00;      memory[11368] <=  8'h00;      memory[11369] <=  8'h00;      memory[11370] <=  8'h00;      memory[11371] <=  8'h00;      memory[11372] <=  8'h00;      memory[11373] <=  8'h00;      memory[11374] <=  8'h00;      memory[11375] <=  8'h00;      memory[11376] <=  8'h00;      memory[11377] <=  8'h00;      memory[11378] <=  8'h00;      memory[11379] <=  8'h00;      memory[11380] <=  8'h00;      memory[11381] <=  8'h00;      memory[11382] <=  8'h00;      memory[11383] <=  8'h00;      memory[11384] <=  8'h00;      memory[11385] <=  8'h00;      memory[11386] <=  8'h00;      memory[11387] <=  8'h00;      memory[11388] <=  8'h00;      memory[11389] <=  8'h00;      memory[11390] <=  8'h00;      memory[11391] <=  8'h00;      memory[11392] <=  8'h00;      memory[11393] <=  8'h00;      memory[11394] <=  8'h00;      memory[11395] <=  8'h00;      memory[11396] <=  8'h00;      memory[11397] <=  8'h00;      memory[11398] <=  8'h00;      memory[11399] <=  8'h00;      memory[11400] <=  8'h00;      memory[11401] <=  8'h00;      memory[11402] <=  8'h00;      memory[11403] <=  8'h00;      memory[11404] <=  8'h00;      memory[11405] <=  8'h00;      memory[11406] <=  8'h00;      memory[11407] <=  8'h00;      memory[11408] <=  8'h00;      memory[11409] <=  8'h00;      memory[11410] <=  8'h00;      memory[11411] <=  8'h00;      memory[11412] <=  8'h00;      memory[11413] <=  8'h00;      memory[11414] <=  8'h00;      memory[11415] <=  8'h00;      memory[11416] <=  8'h00;      memory[11417] <=  8'h00;      memory[11418] <=  8'h00;      memory[11419] <=  8'h00;      memory[11420] <=  8'h00;      memory[11421] <=  8'h00;      memory[11422] <=  8'h00;      memory[11423] <=  8'h00;      memory[11424] <=  8'h00;      memory[11425] <=  8'h00;      memory[11426] <=  8'h00;      memory[11427] <=  8'h00;      memory[11428] <=  8'h00;      memory[11429] <=  8'h00;      memory[11430] <=  8'h00;      memory[11431] <=  8'h00;      memory[11432] <=  8'h00;      memory[11433] <=  8'h00;      memory[11434] <=  8'h00;      memory[11435] <=  8'h00;      memory[11436] <=  8'h00;      memory[11437] <=  8'h00;      memory[11438] <=  8'h00;      memory[11439] <=  8'h00;      memory[11440] <=  8'h00;      memory[11441] <=  8'h00;      memory[11442] <=  8'h00;      memory[11443] <=  8'h00;      memory[11444] <=  8'h00;      memory[11445] <=  8'h00;      memory[11446] <=  8'h00;      memory[11447] <=  8'h00;      memory[11448] <=  8'h00;      memory[11449] <=  8'h00;      memory[11450] <=  8'h00;      memory[11451] <=  8'h00;      memory[11452] <=  8'h00;      memory[11453] <=  8'h00;      memory[11454] <=  8'h00;      memory[11455] <=  8'h00;      memory[11456] <=  8'h00;      memory[11457] <=  8'h00;      memory[11458] <=  8'h00;      memory[11459] <=  8'h00;      memory[11460] <=  8'h00;      memory[11461] <=  8'h00;      memory[11462] <=  8'h00;      memory[11463] <=  8'h00;      memory[11464] <=  8'h00;      memory[11465] <=  8'h00;      memory[11466] <=  8'h00;      memory[11467] <=  8'h00;      memory[11468] <=  8'h00;      memory[11469] <=  8'h00;      memory[11470] <=  8'h00;      memory[11471] <=  8'h00;      memory[11472] <=  8'h00;      memory[11473] <=  8'h00;      memory[11474] <=  8'h00;      memory[11475] <=  8'h00;      memory[11476] <=  8'h00;      memory[11477] <=  8'h00;      memory[11478] <=  8'h00;      memory[11479] <=  8'h00;      memory[11480] <=  8'h00;      memory[11481] <=  8'h00;      memory[11482] <=  8'h00;      memory[11483] <=  8'h00;      memory[11484] <=  8'h00;      memory[11485] <=  8'h00;      memory[11486] <=  8'h00;      memory[11487] <=  8'h00;      memory[11488] <=  8'h00;      memory[11489] <=  8'h00;      memory[11490] <=  8'h00;      memory[11491] <=  8'h00;      memory[11492] <=  8'h00;      memory[11493] <=  8'h00;      memory[11494] <=  8'h00;      memory[11495] <=  8'h00;      memory[11496] <=  8'h00;      memory[11497] <=  8'h00;      memory[11498] <=  8'h00;      memory[11499] <=  8'h00;      memory[11500] <=  8'h00;      memory[11501] <=  8'h00;      memory[11502] <=  8'h00;      memory[11503] <=  8'h00;      memory[11504] <=  8'h00;      memory[11505] <=  8'h00;      memory[11506] <=  8'h00;      memory[11507] <=  8'h00;      memory[11508] <=  8'h00;      memory[11509] <=  8'h00;      memory[11510] <=  8'h00;      memory[11511] <=  8'h00;      memory[11512] <=  8'h00;      memory[11513] <=  8'h00;      memory[11514] <=  8'h00;      memory[11515] <=  8'h00;      memory[11516] <=  8'h00;      memory[11517] <=  8'h00;      memory[11518] <=  8'h00;      memory[11519] <=  8'h00;      memory[11520] <=  8'h00;      memory[11521] <=  8'h00;      memory[11522] <=  8'h00;      memory[11523] <=  8'h00;      memory[11524] <=  8'h00;      memory[11525] <=  8'h00;      memory[11526] <=  8'h00;      memory[11527] <=  8'h00;      memory[11528] <=  8'h00;      memory[11529] <=  8'h00;      memory[11530] <=  8'h00;      memory[11531] <=  8'h00;      memory[11532] <=  8'h00;      memory[11533] <=  8'h00;      memory[11534] <=  8'h00;      memory[11535] <=  8'h00;      memory[11536] <=  8'h00;      memory[11537] <=  8'h00;      memory[11538] <=  8'h00;      memory[11539] <=  8'h00;      memory[11540] <=  8'h00;      memory[11541] <=  8'h00;      memory[11542] <=  8'h00;      memory[11543] <=  8'h00;      memory[11544] <=  8'h00;      memory[11545] <=  8'h00;      memory[11546] <=  8'h00;      memory[11547] <=  8'h00;      memory[11548] <=  8'h00;      memory[11549] <=  8'h00;      memory[11550] <=  8'h00;      memory[11551] <=  8'h00;      memory[11552] <=  8'h00;      memory[11553] <=  8'h00;      memory[11554] <=  8'h00;      memory[11555] <=  8'h00;      memory[11556] <=  8'h00;      memory[11557] <=  8'h00;      memory[11558] <=  8'h00;      memory[11559] <=  8'h00;      memory[11560] <=  8'h00;      memory[11561] <=  8'h00;      memory[11562] <=  8'h00;      memory[11563] <=  8'h00;      memory[11564] <=  8'h00;      memory[11565] <=  8'h00;      memory[11566] <=  8'h00;      memory[11567] <=  8'h00;      memory[11568] <=  8'h00;      memory[11569] <=  8'h00;      memory[11570] <=  8'h00;      memory[11571] <=  8'h00;      memory[11572] <=  8'h00;      memory[11573] <=  8'h00;      memory[11574] <=  8'h00;      memory[11575] <=  8'h00;      memory[11576] <=  8'h00;      memory[11577] <=  8'h00;      memory[11578] <=  8'h00;      memory[11579] <=  8'h00;      memory[11580] <=  8'h00;      memory[11581] <=  8'h00;      memory[11582] <=  8'h00;      memory[11583] <=  8'h00;      memory[11584] <=  8'h00;      memory[11585] <=  8'h00;      memory[11586] <=  8'h00;      memory[11587] <=  8'h00;      memory[11588] <=  8'h00;      memory[11589] <=  8'h00;      memory[11590] <=  8'h00;      memory[11591] <=  8'h00;      memory[11592] <=  8'h00;      memory[11593] <=  8'h00;      memory[11594] <=  8'h00;      memory[11595] <=  8'h00;      memory[11596] <=  8'h00;      memory[11597] <=  8'h00;      memory[11598] <=  8'h00;      memory[11599] <=  8'h00;      memory[11600] <=  8'h00;      memory[11601] <=  8'h00;      memory[11602] <=  8'h00;      memory[11603] <=  8'h00;      memory[11604] <=  8'h00;      memory[11605] <=  8'h00;      memory[11606] <=  8'h00;      memory[11607] <=  8'h00;      memory[11608] <=  8'h00;      memory[11609] <=  8'h00;      memory[11610] <=  8'h00;      memory[11611] <=  8'h00;      memory[11612] <=  8'h00;      memory[11613] <=  8'h00;      memory[11614] <=  8'h00;      memory[11615] <=  8'h00;      memory[11616] <=  8'h00;      memory[11617] <=  8'h00;      memory[11618] <=  8'h00;      memory[11619] <=  8'h00;      memory[11620] <=  8'h00;      memory[11621] <=  8'h00;      memory[11622] <=  8'h00;      memory[11623] <=  8'h00;      memory[11624] <=  8'h00;      memory[11625] <=  8'h00;      memory[11626] <=  8'h00;      memory[11627] <=  8'h00;      memory[11628] <=  8'h00;      memory[11629] <=  8'h00;      memory[11630] <=  8'h00;      memory[11631] <=  8'h00;      memory[11632] <=  8'h00;      memory[11633] <=  8'h00;      memory[11634] <=  8'h00;      memory[11635] <=  8'h00;      memory[11636] <=  8'h00;      memory[11637] <=  8'h00;      memory[11638] <=  8'h00;      memory[11639] <=  8'h00;      memory[11640] <=  8'h00;      memory[11641] <=  8'h00;      memory[11642] <=  8'h00;      memory[11643] <=  8'h00;      memory[11644] <=  8'h00;      memory[11645] <=  8'h00;      memory[11646] <=  8'h00;      memory[11647] <=  8'h00;      memory[11648] <=  8'h00;      memory[11649] <=  8'h00;      memory[11650] <=  8'h00;      memory[11651] <=  8'h00;      memory[11652] <=  8'h00;      memory[11653] <=  8'h00;      memory[11654] <=  8'h00;      memory[11655] <=  8'h00;      memory[11656] <=  8'h00;      memory[11657] <=  8'h00;      memory[11658] <=  8'h00;      memory[11659] <=  8'h00;      memory[11660] <=  8'h00;      memory[11661] <=  8'h00;      memory[11662] <=  8'h00;      memory[11663] <=  8'h00;      memory[11664] <=  8'h00;      memory[11665] <=  8'h00;      memory[11666] <=  8'h00;      memory[11667] <=  8'h00;      memory[11668] <=  8'h00;      memory[11669] <=  8'h00;      memory[11670] <=  8'h00;      memory[11671] <=  8'h00;      memory[11672] <=  8'h00;      memory[11673] <=  8'h00;      memory[11674] <=  8'h00;      memory[11675] <=  8'h00;      memory[11676] <=  8'h00;      memory[11677] <=  8'h00;      memory[11678] <=  8'h00;      memory[11679] <=  8'h00;      memory[11680] <=  8'h00;      memory[11681] <=  8'h00;      memory[11682] <=  8'h00;      memory[11683] <=  8'h00;      memory[11684] <=  8'h00;      memory[11685] <=  8'h00;      memory[11686] <=  8'h00;      memory[11687] <=  8'h00;      memory[11688] <=  8'h00;      memory[11689] <=  8'h00;      memory[11690] <=  8'h00;      memory[11691] <=  8'h00;      memory[11692] <=  8'h00;      memory[11693] <=  8'h00;      memory[11694] <=  8'h00;      memory[11695] <=  8'h00;      memory[11696] <=  8'h00;      memory[11697] <=  8'h00;      memory[11698] <=  8'h00;      memory[11699] <=  8'h00;      memory[11700] <=  8'h00;      memory[11701] <=  8'h00;      memory[11702] <=  8'h00;      memory[11703] <=  8'h00;      memory[11704] <=  8'h00;      memory[11705] <=  8'h00;      memory[11706] <=  8'h00;      memory[11707] <=  8'h00;      memory[11708] <=  8'h00;      memory[11709] <=  8'h00;      memory[11710] <=  8'h00;      memory[11711] <=  8'h00;      memory[11712] <=  8'h00;      memory[11713] <=  8'h00;      memory[11714] <=  8'h00;      memory[11715] <=  8'h00;      memory[11716] <=  8'h00;      memory[11717] <=  8'h00;      memory[11718] <=  8'h00;      memory[11719] <=  8'h00;      memory[11720] <=  8'h00;      memory[11721] <=  8'h00;      memory[11722] <=  8'h00;      memory[11723] <=  8'h00;      memory[11724] <=  8'h00;      memory[11725] <=  8'h00;      memory[11726] <=  8'h00;      memory[11727] <=  8'h00;      memory[11728] <=  8'h00;      memory[11729] <=  8'h00;      memory[11730] <=  8'h00;      memory[11731] <=  8'h00;      memory[11732] <=  8'h00;      memory[11733] <=  8'h00;      memory[11734] <=  8'h00;      memory[11735] <=  8'h00;      memory[11736] <=  8'h00;      memory[11737] <=  8'h00;      memory[11738] <=  8'h00;      memory[11739] <=  8'h00;      memory[11740] <=  8'h00;      memory[11741] <=  8'h00;      memory[11742] <=  8'h00;      memory[11743] <=  8'h00;      memory[11744] <=  8'h00;      memory[11745] <=  8'h00;      memory[11746] <=  8'h00;      memory[11747] <=  8'h00;      memory[11748] <=  8'h00;      memory[11749] <=  8'h00;      memory[11750] <=  8'h00;      memory[11751] <=  8'h00;      memory[11752] <=  8'h00;      memory[11753] <=  8'h00;      memory[11754] <=  8'h00;      memory[11755] <=  8'h00;      memory[11756] <=  8'h00;      memory[11757] <=  8'h00;      memory[11758] <=  8'h00;      memory[11759] <=  8'h00;      memory[11760] <=  8'h00;      memory[11761] <=  8'h00;      memory[11762] <=  8'h00;      memory[11763] <=  8'h00;      memory[11764] <=  8'h00;      memory[11765] <=  8'h00;      memory[11766] <=  8'h00;      memory[11767] <=  8'h00;      memory[11768] <=  8'h00;      memory[11769] <=  8'h00;      memory[11770] <=  8'h00;      memory[11771] <=  8'h00;      memory[11772] <=  8'h00;      memory[11773] <=  8'h00;      memory[11774] <=  8'h00;      memory[11775] <=  8'h00;      memory[11776] <=  8'h00;      memory[11777] <=  8'h00;      memory[11778] <=  8'h00;      memory[11779] <=  8'h00;      memory[11780] <=  8'h00;      memory[11781] <=  8'h00;      memory[11782] <=  8'h00;      memory[11783] <=  8'h00;      memory[11784] <=  8'h00;      memory[11785] <=  8'h00;      memory[11786] <=  8'h00;      memory[11787] <=  8'h00;      memory[11788] <=  8'h00;      memory[11789] <=  8'h00;      memory[11790] <=  8'h00;      memory[11791] <=  8'h00;      memory[11792] <=  8'h00;      memory[11793] <=  8'h00;      memory[11794] <=  8'h00;      memory[11795] <=  8'h00;      memory[11796] <=  8'h00;      memory[11797] <=  8'h00;      memory[11798] <=  8'h00;      memory[11799] <=  8'h00;      memory[11800] <=  8'h00;      memory[11801] <=  8'h00;      memory[11802] <=  8'h00;      memory[11803] <=  8'h00;      memory[11804] <=  8'h00;      memory[11805] <=  8'h00;      memory[11806] <=  8'h00;      memory[11807] <=  8'h00;      memory[11808] <=  8'h00;      memory[11809] <=  8'h00;      memory[11810] <=  8'h00;      memory[11811] <=  8'h00;      memory[11812] <=  8'h00;      memory[11813] <=  8'h00;      memory[11814] <=  8'h00;      memory[11815] <=  8'h00;      memory[11816] <=  8'h00;      memory[11817] <=  8'h00;      memory[11818] <=  8'h00;      memory[11819] <=  8'h00;      memory[11820] <=  8'h00;      memory[11821] <=  8'h00;      memory[11822] <=  8'h00;      memory[11823] <=  8'h00;      memory[11824] <=  8'h00;      memory[11825] <=  8'h00;      memory[11826] <=  8'h00;      memory[11827] <=  8'h00;      memory[11828] <=  8'h00;      memory[11829] <=  8'h00;      memory[11830] <=  8'h00;      memory[11831] <=  8'h00;      memory[11832] <=  8'h00;      memory[11833] <=  8'h00;      memory[11834] <=  8'h00;      memory[11835] <=  8'h00;      memory[11836] <=  8'h00;      memory[11837] <=  8'h00;      memory[11838] <=  8'h00;      memory[11839] <=  8'h00;      memory[11840] <=  8'h00;      memory[11841] <=  8'h00;      memory[11842] <=  8'h00;      memory[11843] <=  8'h00;      memory[11844] <=  8'h00;      memory[11845] <=  8'h00;      memory[11846] <=  8'h00;      memory[11847] <=  8'h00;      memory[11848] <=  8'h00;      memory[11849] <=  8'h00;      memory[11850] <=  8'h00;      memory[11851] <=  8'h00;      memory[11852] <=  8'h00;      memory[11853] <=  8'h00;      memory[11854] <=  8'h00;      memory[11855] <=  8'h00;      memory[11856] <=  8'h00;      memory[11857] <=  8'h00;      memory[11858] <=  8'h00;      memory[11859] <=  8'h00;      memory[11860] <=  8'h00;      memory[11861] <=  8'h00;      memory[11862] <=  8'h00;      memory[11863] <=  8'h00;      memory[11864] <=  8'h00;      memory[11865] <=  8'h00;      memory[11866] <=  8'h00;      memory[11867] <=  8'h00;      memory[11868] <=  8'h00;      memory[11869] <=  8'h00;      memory[11870] <=  8'h00;      memory[11871] <=  8'h00;      memory[11872] <=  8'h00;      memory[11873] <=  8'h00;      memory[11874] <=  8'h00;      memory[11875] <=  8'h00;      memory[11876] <=  8'h00;      memory[11877] <=  8'h00;      memory[11878] <=  8'h00;      memory[11879] <=  8'h00;      memory[11880] <=  8'h00;      memory[11881] <=  8'h00;      memory[11882] <=  8'h00;      memory[11883] <=  8'h00;      memory[11884] <=  8'h00;      memory[11885] <=  8'h00;      memory[11886] <=  8'h00;      memory[11887] <=  8'h00;      memory[11888] <=  8'h00;      memory[11889] <=  8'h00;      memory[11890] <=  8'h00;      memory[11891] <=  8'h00;      memory[11892] <=  8'h00;      memory[11893] <=  8'h00;      memory[11894] <=  8'h00;      memory[11895] <=  8'h00;      memory[11896] <=  8'h00;      memory[11897] <=  8'h00;      memory[11898] <=  8'h00;      memory[11899] <=  8'h00;      memory[11900] <=  8'h00;      memory[11901] <=  8'h00;      memory[11902] <=  8'h00;      memory[11903] <=  8'h00;      memory[11904] <=  8'h00;      memory[11905] <=  8'h00;      memory[11906] <=  8'h00;      memory[11907] <=  8'h00;      memory[11908] <=  8'h00;      memory[11909] <=  8'h00;      memory[11910] <=  8'h00;      memory[11911] <=  8'h00;      memory[11912] <=  8'h00;      memory[11913] <=  8'h00;      memory[11914] <=  8'h00;      memory[11915] <=  8'h00;      memory[11916] <=  8'h00;      memory[11917] <=  8'h00;      memory[11918] <=  8'h00;      memory[11919] <=  8'h00;      memory[11920] <=  8'h00;      memory[11921] <=  8'h00;      memory[11922] <=  8'h00;      memory[11923] <=  8'h00;      memory[11924] <=  8'h00;      memory[11925] <=  8'h00;      memory[11926] <=  8'h00;      memory[11927] <=  8'h00;      memory[11928] <=  8'h00;      memory[11929] <=  8'h00;      memory[11930] <=  8'h00;      memory[11931] <=  8'h00;      memory[11932] <=  8'h00;      memory[11933] <=  8'h00;      memory[11934] <=  8'h00;      memory[11935] <=  8'h00;      memory[11936] <=  8'h00;      memory[11937] <=  8'h00;      memory[11938] <=  8'h00;      memory[11939] <=  8'h00;      memory[11940] <=  8'h00;      memory[11941] <=  8'h00;      memory[11942] <=  8'h00;      memory[11943] <=  8'h00;      memory[11944] <=  8'h00;      memory[11945] <=  8'h00;      memory[11946] <=  8'h00;      memory[11947] <=  8'h00;      memory[11948] <=  8'h00;      memory[11949] <=  8'h00;      memory[11950] <=  8'h00;      memory[11951] <=  8'h00;      memory[11952] <=  8'h00;      memory[11953] <=  8'h00;      memory[11954] <=  8'h00;      memory[11955] <=  8'h00;      memory[11956] <=  8'h00;      memory[11957] <=  8'h00;      memory[11958] <=  8'h00;      memory[11959] <=  8'h00;      memory[11960] <=  8'h00;      memory[11961] <=  8'h00;      memory[11962] <=  8'h00;      memory[11963] <=  8'h00;      memory[11964] <=  8'h00;      memory[11965] <=  8'h00;      memory[11966] <=  8'h00;      memory[11967] <=  8'h00;      memory[11968] <=  8'h00;      memory[11969] <=  8'h00;      memory[11970] <=  8'h00;      memory[11971] <=  8'h00;      memory[11972] <=  8'h00;      memory[11973] <=  8'h00;      memory[11974] <=  8'h00;      memory[11975] <=  8'h00;      memory[11976] <=  8'h00;      memory[11977] <=  8'h00;      memory[11978] <=  8'h00;      memory[11979] <=  8'h00;      memory[11980] <=  8'h00;      memory[11981] <=  8'h00;      memory[11982] <=  8'h00;      memory[11983] <=  8'h00;      memory[11984] <=  8'h00;      memory[11985] <=  8'h00;      memory[11986] <=  8'h00;      memory[11987] <=  8'h00;      memory[11988] <=  8'h00;      memory[11989] <=  8'h00;      memory[11990] <=  8'h00;      memory[11991] <=  8'h00;      memory[11992] <=  8'h00;      memory[11993] <=  8'h00;      memory[11994] <=  8'h00;      memory[11995] <=  8'h00;      memory[11996] <=  8'h00;      memory[11997] <=  8'h00;      memory[11998] <=  8'h00;      memory[11999] <=  8'h00;      memory[12000] <=  8'h00;      memory[12001] <=  8'h00;      memory[12002] <=  8'h00;      memory[12003] <=  8'h00;      memory[12004] <=  8'h00;      memory[12005] <=  8'h00;      memory[12006] <=  8'h00;      memory[12007] <=  8'h00;      memory[12008] <=  8'h00;      memory[12009] <=  8'h00;      memory[12010] <=  8'h00;      memory[12011] <=  8'h00;      memory[12012] <=  8'h00;      memory[12013] <=  8'h00;      memory[12014] <=  8'h00;      memory[12015] <=  8'h00;      memory[12016] <=  8'h00;      memory[12017] <=  8'h00;      memory[12018] <=  8'h00;      memory[12019] <=  8'h00;      memory[12020] <=  8'h00;      memory[12021] <=  8'h00;      memory[12022] <=  8'h00;      memory[12023] <=  8'h00;      memory[12024] <=  8'h00;      memory[12025] <=  8'h00;      memory[12026] <=  8'h00;      memory[12027] <=  8'h00;      memory[12028] <=  8'h00;      memory[12029] <=  8'h00;      memory[12030] <=  8'h00;      memory[12031] <=  8'h00;      memory[12032] <=  8'h00;      memory[12033] <=  8'h00;      memory[12034] <=  8'h00;      memory[12035] <=  8'h00;      memory[12036] <=  8'h00;      memory[12037] <=  8'h00;      memory[12038] <=  8'h00;      memory[12039] <=  8'h00;      memory[12040] <=  8'h00;      memory[12041] <=  8'h00;      memory[12042] <=  8'h00;      memory[12043] <=  8'h00;      memory[12044] <=  8'h00;      memory[12045] <=  8'h00;      memory[12046] <=  8'h00;      memory[12047] <=  8'h00;      memory[12048] <=  8'h00;      memory[12049] <=  8'h00;      memory[12050] <=  8'h00;      memory[12051] <=  8'h00;      memory[12052] <=  8'h00;      memory[12053] <=  8'h00;      memory[12054] <=  8'h00;      memory[12055] <=  8'h00;      memory[12056] <=  8'h00;      memory[12057] <=  8'h00;      memory[12058] <=  8'h00;      memory[12059] <=  8'h00;      memory[12060] <=  8'h00;      memory[12061] <=  8'h00;      memory[12062] <=  8'h00;      memory[12063] <=  8'h00;      memory[12064] <=  8'h00;      memory[12065] <=  8'h00;      memory[12066] <=  8'h00;      memory[12067] <=  8'h00;      memory[12068] <=  8'h00;      memory[12069] <=  8'h00;      memory[12070] <=  8'h00;      memory[12071] <=  8'h00;      memory[12072] <=  8'h00;      memory[12073] <=  8'h00;      memory[12074] <=  8'h00;      memory[12075] <=  8'h00;      memory[12076] <=  8'h00;      memory[12077] <=  8'h00;      memory[12078] <=  8'h00;      memory[12079] <=  8'h00;      memory[12080] <=  8'h00;      memory[12081] <=  8'h00;      memory[12082] <=  8'h00;      memory[12083] <=  8'h00;      memory[12084] <=  8'h00;      memory[12085] <=  8'h00;      memory[12086] <=  8'h00;      memory[12087] <=  8'h00;      memory[12088] <=  8'h00;      memory[12089] <=  8'h00;      memory[12090] <=  8'h00;      memory[12091] <=  8'h00;      memory[12092] <=  8'h00;      memory[12093] <=  8'h00;      memory[12094] <=  8'h00;      memory[12095] <=  8'h00;      memory[12096] <=  8'h00;      memory[12097] <=  8'h00;      memory[12098] <=  8'h00;      memory[12099] <=  8'h00;      memory[12100] <=  8'h00;      memory[12101] <=  8'h00;      memory[12102] <=  8'h00;      memory[12103] <=  8'h00;      memory[12104] <=  8'h00;      memory[12105] <=  8'h00;      memory[12106] <=  8'h00;      memory[12107] <=  8'h00;      memory[12108] <=  8'h00;      memory[12109] <=  8'h00;      memory[12110] <=  8'h00;      memory[12111] <=  8'h00;      memory[12112] <=  8'h00;      memory[12113] <=  8'h00;      memory[12114] <=  8'h00;      memory[12115] <=  8'h00;      memory[12116] <=  8'h00;      memory[12117] <=  8'h00;      memory[12118] <=  8'h00;      memory[12119] <=  8'h00;      memory[12120] <=  8'h00;      memory[12121] <=  8'h00;      memory[12122] <=  8'h00;      memory[12123] <=  8'h00;      memory[12124] <=  8'h00;      memory[12125] <=  8'h00;      memory[12126] <=  8'h00;      memory[12127] <=  8'h00;      memory[12128] <=  8'h00;      memory[12129] <=  8'h00;      memory[12130] <=  8'h00;      memory[12131] <=  8'h00;      memory[12132] <=  8'h00;      memory[12133] <=  8'h00;      memory[12134] <=  8'h00;      memory[12135] <=  8'h00;      memory[12136] <=  8'h00;      memory[12137] <=  8'h00;      memory[12138] <=  8'h00;      memory[12139] <=  8'h00;      memory[12140] <=  8'h00;      memory[12141] <=  8'h00;      memory[12142] <=  8'h00;      memory[12143] <=  8'h00;      memory[12144] <=  8'h00;      memory[12145] <=  8'h00;      memory[12146] <=  8'h00;      memory[12147] <=  8'h00;      memory[12148] <=  8'h00;      memory[12149] <=  8'h00;      memory[12150] <=  8'h00;      memory[12151] <=  8'h00;      memory[12152] <=  8'h00;      memory[12153] <=  8'h00;      memory[12154] <=  8'h00;      memory[12155] <=  8'h00;      memory[12156] <=  8'h00;      memory[12157] <=  8'h00;      memory[12158] <=  8'h00;      memory[12159] <=  8'h00;      memory[12160] <=  8'h00;      memory[12161] <=  8'h00;      memory[12162] <=  8'h00;      memory[12163] <=  8'h00;      memory[12164] <=  8'h00;      memory[12165] <=  8'h00;      memory[12166] <=  8'h00;      memory[12167] <=  8'h00;      memory[12168] <=  8'h00;      memory[12169] <=  8'h00;      memory[12170] <=  8'h00;      memory[12171] <=  8'h00;      memory[12172] <=  8'h00;      memory[12173] <=  8'h00;      memory[12174] <=  8'h00;      memory[12175] <=  8'h00;      memory[12176] <=  8'h00;      memory[12177] <=  8'h00;      memory[12178] <=  8'h00;      memory[12179] <=  8'h00;      memory[12180] <=  8'h00;      memory[12181] <=  8'h00;      memory[12182] <=  8'h00;      memory[12183] <=  8'h00;      memory[12184] <=  8'h00;      memory[12185] <=  8'h00;      memory[12186] <=  8'h00;      memory[12187] <=  8'h00;      memory[12188] <=  8'h00;      memory[12189] <=  8'h00;      memory[12190] <=  8'h00;      memory[12191] <=  8'h00;      memory[12192] <=  8'h00;      memory[12193] <=  8'h00;      memory[12194] <=  8'h00;      memory[12195] <=  8'h00;      memory[12196] <=  8'h00;      memory[12197] <=  8'h00;      memory[12198] <=  8'h00;      memory[12199] <=  8'h00;      memory[12200] <=  8'h00;      memory[12201] <=  8'h00;      memory[12202] <=  8'h00;      memory[12203] <=  8'h00;      memory[12204] <=  8'h00;      memory[12205] <=  8'h00;      memory[12206] <=  8'h00;      memory[12207] <=  8'h00;      memory[12208] <=  8'h00;      memory[12209] <=  8'h00;      memory[12210] <=  8'h00;      memory[12211] <=  8'h00;      memory[12212] <=  8'h00;      memory[12213] <=  8'h00;      memory[12214] <=  8'h00;      memory[12215] <=  8'h00;      memory[12216] <=  8'h00;      memory[12217] <=  8'h00;      memory[12218] <=  8'h00;      memory[12219] <=  8'h00;      memory[12220] <=  8'h00;      memory[12221] <=  8'h00;      memory[12222] <=  8'h00;      memory[12223] <=  8'h00;      memory[12224] <=  8'h00;      memory[12225] <=  8'h00;      memory[12226] <=  8'h00;      memory[12227] <=  8'h00;      memory[12228] <=  8'h00;      memory[12229] <=  8'h00;      memory[12230] <=  8'h00;      memory[12231] <=  8'h00;      memory[12232] <=  8'h00;      memory[12233] <=  8'h00;      memory[12234] <=  8'h00;      memory[12235] <=  8'h00;      memory[12236] <=  8'h00;      memory[12237] <=  8'h00;      memory[12238] <=  8'h00;      memory[12239] <=  8'h00;      memory[12240] <=  8'h00;      memory[12241] <=  8'h00;      memory[12242] <=  8'h00;      memory[12243] <=  8'h00;      memory[12244] <=  8'h00;      memory[12245] <=  8'h00;      memory[12246] <=  8'h00;      memory[12247] <=  8'h00;      memory[12248] <=  8'h00;      memory[12249] <=  8'h00;      memory[12250] <=  8'h00;      memory[12251] <=  8'h00;      memory[12252] <=  8'h00;      memory[12253] <=  8'h00;      memory[12254] <=  8'h00;      memory[12255] <=  8'h00;      memory[12256] <=  8'h00;      memory[12257] <=  8'h00;      memory[12258] <=  8'h00;      memory[12259] <=  8'h00;      memory[12260] <=  8'h00;      memory[12261] <=  8'h00;      memory[12262] <=  8'h00;      memory[12263] <=  8'h00;      memory[12264] <=  8'h00;      memory[12265] <=  8'h00;      memory[12266] <=  8'h00;      memory[12267] <=  8'h00;      memory[12268] <=  8'h00;      memory[12269] <=  8'h00;      memory[12270] <=  8'h00;      memory[12271] <=  8'h00;      memory[12272] <=  8'h00;      memory[12273] <=  8'h00;      memory[12274] <=  8'h00;      memory[12275] <=  8'h00;      memory[12276] <=  8'h00;      memory[12277] <=  8'h00;      memory[12278] <=  8'h00;      memory[12279] <=  8'h00;      memory[12280] <=  8'h00;      memory[12281] <=  8'h00;      memory[12282] <=  8'h00;      memory[12283] <=  8'h00;      memory[12284] <=  8'h00;      memory[12285] <=  8'h00;      memory[12286] <=  8'h00;      memory[12287] <=  8'h00;      memory[12288] <=  8'h00;      memory[12289] <=  8'h00;      memory[12290] <=  8'h00;      memory[12291] <=  8'h00;      memory[12292] <=  8'h00;      memory[12293] <=  8'h00;      memory[12294] <=  8'h00;      memory[12295] <=  8'h00;      memory[12296] <=  8'h00;      memory[12297] <=  8'h00;      memory[12298] <=  8'h00;      memory[12299] <=  8'h00;      memory[12300] <=  8'h00;      memory[12301] <=  8'h00;      memory[12302] <=  8'h00;      memory[12303] <=  8'h00;      memory[12304] <=  8'h00;      memory[12305] <=  8'h00;      memory[12306] <=  8'h00;      memory[12307] <=  8'h00;      memory[12308] <=  8'h00;      memory[12309] <=  8'h00;      memory[12310] <=  8'h00;      memory[12311] <=  8'h00;      memory[12312] <=  8'h00;      memory[12313] <=  8'h00;      memory[12314] <=  8'h00;      memory[12315] <=  8'h00;      memory[12316] <=  8'h00;      memory[12317] <=  8'h00;      memory[12318] <=  8'h00;      memory[12319] <=  8'h00;      memory[12320] <=  8'h00;      memory[12321] <=  8'h00;      memory[12322] <=  8'h00;      memory[12323] <=  8'h00;      memory[12324] <=  8'h00;      memory[12325] <=  8'h00;      memory[12326] <=  8'h00;      memory[12327] <=  8'h00;      memory[12328] <=  8'h00;      memory[12329] <=  8'h00;      memory[12330] <=  8'h00;      memory[12331] <=  8'h00;      memory[12332] <=  8'h00;      memory[12333] <=  8'h00;      memory[12334] <=  8'h00;      memory[12335] <=  8'h00;      memory[12336] <=  8'h00;      memory[12337] <=  8'h00;      memory[12338] <=  8'h00;      memory[12339] <=  8'h00;      memory[12340] <=  8'h00;      memory[12341] <=  8'h00;      memory[12342] <=  8'h00;      memory[12343] <=  8'h00;      memory[12344] <=  8'h00;      memory[12345] <=  8'h00;      memory[12346] <=  8'h00;      memory[12347] <=  8'h00;      memory[12348] <=  8'h00;      memory[12349] <=  8'h00;      memory[12350] <=  8'h00;      memory[12351] <=  8'h00;      memory[12352] <=  8'h00;      memory[12353] <=  8'h00;      memory[12354] <=  8'h00;      memory[12355] <=  8'h00;      memory[12356] <=  8'h00;      memory[12357] <=  8'h00;      memory[12358] <=  8'h00;      memory[12359] <=  8'h00;      memory[12360] <=  8'h00;      memory[12361] <=  8'h00;      memory[12362] <=  8'h00;      memory[12363] <=  8'h00;      memory[12364] <=  8'h00;      memory[12365] <=  8'h00;      memory[12366] <=  8'h00;      memory[12367] <=  8'h00;      memory[12368] <=  8'h00;      memory[12369] <=  8'h00;      memory[12370] <=  8'h00;      memory[12371] <=  8'h00;      memory[12372] <=  8'h00;      memory[12373] <=  8'h00;      memory[12374] <=  8'h00;      memory[12375] <=  8'h00;      memory[12376] <=  8'h00;      memory[12377] <=  8'h00;      memory[12378] <=  8'h00;      memory[12379] <=  8'h00;      memory[12380] <=  8'h00;      memory[12381] <=  8'h00;      memory[12382] <=  8'h00;      memory[12383] <=  8'h00;      memory[12384] <=  8'h00;      memory[12385] <=  8'h00;      memory[12386] <=  8'h00;      memory[12387] <=  8'h00;      memory[12388] <=  8'h00;      memory[12389] <=  8'h00;      memory[12390] <=  8'h00;      memory[12391] <=  8'h00;      memory[12392] <=  8'h00;      memory[12393] <=  8'h00;      memory[12394] <=  8'h00;      memory[12395] <=  8'h00;      memory[12396] <=  8'h00;      memory[12397] <=  8'h00;      memory[12398] <=  8'h00;      memory[12399] <=  8'h00;      memory[12400] <=  8'h00;      memory[12401] <=  8'h00;      memory[12402] <=  8'h00;      memory[12403] <=  8'h00;      memory[12404] <=  8'h00;      memory[12405] <=  8'h00;      memory[12406] <=  8'h00;      memory[12407] <=  8'h00;      memory[12408] <=  8'h00;      memory[12409] <=  8'h00;      memory[12410] <=  8'h00;      memory[12411] <=  8'h00;      memory[12412] <=  8'h00;      memory[12413] <=  8'h00;      memory[12414] <=  8'h00;      memory[12415] <=  8'h00;      memory[12416] <=  8'h00;      memory[12417] <=  8'h00;      memory[12418] <=  8'h00;      memory[12419] <=  8'h00;      memory[12420] <=  8'h00;      memory[12421] <=  8'h00;      memory[12422] <=  8'h00;      memory[12423] <=  8'h00;      memory[12424] <=  8'h00;      memory[12425] <=  8'h00;      memory[12426] <=  8'h00;      memory[12427] <=  8'h00;      memory[12428] <=  8'h00;      memory[12429] <=  8'h00;      memory[12430] <=  8'h00;      memory[12431] <=  8'h00;      memory[12432] <=  8'h00;      memory[12433] <=  8'h00;      memory[12434] <=  8'h00;      memory[12435] <=  8'h00;      memory[12436] <=  8'h00;      memory[12437] <=  8'h00;      memory[12438] <=  8'h00;      memory[12439] <=  8'h00;      memory[12440] <=  8'h00;      memory[12441] <=  8'h00;      memory[12442] <=  8'h00;      memory[12443] <=  8'h00;      memory[12444] <=  8'h00;      memory[12445] <=  8'h00;      memory[12446] <=  8'h00;      memory[12447] <=  8'h00;      memory[12448] <=  8'h00;      memory[12449] <=  8'h00;      memory[12450] <=  8'h00;      memory[12451] <=  8'h00;      memory[12452] <=  8'h00;      memory[12453] <=  8'h00;      memory[12454] <=  8'h00;      memory[12455] <=  8'h00;      memory[12456] <=  8'h00;      memory[12457] <=  8'h00;      memory[12458] <=  8'h00;      memory[12459] <=  8'h00;      memory[12460] <=  8'h00;      memory[12461] <=  8'h00;      memory[12462] <=  8'h00;      memory[12463] <=  8'h00;      memory[12464] <=  8'h00;      memory[12465] <=  8'h00;      memory[12466] <=  8'h00;      memory[12467] <=  8'h00;      memory[12468] <=  8'h00;      memory[12469] <=  8'h00;      memory[12470] <=  8'h00;      memory[12471] <=  8'h00;      memory[12472] <=  8'h00;      memory[12473] <=  8'h00;      memory[12474] <=  8'h00;      memory[12475] <=  8'h00;      memory[12476] <=  8'h00;      memory[12477] <=  8'h00;      memory[12478] <=  8'h00;      memory[12479] <=  8'h00;      memory[12480] <=  8'h00;      memory[12481] <=  8'h00;      memory[12482] <=  8'h00;      memory[12483] <=  8'h00;      memory[12484] <=  8'h00;      memory[12485] <=  8'h00;      memory[12486] <=  8'h00;      memory[12487] <=  8'h00;      memory[12488] <=  8'h00;      memory[12489] <=  8'h00;      memory[12490] <=  8'h00;      memory[12491] <=  8'h00;      memory[12492] <=  8'h00;      memory[12493] <=  8'h00;      memory[12494] <=  8'h00;      memory[12495] <=  8'h00;      memory[12496] <=  8'h00;      memory[12497] <=  8'h00;      memory[12498] <=  8'h00;      memory[12499] <=  8'h00;      memory[12500] <=  8'h00;      memory[12501] <=  8'h00;      memory[12502] <=  8'h00;      memory[12503] <=  8'h00;      memory[12504] <=  8'h00;      memory[12505] <=  8'h00;      memory[12506] <=  8'h00;      memory[12507] <=  8'h00;      memory[12508] <=  8'h00;      memory[12509] <=  8'h00;      memory[12510] <=  8'h00;      memory[12511] <=  8'h00;      memory[12512] <=  8'h00;      memory[12513] <=  8'h00;      memory[12514] <=  8'h00;      memory[12515] <=  8'h00;      memory[12516] <=  8'h00;      memory[12517] <=  8'h00;      memory[12518] <=  8'h00;      memory[12519] <=  8'h00;      memory[12520] <=  8'h00;      memory[12521] <=  8'h00;      memory[12522] <=  8'h00;      memory[12523] <=  8'h00;      memory[12524] <=  8'h00;      memory[12525] <=  8'h00;      memory[12526] <=  8'h00;      memory[12527] <=  8'h00;      memory[12528] <=  8'h00;      memory[12529] <=  8'h00;      memory[12530] <=  8'h00;      memory[12531] <=  8'h00;      memory[12532] <=  8'h00;      memory[12533] <=  8'h00;      memory[12534] <=  8'h00;      memory[12535] <=  8'h00;      memory[12536] <=  8'h00;      memory[12537] <=  8'h00;      memory[12538] <=  8'h00;      memory[12539] <=  8'h00;      memory[12540] <=  8'h00;      memory[12541] <=  8'h00;      memory[12542] <=  8'h00;      memory[12543] <=  8'h00;      memory[12544] <=  8'h00;      memory[12545] <=  8'h00;      memory[12546] <=  8'h00;      memory[12547] <=  8'h00;      memory[12548] <=  8'h00;      memory[12549] <=  8'h00;      memory[12550] <=  8'h00;      memory[12551] <=  8'h00;      memory[12552] <=  8'h00;      memory[12553] <=  8'h00;      memory[12554] <=  8'h00;      memory[12555] <=  8'h00;      memory[12556] <=  8'h00;      memory[12557] <=  8'h00;      memory[12558] <=  8'h00;      memory[12559] <=  8'h00;      memory[12560] <=  8'h00;      memory[12561] <=  8'h00;      memory[12562] <=  8'h00;      memory[12563] <=  8'h00;      memory[12564] <=  8'h00;      memory[12565] <=  8'h00;      memory[12566] <=  8'h00;      memory[12567] <=  8'h00;      memory[12568] <=  8'h00;      memory[12569] <=  8'h00;      memory[12570] <=  8'h00;      memory[12571] <=  8'h00;      memory[12572] <=  8'h00;      memory[12573] <=  8'h00;      memory[12574] <=  8'h00;      memory[12575] <=  8'h00;      memory[12576] <=  8'h00;      memory[12577] <=  8'h00;      memory[12578] <=  8'h00;      memory[12579] <=  8'h00;      memory[12580] <=  8'h00;      memory[12581] <=  8'h00;      memory[12582] <=  8'h00;      memory[12583] <=  8'h00;      memory[12584] <=  8'h00;      memory[12585] <=  8'h00;      memory[12586] <=  8'h00;      memory[12587] <=  8'h00;      memory[12588] <=  8'h00;      memory[12589] <=  8'h00;      memory[12590] <=  8'h00;      memory[12591] <=  8'h00;      memory[12592] <=  8'h00;      memory[12593] <=  8'h00;      memory[12594] <=  8'h00;      memory[12595] <=  8'h00;      memory[12596] <=  8'h00;      memory[12597] <=  8'h00;      memory[12598] <=  8'h00;      memory[12599] <=  8'h00;      memory[12600] <=  8'h00;      memory[12601] <=  8'h00;      memory[12602] <=  8'h00;      memory[12603] <=  8'h00;      memory[12604] <=  8'h00;      memory[12605] <=  8'h00;      memory[12606] <=  8'h00;      memory[12607] <=  8'h00;      memory[12608] <=  8'h00;      memory[12609] <=  8'h00;      memory[12610] <=  8'h00;      memory[12611] <=  8'h00;      memory[12612] <=  8'h00;      memory[12613] <=  8'h00;      memory[12614] <=  8'h00;      memory[12615] <=  8'h00;      memory[12616] <=  8'h00;      memory[12617] <=  8'h00;      memory[12618] <=  8'h00;      memory[12619] <=  8'h00;      memory[12620] <=  8'h00;      memory[12621] <=  8'h00;      memory[12622] <=  8'h00;      memory[12623] <=  8'h00;      memory[12624] <=  8'h00;      memory[12625] <=  8'h00;      memory[12626] <=  8'h00;      memory[12627] <=  8'h00;      memory[12628] <=  8'h00;      memory[12629] <=  8'h00;      memory[12630] <=  8'h00;      memory[12631] <=  8'h00;      memory[12632] <=  8'h00;      memory[12633] <=  8'h00;      memory[12634] <=  8'h00;      memory[12635] <=  8'h00;      memory[12636] <=  8'h00;      memory[12637] <=  8'h00;      memory[12638] <=  8'h00;      memory[12639] <=  8'h00;      memory[12640] <=  8'h00;      memory[12641] <=  8'h00;      memory[12642] <=  8'h00;      memory[12643] <=  8'h00;      memory[12644] <=  8'h00;      memory[12645] <=  8'h00;      memory[12646] <=  8'h00;      memory[12647] <=  8'h00;      memory[12648] <=  8'h00;      memory[12649] <=  8'h00;      memory[12650] <=  8'h00;      memory[12651] <=  8'h00;      memory[12652] <=  8'h00;      memory[12653] <=  8'h00;      memory[12654] <=  8'h00;      memory[12655] <=  8'h00;      memory[12656] <=  8'h00;      memory[12657] <=  8'h00;      memory[12658] <=  8'h00;      memory[12659] <=  8'h00;      memory[12660] <=  8'h00;      memory[12661] <=  8'h00;      memory[12662] <=  8'h00;      memory[12663] <=  8'h00;      memory[12664] <=  8'h00;      memory[12665] <=  8'h00;      memory[12666] <=  8'h00;      memory[12667] <=  8'h00;      memory[12668] <=  8'h00;      memory[12669] <=  8'h00;      memory[12670] <=  8'h00;      memory[12671] <=  8'h00;      memory[12672] <=  8'h00;      memory[12673] <=  8'h00;      memory[12674] <=  8'h00;      memory[12675] <=  8'h00;      memory[12676] <=  8'h00;      memory[12677] <=  8'h00;      memory[12678] <=  8'h00;      memory[12679] <=  8'h00;      memory[12680] <=  8'h00;      memory[12681] <=  8'h00;      memory[12682] <=  8'h00;      memory[12683] <=  8'h00;      memory[12684] <=  8'h00;      memory[12685] <=  8'h00;      memory[12686] <=  8'h00;      memory[12687] <=  8'h00;      memory[12688] <=  8'h00;      memory[12689] <=  8'h00;      memory[12690] <=  8'h00;      memory[12691] <=  8'h00;      memory[12692] <=  8'h00;      memory[12693] <=  8'h00;      memory[12694] <=  8'h00;      memory[12695] <=  8'h00;      memory[12696] <=  8'h00;      memory[12697] <=  8'h00;      memory[12698] <=  8'h00;      memory[12699] <=  8'h00;      memory[12700] <=  8'h00;      memory[12701] <=  8'h00;      memory[12702] <=  8'h00;      memory[12703] <=  8'h00;      memory[12704] <=  8'h00;      memory[12705] <=  8'h00;      memory[12706] <=  8'h00;      memory[12707] <=  8'h00;      memory[12708] <=  8'h00;      memory[12709] <=  8'h00;      memory[12710] <=  8'h00;      memory[12711] <=  8'h00;      memory[12712] <=  8'h00;      memory[12713] <=  8'h00;      memory[12714] <=  8'h00;      memory[12715] <=  8'h00;      memory[12716] <=  8'h00;      memory[12717] <=  8'h00;      memory[12718] <=  8'h00;      memory[12719] <=  8'h00;      memory[12720] <=  8'h00;      memory[12721] <=  8'h00;      memory[12722] <=  8'h00;      memory[12723] <=  8'h00;      memory[12724] <=  8'h00;      memory[12725] <=  8'h00;      memory[12726] <=  8'h00;      memory[12727] <=  8'h00;      memory[12728] <=  8'h00;      memory[12729] <=  8'h00;      memory[12730] <=  8'h00;      memory[12731] <=  8'h00;      memory[12732] <=  8'h00;      memory[12733] <=  8'h00;      memory[12734] <=  8'h00;      memory[12735] <=  8'h00;      memory[12736] <=  8'h00;      memory[12737] <=  8'h00;      memory[12738] <=  8'h00;      memory[12739] <=  8'h00;      memory[12740] <=  8'h00;      memory[12741] <=  8'h00;      memory[12742] <=  8'h00;      memory[12743] <=  8'h00;      memory[12744] <=  8'h00;      memory[12745] <=  8'h00;      memory[12746] <=  8'h00;      memory[12747] <=  8'h00;      memory[12748] <=  8'h00;      memory[12749] <=  8'h00;      memory[12750] <=  8'h00;      memory[12751] <=  8'h00;      memory[12752] <=  8'h00;      memory[12753] <=  8'h00;      memory[12754] <=  8'h00;      memory[12755] <=  8'h00;      memory[12756] <=  8'h00;      memory[12757] <=  8'h00;      memory[12758] <=  8'h00;      memory[12759] <=  8'h00;      memory[12760] <=  8'h00;      memory[12761] <=  8'h00;      memory[12762] <=  8'h00;      memory[12763] <=  8'h00;      memory[12764] <=  8'h00;      memory[12765] <=  8'h00;      memory[12766] <=  8'h00;      memory[12767] <=  8'h00;      memory[12768] <=  8'h00;      memory[12769] <=  8'h00;      memory[12770] <=  8'h00;      memory[12771] <=  8'h00;      memory[12772] <=  8'h00;      memory[12773] <=  8'h00;      memory[12774] <=  8'h00;      memory[12775] <=  8'h00;      memory[12776] <=  8'h00;      memory[12777] <=  8'h00;      memory[12778] <=  8'h00;      memory[12779] <=  8'h00;      memory[12780] <=  8'h00;      memory[12781] <=  8'h00;      memory[12782] <=  8'h00;      memory[12783] <=  8'h00;      memory[12784] <=  8'h00;      memory[12785] <=  8'h00;      memory[12786] <=  8'h00;      memory[12787] <=  8'h00;      memory[12788] <=  8'h00;      memory[12789] <=  8'h00;      memory[12790] <=  8'h00;      memory[12791] <=  8'h00;      memory[12792] <=  8'h00;      memory[12793] <=  8'h00;      memory[12794] <=  8'h00;      memory[12795] <=  8'h00;      memory[12796] <=  8'h00;      memory[12797] <=  8'h00;      memory[12798] <=  8'h00;      memory[12799] <=  8'h00;      memory[12800] <=  8'h00;      memory[12801] <=  8'h00;      memory[12802] <=  8'h00;      memory[12803] <=  8'h00;      memory[12804] <=  8'h00;      memory[12805] <=  8'h00;      memory[12806] <=  8'h00;      memory[12807] <=  8'h00;      memory[12808] <=  8'h00;      memory[12809] <=  8'h00;      memory[12810] <=  8'h00;      memory[12811] <=  8'h00;      memory[12812] <=  8'h00;      memory[12813] <=  8'h00;      memory[12814] <=  8'h00;      memory[12815] <=  8'h00;      memory[12816] <=  8'h00;      memory[12817] <=  8'h00;      memory[12818] <=  8'h00;      memory[12819] <=  8'h00;      memory[12820] <=  8'h00;      memory[12821] <=  8'h00;      memory[12822] <=  8'h00;      memory[12823] <=  8'h00;      memory[12824] <=  8'h00;      memory[12825] <=  8'h00;      memory[12826] <=  8'h00;      memory[12827] <=  8'h00;      memory[12828] <=  8'h00;      memory[12829] <=  8'h00;      memory[12830] <=  8'h00;      memory[12831] <=  8'h00;      memory[12832] <=  8'h00;      memory[12833] <=  8'h00;      memory[12834] <=  8'h00;      memory[12835] <=  8'h00;      memory[12836] <=  8'h00;      memory[12837] <=  8'h00;      memory[12838] <=  8'h00;      memory[12839] <=  8'h00;      memory[12840] <=  8'h00;      memory[12841] <=  8'h00;      memory[12842] <=  8'h00;      memory[12843] <=  8'h00;      memory[12844] <=  8'h00;      memory[12845] <=  8'h00;      memory[12846] <=  8'h00;      memory[12847] <=  8'h00;      memory[12848] <=  8'h00;      memory[12849] <=  8'h00;      memory[12850] <=  8'h00;      memory[12851] <=  8'h00;      memory[12852] <=  8'h00;      memory[12853] <=  8'h00;      memory[12854] <=  8'h00;      memory[12855] <=  8'h00;      memory[12856] <=  8'h00;      memory[12857] <=  8'h00;      memory[12858] <=  8'h00;      memory[12859] <=  8'h00;      memory[12860] <=  8'h00;      memory[12861] <=  8'h00;      memory[12862] <=  8'h00;      memory[12863] <=  8'h00;      memory[12864] <=  8'h00;      memory[12865] <=  8'h00;      memory[12866] <=  8'h00;      memory[12867] <=  8'h00;      memory[12868] <=  8'h00;      memory[12869] <=  8'h00;      memory[12870] <=  8'h00;      memory[12871] <=  8'h00;      memory[12872] <=  8'h00;      memory[12873] <=  8'h00;      memory[12874] <=  8'h00;      memory[12875] <=  8'h00;      memory[12876] <=  8'h00;      memory[12877] <=  8'h00;      memory[12878] <=  8'h00;      memory[12879] <=  8'h00;      memory[12880] <=  8'h00;      memory[12881] <=  8'h00;      memory[12882] <=  8'h00;      memory[12883] <=  8'h00;      memory[12884] <=  8'h00;      memory[12885] <=  8'h00;      memory[12886] <=  8'h00;      memory[12887] <=  8'h00;      memory[12888] <=  8'h00;      memory[12889] <=  8'h00;      memory[12890] <=  8'h00;      memory[12891] <=  8'h00;      memory[12892] <=  8'h00;      memory[12893] <=  8'h00;      memory[12894] <=  8'h00;      memory[12895] <=  8'h00;      memory[12896] <=  8'h00;      memory[12897] <=  8'h00;      memory[12898] <=  8'h00;      memory[12899] <=  8'h00;      memory[12900] <=  8'h00;      memory[12901] <=  8'h00;      memory[12902] <=  8'h00;      memory[12903] <=  8'h00;      memory[12904] <=  8'h00;      memory[12905] <=  8'h00;      memory[12906] <=  8'h00;      memory[12907] <=  8'h00;      memory[12908] <=  8'h00;      memory[12909] <=  8'h00;      memory[12910] <=  8'h00;      memory[12911] <=  8'h00;      memory[12912] <=  8'h00;      memory[12913] <=  8'h00;      memory[12914] <=  8'h00;      memory[12915] <=  8'h00;      memory[12916] <=  8'h00;      memory[12917] <=  8'h00;      memory[12918] <=  8'h00;      memory[12919] <=  8'h00;      memory[12920] <=  8'h00;      memory[12921] <=  8'h00;      memory[12922] <=  8'h00;      memory[12923] <=  8'h00;      memory[12924] <=  8'h00;      memory[12925] <=  8'h00;      memory[12926] <=  8'h00;      memory[12927] <=  8'h00;      memory[12928] <=  8'h00;      memory[12929] <=  8'h00;      memory[12930] <=  8'h00;      memory[12931] <=  8'h00;      memory[12932] <=  8'h00;      memory[12933] <=  8'h00;      memory[12934] <=  8'h00;      memory[12935] <=  8'h00;      memory[12936] <=  8'h00;      memory[12937] <=  8'h00;      memory[12938] <=  8'h00;      memory[12939] <=  8'h00;      memory[12940] <=  8'h00;      memory[12941] <=  8'h00;      memory[12942] <=  8'h00;      memory[12943] <=  8'h00;      memory[12944] <=  8'h00;      memory[12945] <=  8'h00;      memory[12946] <=  8'h00;      memory[12947] <=  8'h00;      memory[12948] <=  8'h00;      memory[12949] <=  8'h00;      memory[12950] <=  8'h00;      memory[12951] <=  8'h00;      memory[12952] <=  8'h00;      memory[12953] <=  8'h00;      memory[12954] <=  8'h00;      memory[12955] <=  8'h00;      memory[12956] <=  8'h00;      memory[12957] <=  8'h00;      memory[12958] <=  8'h00;      memory[12959] <=  8'h00;      memory[12960] <=  8'h00;      memory[12961] <=  8'h00;      memory[12962] <=  8'h00;      memory[12963] <=  8'h00;      memory[12964] <=  8'h00;      memory[12965] <=  8'h00;      memory[12966] <=  8'h00;      memory[12967] <=  8'h00;      memory[12968] <=  8'h00;      memory[12969] <=  8'h00;      memory[12970] <=  8'h00;      memory[12971] <=  8'h00;      memory[12972] <=  8'h00;      memory[12973] <=  8'h00;      memory[12974] <=  8'h00;      memory[12975] <=  8'h00;      memory[12976] <=  8'h00;      memory[12977] <=  8'h00;      memory[12978] <=  8'h00;      memory[12979] <=  8'h00;      memory[12980] <=  8'h00;      memory[12981] <=  8'h00;      memory[12982] <=  8'h00;      memory[12983] <=  8'h00;      memory[12984] <=  8'h00;      memory[12985] <=  8'h00;      memory[12986] <=  8'h00;      memory[12987] <=  8'h00;      memory[12988] <=  8'h00;      memory[12989] <=  8'h00;      memory[12990] <=  8'h00;      memory[12991] <=  8'h00;      memory[12992] <=  8'h00;      memory[12993] <=  8'h00;      memory[12994] <=  8'h00;      memory[12995] <=  8'h00;      memory[12996] <=  8'h00;      memory[12997] <=  8'h00;      memory[12998] <=  8'h00;      memory[12999] <=  8'h00;      memory[13000] <=  8'h00;      memory[13001] <=  8'h00;      memory[13002] <=  8'h00;      memory[13003] <=  8'h00;      memory[13004] <=  8'h00;      memory[13005] <=  8'h00;      memory[13006] <=  8'h00;      memory[13007] <=  8'h00;      memory[13008] <=  8'h00;      memory[13009] <=  8'h00;      memory[13010] <=  8'h00;      memory[13011] <=  8'h00;      memory[13012] <=  8'h00;      memory[13013] <=  8'h00;      memory[13014] <=  8'h00;      memory[13015] <=  8'h00;      memory[13016] <=  8'h00;      memory[13017] <=  8'h00;      memory[13018] <=  8'h00;      memory[13019] <=  8'h00;      memory[13020] <=  8'h00;      memory[13021] <=  8'h00;      memory[13022] <=  8'h00;      memory[13023] <=  8'h00;      memory[13024] <=  8'h00;      memory[13025] <=  8'h00;      memory[13026] <=  8'h00;      memory[13027] <=  8'h00;      memory[13028] <=  8'h00;      memory[13029] <=  8'h00;      memory[13030] <=  8'h00;      memory[13031] <=  8'h00;      memory[13032] <=  8'h00;      memory[13033] <=  8'h00;      memory[13034] <=  8'h00;      memory[13035] <=  8'h00;      memory[13036] <=  8'h00;      memory[13037] <=  8'h00;      memory[13038] <=  8'h00;      memory[13039] <=  8'h00;      memory[13040] <=  8'h00;      memory[13041] <=  8'h00;      memory[13042] <=  8'h00;      memory[13043] <=  8'h00;      memory[13044] <=  8'h00;      memory[13045] <=  8'h00;      memory[13046] <=  8'h00;      memory[13047] <=  8'h00;      memory[13048] <=  8'h00;      memory[13049] <=  8'h00;      memory[13050] <=  8'h00;      memory[13051] <=  8'h00;      memory[13052] <=  8'h00;      memory[13053] <=  8'h00;      memory[13054] <=  8'h00;      memory[13055] <=  8'h00;      memory[13056] <=  8'h00;      memory[13057] <=  8'h00;      memory[13058] <=  8'h00;      memory[13059] <=  8'h00;      memory[13060] <=  8'h00;      memory[13061] <=  8'h00;      memory[13062] <=  8'h00;      memory[13063] <=  8'h00;      memory[13064] <=  8'h00;      memory[13065] <=  8'h00;      memory[13066] <=  8'h00;      memory[13067] <=  8'h00;      memory[13068] <=  8'h00;      memory[13069] <=  8'h00;      memory[13070] <=  8'h00;      memory[13071] <=  8'h00;      memory[13072] <=  8'h00;      memory[13073] <=  8'h00;      memory[13074] <=  8'h00;      memory[13075] <=  8'h00;      memory[13076] <=  8'h00;      memory[13077] <=  8'h00;      memory[13078] <=  8'h00;      memory[13079] <=  8'h00;      memory[13080] <=  8'h00;      memory[13081] <=  8'h00;      memory[13082] <=  8'h00;      memory[13083] <=  8'h00;      memory[13084] <=  8'h00;      memory[13085] <=  8'h00;      memory[13086] <=  8'h00;      memory[13087] <=  8'h00;      memory[13088] <=  8'h00;      memory[13089] <=  8'h00;      memory[13090] <=  8'h00;      memory[13091] <=  8'h00;      memory[13092] <=  8'h00;      memory[13093] <=  8'h00;      memory[13094] <=  8'h00;      memory[13095] <=  8'h00;      memory[13096] <=  8'h00;      memory[13097] <=  8'h00;      memory[13098] <=  8'h00;      memory[13099] <=  8'h00;      memory[13100] <=  8'h00;      memory[13101] <=  8'h00;      memory[13102] <=  8'h00;      memory[13103] <=  8'h00;      memory[13104] <=  8'h00;      memory[13105] <=  8'h00;      memory[13106] <=  8'h00;      memory[13107] <=  8'h00;      memory[13108] <=  8'h00;      memory[13109] <=  8'h00;      memory[13110] <=  8'h00;      memory[13111] <=  8'h00;      memory[13112] <=  8'h00;      memory[13113] <=  8'h00;      memory[13114] <=  8'h00;      memory[13115] <=  8'h00;      memory[13116] <=  8'h00;      memory[13117] <=  8'h00;      memory[13118] <=  8'h00;      memory[13119] <=  8'h00;      memory[13120] <=  8'h00;      memory[13121] <=  8'h00;      memory[13122] <=  8'h00;      memory[13123] <=  8'h00;      memory[13124] <=  8'h00;      memory[13125] <=  8'h00;      memory[13126] <=  8'h00;      memory[13127] <=  8'h00;      memory[13128] <=  8'h00;      memory[13129] <=  8'h00;      memory[13130] <=  8'h00;      memory[13131] <=  8'h00;      memory[13132] <=  8'h00;      memory[13133] <=  8'h00;      memory[13134] <=  8'h00;      memory[13135] <=  8'h00;      memory[13136] <=  8'h00;      memory[13137] <=  8'h00;      memory[13138] <=  8'h00;      memory[13139] <=  8'h00;      memory[13140] <=  8'h00;      memory[13141] <=  8'h00;      memory[13142] <=  8'h00;      memory[13143] <=  8'h00;      memory[13144] <=  8'h00;      memory[13145] <=  8'h00;      memory[13146] <=  8'h00;      memory[13147] <=  8'h00;      memory[13148] <=  8'h00;      memory[13149] <=  8'h00;      memory[13150] <=  8'h00;      memory[13151] <=  8'h00;      memory[13152] <=  8'h00;      memory[13153] <=  8'h00;      memory[13154] <=  8'h00;      memory[13155] <=  8'h00;      memory[13156] <=  8'h00;      memory[13157] <=  8'h00;      memory[13158] <=  8'h00;      memory[13159] <=  8'h00;      memory[13160] <=  8'h00;      memory[13161] <=  8'h00;      memory[13162] <=  8'h00;      memory[13163] <=  8'h00;      memory[13164] <=  8'h00;      memory[13165] <=  8'h00;      memory[13166] <=  8'h00;      memory[13167] <=  8'h00;      memory[13168] <=  8'h00;      memory[13169] <=  8'h00;      memory[13170] <=  8'h00;      memory[13171] <=  8'h00;      memory[13172] <=  8'h00;      memory[13173] <=  8'h00;      memory[13174] <=  8'h00;      memory[13175] <=  8'h00;      memory[13176] <=  8'h00;      memory[13177] <=  8'h00;      memory[13178] <=  8'h00;      memory[13179] <=  8'h00;      memory[13180] <=  8'h00;      memory[13181] <=  8'h00;      memory[13182] <=  8'h00;      memory[13183] <=  8'h00;      memory[13184] <=  8'h00;      memory[13185] <=  8'h00;      memory[13186] <=  8'h00;      memory[13187] <=  8'h00;      memory[13188] <=  8'h00;      memory[13189] <=  8'h00;      memory[13190] <=  8'h00;      memory[13191] <=  8'h00;      memory[13192] <=  8'h00;      memory[13193] <=  8'h00;      memory[13194] <=  8'h00;      memory[13195] <=  8'h00;      memory[13196] <=  8'h00;      memory[13197] <=  8'h00;      memory[13198] <=  8'h00;      memory[13199] <=  8'h00;      memory[13200] <=  8'h00;      memory[13201] <=  8'h00;      memory[13202] <=  8'h00;      memory[13203] <=  8'h00;      memory[13204] <=  8'h00;      memory[13205] <=  8'h00;      memory[13206] <=  8'h00;      memory[13207] <=  8'h00;      memory[13208] <=  8'h00;      memory[13209] <=  8'h00;      memory[13210] <=  8'h00;      memory[13211] <=  8'h00;      memory[13212] <=  8'h00;      memory[13213] <=  8'h00;      memory[13214] <=  8'h00;      memory[13215] <=  8'h00;      memory[13216] <=  8'h00;      memory[13217] <=  8'h00;      memory[13218] <=  8'h00;      memory[13219] <=  8'h00;      memory[13220] <=  8'h00;      memory[13221] <=  8'h00;      memory[13222] <=  8'h00;      memory[13223] <=  8'h00;      memory[13224] <=  8'h00;      memory[13225] <=  8'h00;      memory[13226] <=  8'h00;      memory[13227] <=  8'h00;      memory[13228] <=  8'h00;      memory[13229] <=  8'h00;      memory[13230] <=  8'h00;      memory[13231] <=  8'h00;      memory[13232] <=  8'h00;      memory[13233] <=  8'h00;      memory[13234] <=  8'h00;      memory[13235] <=  8'h00;      memory[13236] <=  8'h00;      memory[13237] <=  8'h00;      memory[13238] <=  8'h00;      memory[13239] <=  8'h00;      memory[13240] <=  8'h00;      memory[13241] <=  8'h00;      memory[13242] <=  8'h00;      memory[13243] <=  8'h00;      memory[13244] <=  8'h00;      memory[13245] <=  8'h00;      memory[13246] <=  8'h00;      memory[13247] <=  8'h00;      memory[13248] <=  8'h00;      memory[13249] <=  8'h00;      memory[13250] <=  8'h00;      memory[13251] <=  8'h00;      memory[13252] <=  8'h00;      memory[13253] <=  8'h00;      memory[13254] <=  8'h00;      memory[13255] <=  8'h00;      memory[13256] <=  8'h00;      memory[13257] <=  8'h00;      memory[13258] <=  8'h00;      memory[13259] <=  8'h00;      memory[13260] <=  8'h00;      memory[13261] <=  8'h00;      memory[13262] <=  8'h00;      memory[13263] <=  8'h00;      memory[13264] <=  8'h00;      memory[13265] <=  8'h00;      memory[13266] <=  8'h00;      memory[13267] <=  8'h00;      memory[13268] <=  8'h00;      memory[13269] <=  8'h00;      memory[13270] <=  8'h00;      memory[13271] <=  8'h00;      memory[13272] <=  8'h00;      memory[13273] <=  8'h00;      memory[13274] <=  8'h00;      memory[13275] <=  8'h00;      memory[13276] <=  8'h00;      memory[13277] <=  8'h00;      memory[13278] <=  8'h00;      memory[13279] <=  8'h00;      memory[13280] <=  8'h00;      memory[13281] <=  8'h00;      memory[13282] <=  8'h00;      memory[13283] <=  8'h00;      memory[13284] <=  8'h00;      memory[13285] <=  8'h00;      memory[13286] <=  8'h00;      memory[13287] <=  8'h00;      memory[13288] <=  8'h00;      memory[13289] <=  8'h00;      memory[13290] <=  8'h00;      memory[13291] <=  8'h00;      memory[13292] <=  8'h00;      memory[13293] <=  8'h00;      memory[13294] <=  8'h00;      memory[13295] <=  8'h00;      memory[13296] <=  8'h00;      memory[13297] <=  8'h00;      memory[13298] <=  8'h00;      memory[13299] <=  8'h00;      memory[13300] <=  8'h00;      memory[13301] <=  8'h00;      memory[13302] <=  8'h00;      memory[13303] <=  8'h00;      memory[13304] <=  8'h00;      memory[13305] <=  8'h00;      memory[13306] <=  8'h00;      memory[13307] <=  8'h00;      memory[13308] <=  8'h00;      memory[13309] <=  8'h00;      memory[13310] <=  8'h00;      memory[13311] <=  8'h00;      memory[13312] <=  8'h00;      memory[13313] <=  8'h00;      memory[13314] <=  8'h00;      memory[13315] <=  8'h00;      memory[13316] <=  8'h00;      memory[13317] <=  8'h00;      memory[13318] <=  8'h00;      memory[13319] <=  8'h00;      memory[13320] <=  8'h00;      memory[13321] <=  8'h00;      memory[13322] <=  8'h00;      memory[13323] <=  8'h00;      memory[13324] <=  8'h00;      memory[13325] <=  8'h00;      memory[13326] <=  8'h00;      memory[13327] <=  8'h00;      memory[13328] <=  8'h00;      memory[13329] <=  8'h00;      memory[13330] <=  8'h00;      memory[13331] <=  8'h00;      memory[13332] <=  8'h00;      memory[13333] <=  8'h00;      memory[13334] <=  8'h00;      memory[13335] <=  8'h00;      memory[13336] <=  8'h00;      memory[13337] <=  8'h00;      memory[13338] <=  8'h00;      memory[13339] <=  8'h00;      memory[13340] <=  8'h00;      memory[13341] <=  8'h00;      memory[13342] <=  8'h00;      memory[13343] <=  8'h00;      memory[13344] <=  8'h00;      memory[13345] <=  8'h00;      memory[13346] <=  8'h00;      memory[13347] <=  8'h00;      memory[13348] <=  8'h00;      memory[13349] <=  8'h00;      memory[13350] <=  8'h00;      memory[13351] <=  8'h00;      memory[13352] <=  8'h00;      memory[13353] <=  8'h00;      memory[13354] <=  8'h00;      memory[13355] <=  8'h00;      memory[13356] <=  8'h00;      memory[13357] <=  8'h00;      memory[13358] <=  8'h00;      memory[13359] <=  8'h00;      memory[13360] <=  8'h00;      memory[13361] <=  8'h00;      memory[13362] <=  8'h00;      memory[13363] <=  8'h00;      memory[13364] <=  8'h00;      memory[13365] <=  8'h00;      memory[13366] <=  8'h00;      memory[13367] <=  8'h00;      memory[13368] <=  8'h00;      memory[13369] <=  8'h00;      memory[13370] <=  8'h00;      memory[13371] <=  8'h00;      memory[13372] <=  8'h00;      memory[13373] <=  8'h00;      memory[13374] <=  8'h00;      memory[13375] <=  8'h00;      memory[13376] <=  8'h00;      memory[13377] <=  8'h00;      memory[13378] <=  8'h00;      memory[13379] <=  8'h00;      memory[13380] <=  8'h00;      memory[13381] <=  8'h00;      memory[13382] <=  8'h00;      memory[13383] <=  8'h00;      memory[13384] <=  8'h00;      memory[13385] <=  8'h00;      memory[13386] <=  8'h00;      memory[13387] <=  8'h00;      memory[13388] <=  8'h00;      memory[13389] <=  8'h00;      memory[13390] <=  8'h00;      memory[13391] <=  8'h00;      memory[13392] <=  8'h00;      memory[13393] <=  8'h00;      memory[13394] <=  8'h00;      memory[13395] <=  8'h00;      memory[13396] <=  8'h00;      memory[13397] <=  8'h00;      memory[13398] <=  8'h00;      memory[13399] <=  8'h00;      memory[13400] <=  8'h00;      memory[13401] <=  8'h00;      memory[13402] <=  8'h00;      memory[13403] <=  8'h00;      memory[13404] <=  8'h00;      memory[13405] <=  8'h00;      memory[13406] <=  8'h00;      memory[13407] <=  8'h00;      memory[13408] <=  8'h00;      memory[13409] <=  8'h00;      memory[13410] <=  8'h00;      memory[13411] <=  8'h00;      memory[13412] <=  8'h00;      memory[13413] <=  8'h00;      memory[13414] <=  8'h00;      memory[13415] <=  8'h00;      memory[13416] <=  8'h00;      memory[13417] <=  8'h00;      memory[13418] <=  8'h00;      memory[13419] <=  8'h00;      memory[13420] <=  8'h00;      memory[13421] <=  8'h00;      memory[13422] <=  8'h00;      memory[13423] <=  8'h00;      memory[13424] <=  8'h00;      memory[13425] <=  8'h00;      memory[13426] <=  8'h00;      memory[13427] <=  8'h00;      memory[13428] <=  8'h00;      memory[13429] <=  8'h00;      memory[13430] <=  8'h00;      memory[13431] <=  8'h00;      memory[13432] <=  8'h00;      memory[13433] <=  8'h00;      memory[13434] <=  8'h00;      memory[13435] <=  8'h00;      memory[13436] <=  8'h00;      memory[13437] <=  8'h00;      memory[13438] <=  8'h00;      memory[13439] <=  8'h00;      memory[13440] <=  8'h00;      memory[13441] <=  8'h00;      memory[13442] <=  8'h00;      memory[13443] <=  8'h00;      memory[13444] <=  8'h00;      memory[13445] <=  8'h00;      memory[13446] <=  8'h00;      memory[13447] <=  8'h00;      memory[13448] <=  8'h00;      memory[13449] <=  8'h00;      memory[13450] <=  8'h00;      memory[13451] <=  8'h00;      memory[13452] <=  8'h00;      memory[13453] <=  8'h00;      memory[13454] <=  8'h00;      memory[13455] <=  8'h00;      memory[13456] <=  8'h00;      memory[13457] <=  8'h00;      memory[13458] <=  8'h00;      memory[13459] <=  8'h00;      memory[13460] <=  8'h00;      memory[13461] <=  8'h00;      memory[13462] <=  8'h00;      memory[13463] <=  8'h00;      memory[13464] <=  8'h00;      memory[13465] <=  8'h00;      memory[13466] <=  8'h00;      memory[13467] <=  8'h00;      memory[13468] <=  8'h00;      memory[13469] <=  8'h00;      memory[13470] <=  8'h00;      memory[13471] <=  8'h00;      memory[13472] <=  8'h00;      memory[13473] <=  8'h00;      memory[13474] <=  8'h00;      memory[13475] <=  8'h00;      memory[13476] <=  8'h00;      memory[13477] <=  8'h00;      memory[13478] <=  8'h00;      memory[13479] <=  8'h00;      memory[13480] <=  8'h00;      memory[13481] <=  8'h00;      memory[13482] <=  8'h00;      memory[13483] <=  8'h00;      memory[13484] <=  8'h00;      memory[13485] <=  8'h00;      memory[13486] <=  8'h00;      memory[13487] <=  8'h00;      memory[13488] <=  8'h00;      memory[13489] <=  8'h00;      memory[13490] <=  8'h00;      memory[13491] <=  8'h00;      memory[13492] <=  8'h00;      memory[13493] <=  8'h00;      memory[13494] <=  8'h00;      memory[13495] <=  8'h00;      memory[13496] <=  8'h00;      memory[13497] <=  8'h00;      memory[13498] <=  8'h00;      memory[13499] <=  8'h00;      memory[13500] <=  8'h00;      memory[13501] <=  8'h00;      memory[13502] <=  8'h00;      memory[13503] <=  8'h00;      memory[13504] <=  8'h00;      memory[13505] <=  8'h00;      memory[13506] <=  8'h00;      memory[13507] <=  8'h00;      memory[13508] <=  8'h00;      memory[13509] <=  8'h00;      memory[13510] <=  8'h00;      memory[13511] <=  8'h00;      memory[13512] <=  8'h00;      memory[13513] <=  8'h00;      memory[13514] <=  8'h00;      memory[13515] <=  8'h00;      memory[13516] <=  8'h00;      memory[13517] <=  8'h00;      memory[13518] <=  8'h00;      memory[13519] <=  8'h00;      memory[13520] <=  8'h00;      memory[13521] <=  8'h00;      memory[13522] <=  8'h00;      memory[13523] <=  8'h00;      memory[13524] <=  8'h00;      memory[13525] <=  8'h00;      memory[13526] <=  8'h00;      memory[13527] <=  8'h00;      memory[13528] <=  8'h00;      memory[13529] <=  8'h00;      memory[13530] <=  8'h00;      memory[13531] <=  8'h00;      memory[13532] <=  8'h00;      memory[13533] <=  8'h00;      memory[13534] <=  8'h00;      memory[13535] <=  8'h00;      memory[13536] <=  8'h00;      memory[13537] <=  8'h00;      memory[13538] <=  8'h00;      memory[13539] <=  8'h00;      memory[13540] <=  8'h00;      memory[13541] <=  8'h00;      memory[13542] <=  8'h00;      memory[13543] <=  8'h00;      memory[13544] <=  8'h00;      memory[13545] <=  8'h00;      memory[13546] <=  8'h00;      memory[13547] <=  8'h00;      memory[13548] <=  8'h00;      memory[13549] <=  8'h00;      memory[13550] <=  8'h00;      memory[13551] <=  8'h00;      memory[13552] <=  8'h00;      memory[13553] <=  8'h00;      memory[13554] <=  8'h00;      memory[13555] <=  8'h00;      memory[13556] <=  8'h00;      memory[13557] <=  8'h00;      memory[13558] <=  8'h00;      memory[13559] <=  8'h00;      memory[13560] <=  8'h00;      memory[13561] <=  8'h00;      memory[13562] <=  8'h00;      memory[13563] <=  8'h00;      memory[13564] <=  8'h00;      memory[13565] <=  8'h00;      memory[13566] <=  8'h00;      memory[13567] <=  8'h00;      memory[13568] <=  8'h00;      memory[13569] <=  8'h00;      memory[13570] <=  8'h00;      memory[13571] <=  8'h00;      memory[13572] <=  8'h00;      memory[13573] <=  8'h00;      memory[13574] <=  8'h00;      memory[13575] <=  8'h00;      memory[13576] <=  8'h00;      memory[13577] <=  8'h00;      memory[13578] <=  8'h00;      memory[13579] <=  8'h00;      memory[13580] <=  8'h00;      memory[13581] <=  8'h00;      memory[13582] <=  8'h00;      memory[13583] <=  8'h00;      memory[13584] <=  8'h00;      memory[13585] <=  8'h00;      memory[13586] <=  8'h00;      memory[13587] <=  8'h00;      memory[13588] <=  8'h00;      memory[13589] <=  8'h00;      memory[13590] <=  8'h00;      memory[13591] <=  8'h00;      memory[13592] <=  8'h00;      memory[13593] <=  8'h00;      memory[13594] <=  8'h00;      memory[13595] <=  8'h00;      memory[13596] <=  8'h00;      memory[13597] <=  8'h00;      memory[13598] <=  8'h00;      memory[13599] <=  8'h00;      memory[13600] <=  8'h00;      memory[13601] <=  8'h00;      memory[13602] <=  8'h00;      memory[13603] <=  8'h00;      memory[13604] <=  8'h00;      memory[13605] <=  8'h00;      memory[13606] <=  8'h00;      memory[13607] <=  8'h00;      memory[13608] <=  8'h00;      memory[13609] <=  8'h00;      memory[13610] <=  8'h00;      memory[13611] <=  8'h00;      memory[13612] <=  8'h00;      memory[13613] <=  8'h00;      memory[13614] <=  8'h00;      memory[13615] <=  8'h00;      memory[13616] <=  8'h00;      memory[13617] <=  8'h00;      memory[13618] <=  8'h00;      memory[13619] <=  8'h00;      memory[13620] <=  8'h00;      memory[13621] <=  8'h00;      memory[13622] <=  8'h00;      memory[13623] <=  8'h00;      memory[13624] <=  8'h00;      memory[13625] <=  8'h00;      memory[13626] <=  8'h00;      memory[13627] <=  8'h00;      memory[13628] <=  8'h00;      memory[13629] <=  8'h00;      memory[13630] <=  8'h00;      memory[13631] <=  8'h00;      memory[13632] <=  8'h00;      memory[13633] <=  8'h00;      memory[13634] <=  8'h00;      memory[13635] <=  8'h00;      memory[13636] <=  8'h00;      memory[13637] <=  8'h00;      memory[13638] <=  8'h00;      memory[13639] <=  8'h00;      memory[13640] <=  8'h00;      memory[13641] <=  8'h00;      memory[13642] <=  8'h00;      memory[13643] <=  8'h00;      memory[13644] <=  8'h00;      memory[13645] <=  8'h00;      memory[13646] <=  8'h00;      memory[13647] <=  8'h00;      memory[13648] <=  8'h00;      memory[13649] <=  8'h00;      memory[13650] <=  8'h00;      memory[13651] <=  8'h00;      memory[13652] <=  8'h00;      memory[13653] <=  8'h00;      memory[13654] <=  8'h00;      memory[13655] <=  8'h00;      memory[13656] <=  8'h00;      memory[13657] <=  8'h00;      memory[13658] <=  8'h00;      memory[13659] <=  8'h00;      memory[13660] <=  8'h00;      memory[13661] <=  8'h00;      memory[13662] <=  8'h00;      memory[13663] <=  8'h00;      memory[13664] <=  8'h00;      memory[13665] <=  8'h00;      memory[13666] <=  8'h00;      memory[13667] <=  8'h00;      memory[13668] <=  8'h00;      memory[13669] <=  8'h00;      memory[13670] <=  8'h00;      memory[13671] <=  8'h00;      memory[13672] <=  8'h00;      memory[13673] <=  8'h00;      memory[13674] <=  8'h00;      memory[13675] <=  8'h00;      memory[13676] <=  8'h00;      memory[13677] <=  8'h00;      memory[13678] <=  8'h00;      memory[13679] <=  8'h00;      memory[13680] <=  8'h00;      memory[13681] <=  8'h00;      memory[13682] <=  8'h00;      memory[13683] <=  8'h00;      memory[13684] <=  8'h00;      memory[13685] <=  8'h00;      memory[13686] <=  8'h00;      memory[13687] <=  8'h00;      memory[13688] <=  8'h00;      memory[13689] <=  8'h00;      memory[13690] <=  8'h00;      memory[13691] <=  8'h00;      memory[13692] <=  8'h00;      memory[13693] <=  8'h00;      memory[13694] <=  8'h00;      memory[13695] <=  8'h00;      memory[13696] <=  8'h00;      memory[13697] <=  8'h00;      memory[13698] <=  8'h00;      memory[13699] <=  8'h00;      memory[13700] <=  8'h00;      memory[13701] <=  8'h00;      memory[13702] <=  8'h00;      memory[13703] <=  8'h00;      memory[13704] <=  8'h00;      memory[13705] <=  8'h00;      memory[13706] <=  8'h00;      memory[13707] <=  8'h00;      memory[13708] <=  8'h00;      memory[13709] <=  8'h00;      memory[13710] <=  8'h00;      memory[13711] <=  8'h00;      memory[13712] <=  8'h00;      memory[13713] <=  8'h00;      memory[13714] <=  8'h00;      memory[13715] <=  8'h00;      memory[13716] <=  8'h00;      memory[13717] <=  8'h00;      memory[13718] <=  8'h00;      memory[13719] <=  8'h00;      memory[13720] <=  8'h00;      memory[13721] <=  8'h00;      memory[13722] <=  8'h00;      memory[13723] <=  8'h00;      memory[13724] <=  8'h00;      memory[13725] <=  8'h00;      memory[13726] <=  8'h00;      memory[13727] <=  8'h00;      memory[13728] <=  8'h00;      memory[13729] <=  8'h00;      memory[13730] <=  8'h00;      memory[13731] <=  8'h00;      memory[13732] <=  8'h00;      memory[13733] <=  8'h00;      memory[13734] <=  8'h00;      memory[13735] <=  8'h00;      memory[13736] <=  8'h00;      memory[13737] <=  8'h00;      memory[13738] <=  8'h00;      memory[13739] <=  8'h00;      memory[13740] <=  8'h00;      memory[13741] <=  8'h00;      memory[13742] <=  8'h00;      memory[13743] <=  8'h00;      memory[13744] <=  8'h00;      memory[13745] <=  8'h00;      memory[13746] <=  8'h00;      memory[13747] <=  8'h00;      memory[13748] <=  8'h00;      memory[13749] <=  8'h00;      memory[13750] <=  8'h00;      memory[13751] <=  8'h00;      memory[13752] <=  8'h00;      memory[13753] <=  8'h00;      memory[13754] <=  8'h00;      memory[13755] <=  8'h00;      memory[13756] <=  8'h00;      memory[13757] <=  8'h00;      memory[13758] <=  8'h00;      memory[13759] <=  8'h00;      memory[13760] <=  8'h00;      memory[13761] <=  8'h00;      memory[13762] <=  8'h00;      memory[13763] <=  8'h00;      memory[13764] <=  8'h00;      memory[13765] <=  8'h00;      memory[13766] <=  8'h00;      memory[13767] <=  8'h00;      memory[13768] <=  8'h00;      memory[13769] <=  8'h00;      memory[13770] <=  8'h00;      memory[13771] <=  8'h00;      memory[13772] <=  8'h00;      memory[13773] <=  8'h00;      memory[13774] <=  8'h00;      memory[13775] <=  8'h00;      memory[13776] <=  8'h00;      memory[13777] <=  8'h00;      memory[13778] <=  8'h00;      memory[13779] <=  8'h00;      memory[13780] <=  8'h00;      memory[13781] <=  8'h00;      memory[13782] <=  8'h00;      memory[13783] <=  8'h00;      memory[13784] <=  8'h00;      memory[13785] <=  8'h00;      memory[13786] <=  8'h00;      memory[13787] <=  8'h00;      memory[13788] <=  8'h00;      memory[13789] <=  8'h00;      memory[13790] <=  8'h00;      memory[13791] <=  8'h00;      memory[13792] <=  8'h00;      memory[13793] <=  8'h00;      memory[13794] <=  8'h00;      memory[13795] <=  8'h00;      memory[13796] <=  8'h00;      memory[13797] <=  8'h00;      memory[13798] <=  8'h00;      memory[13799] <=  8'h00;      memory[13800] <=  8'h00;      memory[13801] <=  8'h00;      memory[13802] <=  8'h00;      memory[13803] <=  8'h00;      memory[13804] <=  8'h00;      memory[13805] <=  8'h00;      memory[13806] <=  8'h00;      memory[13807] <=  8'h00;      memory[13808] <=  8'h00;      memory[13809] <=  8'h00;      memory[13810] <=  8'h00;      memory[13811] <=  8'h00;      memory[13812] <=  8'h00;      memory[13813] <=  8'h00;      memory[13814] <=  8'h00;      memory[13815] <=  8'h00;      memory[13816] <=  8'h00;      memory[13817] <=  8'h00;      memory[13818] <=  8'h00;      memory[13819] <=  8'h00;      memory[13820] <=  8'h00;      memory[13821] <=  8'h00;      memory[13822] <=  8'h00;      memory[13823] <=  8'h00;      memory[13824] <=  8'h00;      memory[13825] <=  8'h00;      memory[13826] <=  8'h00;      memory[13827] <=  8'h00;      memory[13828] <=  8'h00;      memory[13829] <=  8'h00;      memory[13830] <=  8'h00;      memory[13831] <=  8'h00;      memory[13832] <=  8'h00;      memory[13833] <=  8'h00;      memory[13834] <=  8'h00;      memory[13835] <=  8'h00;      memory[13836] <=  8'h00;      memory[13837] <=  8'h00;      memory[13838] <=  8'h00;      memory[13839] <=  8'h00;      memory[13840] <=  8'h00;      memory[13841] <=  8'h00;      memory[13842] <=  8'h00;      memory[13843] <=  8'h00;      memory[13844] <=  8'h00;      memory[13845] <=  8'h00;      memory[13846] <=  8'h00;      memory[13847] <=  8'h00;      memory[13848] <=  8'h00;      memory[13849] <=  8'h00;      memory[13850] <=  8'h00;      memory[13851] <=  8'h00;      memory[13852] <=  8'h00;      memory[13853] <=  8'h00;      memory[13854] <=  8'h00;      memory[13855] <=  8'h00;      memory[13856] <=  8'h00;      memory[13857] <=  8'h00;      memory[13858] <=  8'h00;      memory[13859] <=  8'h00;      memory[13860] <=  8'h00;      memory[13861] <=  8'h00;      memory[13862] <=  8'h00;      memory[13863] <=  8'h00;      memory[13864] <=  8'h00;      memory[13865] <=  8'h00;      memory[13866] <=  8'h00;      memory[13867] <=  8'h00;      memory[13868] <=  8'h00;      memory[13869] <=  8'h00;      memory[13870] <=  8'h00;      memory[13871] <=  8'h00;      memory[13872] <=  8'h00;      memory[13873] <=  8'h00;      memory[13874] <=  8'h00;      memory[13875] <=  8'h00;      memory[13876] <=  8'h00;      memory[13877] <=  8'h00;      memory[13878] <=  8'h00;      memory[13879] <=  8'h00;      memory[13880] <=  8'h00;      memory[13881] <=  8'h00;      memory[13882] <=  8'h00;      memory[13883] <=  8'h00;      memory[13884] <=  8'h00;      memory[13885] <=  8'h00;      memory[13886] <=  8'h00;      memory[13887] <=  8'h00;      memory[13888] <=  8'h00;      memory[13889] <=  8'h00;      memory[13890] <=  8'h00;      memory[13891] <=  8'h00;      memory[13892] <=  8'h00;      memory[13893] <=  8'h00;      memory[13894] <=  8'h00;      memory[13895] <=  8'h00;      memory[13896] <=  8'h00;      memory[13897] <=  8'h00;      memory[13898] <=  8'h00;      memory[13899] <=  8'h00;      memory[13900] <=  8'h00;      memory[13901] <=  8'h00;      memory[13902] <=  8'h00;      memory[13903] <=  8'h00;      memory[13904] <=  8'h00;      memory[13905] <=  8'h00;      memory[13906] <=  8'h00;      memory[13907] <=  8'h00;      memory[13908] <=  8'h00;      memory[13909] <=  8'h00;      memory[13910] <=  8'h00;      memory[13911] <=  8'h00;      memory[13912] <=  8'h00;      memory[13913] <=  8'h00;      memory[13914] <=  8'h00;      memory[13915] <=  8'h00;      memory[13916] <=  8'h00;      memory[13917] <=  8'h00;      memory[13918] <=  8'h00;      memory[13919] <=  8'h00;      memory[13920] <=  8'h00;      memory[13921] <=  8'h00;      memory[13922] <=  8'h00;      memory[13923] <=  8'h00;      memory[13924] <=  8'h00;      memory[13925] <=  8'h00;      memory[13926] <=  8'h00;      memory[13927] <=  8'h00;      memory[13928] <=  8'h00;      memory[13929] <=  8'h00;      memory[13930] <=  8'h00;      memory[13931] <=  8'h00;      memory[13932] <=  8'h00;      memory[13933] <=  8'h00;      memory[13934] <=  8'h00;      memory[13935] <=  8'h00;      memory[13936] <=  8'h00;      memory[13937] <=  8'h00;      memory[13938] <=  8'h00;      memory[13939] <=  8'h00;      memory[13940] <=  8'h00;      memory[13941] <=  8'h00;      memory[13942] <=  8'h00;      memory[13943] <=  8'h00;      memory[13944] <=  8'h00;      memory[13945] <=  8'h00;      memory[13946] <=  8'h00;      memory[13947] <=  8'h00;      memory[13948] <=  8'h00;      memory[13949] <=  8'h00;      memory[13950] <=  8'h00;      memory[13951] <=  8'h00;      memory[13952] <=  8'h00;      memory[13953] <=  8'h00;      memory[13954] <=  8'h00;      memory[13955] <=  8'h00;      memory[13956] <=  8'h00;      memory[13957] <=  8'h00;      memory[13958] <=  8'h00;      memory[13959] <=  8'h00;      memory[13960] <=  8'h00;      memory[13961] <=  8'h00;      memory[13962] <=  8'h00;      memory[13963] <=  8'h00;      memory[13964] <=  8'h00;      memory[13965] <=  8'h00;      memory[13966] <=  8'h00;      memory[13967] <=  8'h00;      memory[13968] <=  8'h00;      memory[13969] <=  8'h00;      memory[13970] <=  8'h00;      memory[13971] <=  8'h00;      memory[13972] <=  8'h00;      memory[13973] <=  8'h00;      memory[13974] <=  8'h00;      memory[13975] <=  8'h00;      memory[13976] <=  8'h00;      memory[13977] <=  8'h00;      memory[13978] <=  8'h00;      memory[13979] <=  8'h00;      memory[13980] <=  8'h00;      memory[13981] <=  8'h00;      memory[13982] <=  8'h00;      memory[13983] <=  8'h00;      memory[13984] <=  8'h00;      memory[13985] <=  8'h00;      memory[13986] <=  8'h00;      memory[13987] <=  8'h00;      memory[13988] <=  8'h00;      memory[13989] <=  8'h00;      memory[13990] <=  8'h00;      memory[13991] <=  8'h00;      memory[13992] <=  8'h00;      memory[13993] <=  8'h00;      memory[13994] <=  8'h00;      memory[13995] <=  8'h00;      memory[13996] <=  8'h00;      memory[13997] <=  8'h00;      memory[13998] <=  8'h00;      memory[13999] <=  8'h00;      memory[14000] <=  8'h00;      memory[14001] <=  8'h00;      memory[14002] <=  8'h00;      memory[14003] <=  8'h00;      memory[14004] <=  8'h00;      memory[14005] <=  8'h00;      memory[14006] <=  8'h00;      memory[14007] <=  8'h00;      memory[14008] <=  8'h00;      memory[14009] <=  8'h00;      memory[14010] <=  8'h00;      memory[14011] <=  8'h00;      memory[14012] <=  8'h00;      memory[14013] <=  8'h00;      memory[14014] <=  8'h00;      memory[14015] <=  8'h00;      memory[14016] <=  8'h00;      memory[14017] <=  8'h00;      memory[14018] <=  8'h00;      memory[14019] <=  8'h00;      memory[14020] <=  8'h00;      memory[14021] <=  8'h00;      memory[14022] <=  8'h00;      memory[14023] <=  8'h00;      memory[14024] <=  8'h00;      memory[14025] <=  8'h00;      memory[14026] <=  8'h00;      memory[14027] <=  8'h00;      memory[14028] <=  8'h00;      memory[14029] <=  8'h00;      memory[14030] <=  8'h00;      memory[14031] <=  8'h00;      memory[14032] <=  8'h00;      memory[14033] <=  8'h00;      memory[14034] <=  8'h00;      memory[14035] <=  8'h00;      memory[14036] <=  8'h00;      memory[14037] <=  8'h00;      memory[14038] <=  8'h00;      memory[14039] <=  8'h00;      memory[14040] <=  8'h00;      memory[14041] <=  8'h00;      memory[14042] <=  8'h00;      memory[14043] <=  8'h00;      memory[14044] <=  8'h00;      memory[14045] <=  8'h00;      memory[14046] <=  8'h00;      memory[14047] <=  8'h00;      memory[14048] <=  8'h00;      memory[14049] <=  8'h00;      memory[14050] <=  8'h00;      memory[14051] <=  8'h00;      memory[14052] <=  8'h00;      memory[14053] <=  8'h00;      memory[14054] <=  8'h00;      memory[14055] <=  8'h00;      memory[14056] <=  8'h00;      memory[14057] <=  8'h00;      memory[14058] <=  8'h00;      memory[14059] <=  8'h00;      memory[14060] <=  8'h00;      memory[14061] <=  8'h00;      memory[14062] <=  8'h00;      memory[14063] <=  8'h00;      memory[14064] <=  8'h00;      memory[14065] <=  8'h00;      memory[14066] <=  8'h00;      memory[14067] <=  8'h00;      memory[14068] <=  8'h00;      memory[14069] <=  8'h00;      memory[14070] <=  8'h00;      memory[14071] <=  8'h00;      memory[14072] <=  8'h00;      memory[14073] <=  8'h00;      memory[14074] <=  8'h00;      memory[14075] <=  8'h00;      memory[14076] <=  8'h00;      memory[14077] <=  8'h00;      memory[14078] <=  8'h00;      memory[14079] <=  8'h00;      memory[14080] <=  8'h00;      memory[14081] <=  8'h00;      memory[14082] <=  8'h00;      memory[14083] <=  8'h00;      memory[14084] <=  8'h00;      memory[14085] <=  8'h00;      memory[14086] <=  8'h00;      memory[14087] <=  8'h00;      memory[14088] <=  8'h00;      memory[14089] <=  8'h00;      memory[14090] <=  8'h00;      memory[14091] <=  8'h00;      memory[14092] <=  8'h00;      memory[14093] <=  8'h00;      memory[14094] <=  8'h00;      memory[14095] <=  8'h00;      memory[14096] <=  8'h00;      memory[14097] <=  8'h00;      memory[14098] <=  8'h00;      memory[14099] <=  8'h00;      memory[14100] <=  8'h00;      memory[14101] <=  8'h00;      memory[14102] <=  8'h00;      memory[14103] <=  8'h00;      memory[14104] <=  8'h00;      memory[14105] <=  8'h00;      memory[14106] <=  8'h00;      memory[14107] <=  8'h00;      memory[14108] <=  8'h00;      memory[14109] <=  8'h00;      memory[14110] <=  8'h00;      memory[14111] <=  8'h00;      memory[14112] <=  8'h00;      memory[14113] <=  8'h00;      memory[14114] <=  8'h00;      memory[14115] <=  8'h00;      memory[14116] <=  8'h00;      memory[14117] <=  8'h00;      memory[14118] <=  8'h00;      memory[14119] <=  8'h00;      memory[14120] <=  8'h00;      memory[14121] <=  8'h00;      memory[14122] <=  8'h00;      memory[14123] <=  8'h00;      memory[14124] <=  8'h00;      memory[14125] <=  8'h00;      memory[14126] <=  8'h00;      memory[14127] <=  8'h00;      memory[14128] <=  8'h00;      memory[14129] <=  8'h00;      memory[14130] <=  8'h00;      memory[14131] <=  8'h00;      memory[14132] <=  8'h00;      memory[14133] <=  8'h00;      memory[14134] <=  8'h00;      memory[14135] <=  8'h00;      memory[14136] <=  8'h00;      memory[14137] <=  8'h00;      memory[14138] <=  8'h00;      memory[14139] <=  8'h00;      memory[14140] <=  8'h00;      memory[14141] <=  8'h00;      memory[14142] <=  8'h00;      memory[14143] <=  8'h00;      memory[14144] <=  8'h00;      memory[14145] <=  8'h00;      memory[14146] <=  8'h00;      memory[14147] <=  8'h00;      memory[14148] <=  8'h00;      memory[14149] <=  8'h00;      memory[14150] <=  8'h00;      memory[14151] <=  8'h00;      memory[14152] <=  8'h00;      memory[14153] <=  8'h00;      memory[14154] <=  8'h00;      memory[14155] <=  8'h00;      memory[14156] <=  8'h00;      memory[14157] <=  8'h00;      memory[14158] <=  8'h00;      memory[14159] <=  8'h00;      memory[14160] <=  8'h00;      memory[14161] <=  8'h00;      memory[14162] <=  8'h00;      memory[14163] <=  8'h00;      memory[14164] <=  8'h00;      memory[14165] <=  8'h00;      memory[14166] <=  8'h00;      memory[14167] <=  8'h00;      memory[14168] <=  8'h00;      memory[14169] <=  8'h00;      memory[14170] <=  8'h00;      memory[14171] <=  8'h00;      memory[14172] <=  8'h00;      memory[14173] <=  8'h00;      memory[14174] <=  8'h00;      memory[14175] <=  8'h00;      memory[14176] <=  8'h00;      memory[14177] <=  8'h00;      memory[14178] <=  8'h00;      memory[14179] <=  8'h00;      memory[14180] <=  8'h00;      memory[14181] <=  8'h00;      memory[14182] <=  8'h00;      memory[14183] <=  8'h00;      memory[14184] <=  8'h00;      memory[14185] <=  8'h00;      memory[14186] <=  8'h00;      memory[14187] <=  8'h00;      memory[14188] <=  8'h00;      memory[14189] <=  8'h00;      memory[14190] <=  8'h00;      memory[14191] <=  8'h00;      memory[14192] <=  8'h00;      memory[14193] <=  8'h00;      memory[14194] <=  8'h00;      memory[14195] <=  8'h00;      memory[14196] <=  8'h00;      memory[14197] <=  8'h00;      memory[14198] <=  8'h00;      memory[14199] <=  8'h00;      memory[14200] <=  8'h00;      memory[14201] <=  8'h00;      memory[14202] <=  8'h00;      memory[14203] <=  8'h00;      memory[14204] <=  8'h00;      memory[14205] <=  8'h00;      memory[14206] <=  8'h00;      memory[14207] <=  8'h00;      memory[14208] <=  8'h00;      memory[14209] <=  8'h00;      memory[14210] <=  8'h00;      memory[14211] <=  8'h00;      memory[14212] <=  8'h00;      memory[14213] <=  8'h00;      memory[14214] <=  8'h00;      memory[14215] <=  8'h00;      memory[14216] <=  8'h00;      memory[14217] <=  8'h00;      memory[14218] <=  8'h00;      memory[14219] <=  8'h00;      memory[14220] <=  8'h00;      memory[14221] <=  8'h00;      memory[14222] <=  8'h00;      memory[14223] <=  8'h00;      memory[14224] <=  8'h00;      memory[14225] <=  8'h00;      memory[14226] <=  8'h00;      memory[14227] <=  8'h00;      memory[14228] <=  8'h00;      memory[14229] <=  8'h00;      memory[14230] <=  8'h00;      memory[14231] <=  8'h00;      memory[14232] <=  8'h00;      memory[14233] <=  8'h00;      memory[14234] <=  8'h00;      memory[14235] <=  8'h00;      memory[14236] <=  8'h00;      memory[14237] <=  8'h00;      memory[14238] <=  8'h00;      memory[14239] <=  8'h00;      memory[14240] <=  8'h00;      memory[14241] <=  8'h00;      memory[14242] <=  8'h00;      memory[14243] <=  8'h00;      memory[14244] <=  8'h00;      memory[14245] <=  8'h00;      memory[14246] <=  8'h00;      memory[14247] <=  8'h00;      memory[14248] <=  8'h00;      memory[14249] <=  8'h00;      memory[14250] <=  8'h00;      memory[14251] <=  8'h00;      memory[14252] <=  8'h00;      memory[14253] <=  8'h00;      memory[14254] <=  8'h00;      memory[14255] <=  8'h00;      memory[14256] <=  8'h00;      memory[14257] <=  8'h00;      memory[14258] <=  8'h00;      memory[14259] <=  8'h00;      memory[14260] <=  8'h00;      memory[14261] <=  8'h00;      memory[14262] <=  8'h00;      memory[14263] <=  8'h00;      memory[14264] <=  8'h00;      memory[14265] <=  8'h00;      memory[14266] <=  8'h00;      memory[14267] <=  8'h00;      memory[14268] <=  8'h00;      memory[14269] <=  8'h00;      memory[14270] <=  8'h00;      memory[14271] <=  8'h00;      memory[14272] <=  8'h00;      memory[14273] <=  8'h00;      memory[14274] <=  8'h00;      memory[14275] <=  8'h00;      memory[14276] <=  8'h00;      memory[14277] <=  8'h00;      memory[14278] <=  8'h00;      memory[14279] <=  8'h00;      memory[14280] <=  8'h00;      memory[14281] <=  8'h00;      memory[14282] <=  8'h00;      memory[14283] <=  8'h00;      memory[14284] <=  8'h00;      memory[14285] <=  8'h00;      memory[14286] <=  8'h00;      memory[14287] <=  8'h00;      memory[14288] <=  8'h00;      memory[14289] <=  8'h00;      memory[14290] <=  8'h00;      memory[14291] <=  8'h00;      memory[14292] <=  8'h00;      memory[14293] <=  8'h00;      memory[14294] <=  8'h00;      memory[14295] <=  8'h00;      memory[14296] <=  8'h00;      memory[14297] <=  8'h00;      memory[14298] <=  8'h00;      memory[14299] <=  8'h00;      memory[14300] <=  8'h00;      memory[14301] <=  8'h00;      memory[14302] <=  8'h00;      memory[14303] <=  8'h00;      memory[14304] <=  8'h00;      memory[14305] <=  8'h00;      memory[14306] <=  8'h00;      memory[14307] <=  8'h00;      memory[14308] <=  8'h00;      memory[14309] <=  8'h00;      memory[14310] <=  8'h00;      memory[14311] <=  8'h00;      memory[14312] <=  8'h00;      memory[14313] <=  8'h00;      memory[14314] <=  8'h00;      memory[14315] <=  8'h00;      memory[14316] <=  8'h00;      memory[14317] <=  8'h00;      memory[14318] <=  8'h00;      memory[14319] <=  8'h00;      memory[14320] <=  8'h00;      memory[14321] <=  8'h00;      memory[14322] <=  8'h00;      memory[14323] <=  8'h00;      memory[14324] <=  8'h00;      memory[14325] <=  8'h00;      memory[14326] <=  8'h00;      memory[14327] <=  8'h00;      memory[14328] <=  8'h00;      memory[14329] <=  8'h00;      memory[14330] <=  8'h00;      memory[14331] <=  8'h00;      memory[14332] <=  8'h00;      memory[14333] <=  8'h00;      memory[14334] <=  8'h00;      memory[14335] <=  8'h00;      memory[14336] <=  8'h00;      memory[14337] <=  8'h00;      memory[14338] <=  8'h00;      memory[14339] <=  8'h00;      memory[14340] <=  8'h00;      memory[14341] <=  8'h00;      memory[14342] <=  8'h00;      memory[14343] <=  8'h00;      memory[14344] <=  8'h00;      memory[14345] <=  8'h00;      memory[14346] <=  8'h00;      memory[14347] <=  8'h00;      memory[14348] <=  8'h00;      memory[14349] <=  8'h00;      memory[14350] <=  8'h00;      memory[14351] <=  8'h00;      memory[14352] <=  8'h00;      memory[14353] <=  8'h00;      memory[14354] <=  8'h00;      memory[14355] <=  8'h00;      memory[14356] <=  8'h00;      memory[14357] <=  8'h00;      memory[14358] <=  8'h00;      memory[14359] <=  8'h00;      memory[14360] <=  8'h00;      memory[14361] <=  8'h00;      memory[14362] <=  8'h00;      memory[14363] <=  8'h00;      memory[14364] <=  8'h00;      memory[14365] <=  8'h00;      memory[14366] <=  8'h00;      memory[14367] <=  8'h00;      memory[14368] <=  8'h00;      memory[14369] <=  8'h00;      memory[14370] <=  8'h00;      memory[14371] <=  8'h00;      memory[14372] <=  8'h00;      memory[14373] <=  8'h00;      memory[14374] <=  8'h00;      memory[14375] <=  8'h00;      memory[14376] <=  8'h00;      memory[14377] <=  8'h00;      memory[14378] <=  8'h00;      memory[14379] <=  8'h00;      memory[14380] <=  8'h00;      memory[14381] <=  8'h00;      memory[14382] <=  8'h00;      memory[14383] <=  8'h00;      memory[14384] <=  8'h00;      memory[14385] <=  8'h00;      memory[14386] <=  8'h00;      memory[14387] <=  8'h00;      memory[14388] <=  8'h00;      memory[14389] <=  8'h00;      memory[14390] <=  8'h00;      memory[14391] <=  8'h00;      memory[14392] <=  8'h00;      memory[14393] <=  8'h00;      memory[14394] <=  8'h00;      memory[14395] <=  8'h00;      memory[14396] <=  8'h00;      memory[14397] <=  8'h00;      memory[14398] <=  8'h00;      memory[14399] <=  8'h00;      memory[14400] <=  8'h00;      memory[14401] <=  8'h00;      memory[14402] <=  8'h00;      memory[14403] <=  8'h00;      memory[14404] <=  8'h00;      memory[14405] <=  8'h00;      memory[14406] <=  8'h00;      memory[14407] <=  8'h00;      memory[14408] <=  8'h00;      memory[14409] <=  8'h00;      memory[14410] <=  8'h00;      memory[14411] <=  8'h00;      memory[14412] <=  8'h00;      memory[14413] <=  8'h00;      memory[14414] <=  8'h00;      memory[14415] <=  8'h00;      memory[14416] <=  8'h00;      memory[14417] <=  8'h00;      memory[14418] <=  8'h00;      memory[14419] <=  8'h00;      memory[14420] <=  8'h00;      memory[14421] <=  8'h00;      memory[14422] <=  8'h00;      memory[14423] <=  8'h00;      memory[14424] <=  8'h00;      memory[14425] <=  8'h00;      memory[14426] <=  8'h00;      memory[14427] <=  8'h00;      memory[14428] <=  8'h00;      memory[14429] <=  8'h00;      memory[14430] <=  8'h00;      memory[14431] <=  8'h00;      memory[14432] <=  8'h00;      memory[14433] <=  8'h00;      memory[14434] <=  8'h00;      memory[14435] <=  8'h00;      memory[14436] <=  8'h00;      memory[14437] <=  8'h00;      memory[14438] <=  8'h00;      memory[14439] <=  8'h00;      memory[14440] <=  8'h00;      memory[14441] <=  8'h00;      memory[14442] <=  8'h00;      memory[14443] <=  8'h00;      memory[14444] <=  8'h00;      memory[14445] <=  8'h00;      memory[14446] <=  8'h00;      memory[14447] <=  8'h00;      memory[14448] <=  8'h00;      memory[14449] <=  8'h00;      memory[14450] <=  8'h00;      memory[14451] <=  8'h00;      memory[14452] <=  8'h00;      memory[14453] <=  8'h00;      memory[14454] <=  8'h00;      memory[14455] <=  8'h00;      memory[14456] <=  8'h00;      memory[14457] <=  8'h00;      memory[14458] <=  8'h00;      memory[14459] <=  8'h00;      memory[14460] <=  8'h00;      memory[14461] <=  8'h00;      memory[14462] <=  8'h00;      memory[14463] <=  8'h00;      memory[14464] <=  8'h00;      memory[14465] <=  8'h00;      memory[14466] <=  8'h00;      memory[14467] <=  8'h00;      memory[14468] <=  8'h00;      memory[14469] <=  8'h00;      memory[14470] <=  8'h00;      memory[14471] <=  8'h00;      memory[14472] <=  8'h00;      memory[14473] <=  8'h00;      memory[14474] <=  8'h00;      memory[14475] <=  8'h00;      memory[14476] <=  8'h00;      memory[14477] <=  8'h00;      memory[14478] <=  8'h00;      memory[14479] <=  8'h00;      memory[14480] <=  8'h00;      memory[14481] <=  8'h00;      memory[14482] <=  8'h00;      memory[14483] <=  8'h00;      memory[14484] <=  8'h00;      memory[14485] <=  8'h00;      memory[14486] <=  8'h00;      memory[14487] <=  8'h00;      memory[14488] <=  8'h00;      memory[14489] <=  8'h00;      memory[14490] <=  8'h00;      memory[14491] <=  8'h00;      memory[14492] <=  8'h00;      memory[14493] <=  8'h00;      memory[14494] <=  8'h00;      memory[14495] <=  8'h00;      memory[14496] <=  8'h00;      memory[14497] <=  8'h00;      memory[14498] <=  8'h00;      memory[14499] <=  8'h00;      memory[14500] <=  8'h00;      memory[14501] <=  8'h00;      memory[14502] <=  8'h00;      memory[14503] <=  8'h00;      memory[14504] <=  8'h00;      memory[14505] <=  8'h00;      memory[14506] <=  8'h00;      memory[14507] <=  8'h00;      memory[14508] <=  8'h00;      memory[14509] <=  8'h00;      memory[14510] <=  8'h00;      memory[14511] <=  8'h00;      memory[14512] <=  8'h00;      memory[14513] <=  8'h00;      memory[14514] <=  8'h00;      memory[14515] <=  8'h00;      memory[14516] <=  8'h00;      memory[14517] <=  8'h00;      memory[14518] <=  8'h00;      memory[14519] <=  8'h00;      memory[14520] <=  8'h00;      memory[14521] <=  8'h00;      memory[14522] <=  8'h00;      memory[14523] <=  8'h00;      memory[14524] <=  8'h00;      memory[14525] <=  8'h00;      memory[14526] <=  8'h00;      memory[14527] <=  8'h00;      memory[14528] <=  8'h00;      memory[14529] <=  8'h00;      memory[14530] <=  8'h00;      memory[14531] <=  8'h00;      memory[14532] <=  8'h00;      memory[14533] <=  8'h00;      memory[14534] <=  8'h00;      memory[14535] <=  8'h00;      memory[14536] <=  8'h00;      memory[14537] <=  8'h00;      memory[14538] <=  8'h00;      memory[14539] <=  8'h00;      memory[14540] <=  8'h00;      memory[14541] <=  8'h00;      memory[14542] <=  8'h00;      memory[14543] <=  8'h00;      memory[14544] <=  8'h00;      memory[14545] <=  8'h00;      memory[14546] <=  8'h00;      memory[14547] <=  8'h00;      memory[14548] <=  8'h00;      memory[14549] <=  8'h00;      memory[14550] <=  8'h00;      memory[14551] <=  8'h00;      memory[14552] <=  8'h00;      memory[14553] <=  8'h00;      memory[14554] <=  8'h00;      memory[14555] <=  8'h00;      memory[14556] <=  8'h00;      memory[14557] <=  8'h00;      memory[14558] <=  8'h00;      memory[14559] <=  8'h00;      memory[14560] <=  8'h00;      memory[14561] <=  8'h00;      memory[14562] <=  8'h00;      memory[14563] <=  8'h00;      memory[14564] <=  8'h00;      memory[14565] <=  8'h00;      memory[14566] <=  8'h00;      memory[14567] <=  8'h00;      memory[14568] <=  8'h00;      memory[14569] <=  8'h00;      memory[14570] <=  8'h00;      memory[14571] <=  8'h00;      memory[14572] <=  8'h00;      memory[14573] <=  8'h00;      memory[14574] <=  8'h00;      memory[14575] <=  8'h00;      memory[14576] <=  8'h00;      memory[14577] <=  8'h00;      memory[14578] <=  8'h00;      memory[14579] <=  8'h00;      memory[14580] <=  8'h00;      memory[14581] <=  8'h00;      memory[14582] <=  8'h00;      memory[14583] <=  8'h00;      memory[14584] <=  8'h00;      memory[14585] <=  8'h00;      memory[14586] <=  8'h00;      memory[14587] <=  8'h00;      memory[14588] <=  8'h00;      memory[14589] <=  8'h00;      memory[14590] <=  8'h00;      memory[14591] <=  8'h00;      memory[14592] <=  8'h00;      memory[14593] <=  8'h00;      memory[14594] <=  8'h00;      memory[14595] <=  8'h00;      memory[14596] <=  8'h00;      memory[14597] <=  8'h00;      memory[14598] <=  8'h00;      memory[14599] <=  8'h00;      memory[14600] <=  8'h00;      memory[14601] <=  8'h00;      memory[14602] <=  8'h00;      memory[14603] <=  8'h00;      memory[14604] <=  8'h00;      memory[14605] <=  8'h00;      memory[14606] <=  8'h00;      memory[14607] <=  8'h00;      memory[14608] <=  8'h00;      memory[14609] <=  8'h00;      memory[14610] <=  8'h00;      memory[14611] <=  8'h00;      memory[14612] <=  8'h00;      memory[14613] <=  8'h00;      memory[14614] <=  8'h00;      memory[14615] <=  8'h00;      memory[14616] <=  8'h00;      memory[14617] <=  8'h00;      memory[14618] <=  8'h00;      memory[14619] <=  8'h00;      memory[14620] <=  8'h00;      memory[14621] <=  8'h00;      memory[14622] <=  8'h00;      memory[14623] <=  8'h00;      memory[14624] <=  8'h00;      memory[14625] <=  8'h00;      memory[14626] <=  8'h00;      memory[14627] <=  8'h00;      memory[14628] <=  8'h00;      memory[14629] <=  8'h00;      memory[14630] <=  8'h00;      memory[14631] <=  8'h00;      memory[14632] <=  8'h00;      memory[14633] <=  8'h00;      memory[14634] <=  8'h00;      memory[14635] <=  8'h00;      memory[14636] <=  8'h00;      memory[14637] <=  8'h00;      memory[14638] <=  8'h00;      memory[14639] <=  8'h00;      memory[14640] <=  8'h00;      memory[14641] <=  8'h00;      memory[14642] <=  8'h00;      memory[14643] <=  8'h00;      memory[14644] <=  8'h00;      memory[14645] <=  8'h00;      memory[14646] <=  8'h00;      memory[14647] <=  8'h00;      memory[14648] <=  8'h00;      memory[14649] <=  8'h00;      memory[14650] <=  8'h00;      memory[14651] <=  8'h00;      memory[14652] <=  8'h00;      memory[14653] <=  8'h00;      memory[14654] <=  8'h00;      memory[14655] <=  8'h00;      memory[14656] <=  8'h00;      memory[14657] <=  8'h00;      memory[14658] <=  8'h00;      memory[14659] <=  8'h00;      memory[14660] <=  8'h00;      memory[14661] <=  8'h00;      memory[14662] <=  8'h00;      memory[14663] <=  8'h00;      memory[14664] <=  8'h00;      memory[14665] <=  8'h00;      memory[14666] <=  8'h00;      memory[14667] <=  8'h00;      memory[14668] <=  8'h00;      memory[14669] <=  8'h00;      memory[14670] <=  8'h00;      memory[14671] <=  8'h00;      memory[14672] <=  8'h00;      memory[14673] <=  8'h00;      memory[14674] <=  8'h00;      memory[14675] <=  8'h00;      memory[14676] <=  8'h00;      memory[14677] <=  8'h00;      memory[14678] <=  8'h00;      memory[14679] <=  8'h00;      memory[14680] <=  8'h00;      memory[14681] <=  8'h00;      memory[14682] <=  8'h00;      memory[14683] <=  8'h00;      memory[14684] <=  8'h00;      memory[14685] <=  8'h00;      memory[14686] <=  8'h00;      memory[14687] <=  8'h00;      memory[14688] <=  8'h00;      memory[14689] <=  8'h00;      memory[14690] <=  8'h00;      memory[14691] <=  8'h00;      memory[14692] <=  8'h00;      memory[14693] <=  8'h00;      memory[14694] <=  8'h00;      memory[14695] <=  8'h00;      memory[14696] <=  8'h00;      memory[14697] <=  8'h00;      memory[14698] <=  8'h00;      memory[14699] <=  8'h00;      memory[14700] <=  8'h00;      memory[14701] <=  8'h00;      memory[14702] <=  8'h00;      memory[14703] <=  8'h00;      memory[14704] <=  8'h00;      memory[14705] <=  8'h00;      memory[14706] <=  8'h00;      memory[14707] <=  8'h00;      memory[14708] <=  8'h00;      memory[14709] <=  8'h00;      memory[14710] <=  8'h00;      memory[14711] <=  8'h00;      memory[14712] <=  8'h00;      memory[14713] <=  8'h00;      memory[14714] <=  8'h00;      memory[14715] <=  8'h00;      memory[14716] <=  8'h00;      memory[14717] <=  8'h00;      memory[14718] <=  8'h00;      memory[14719] <=  8'h00;      memory[14720] <=  8'h00;      memory[14721] <=  8'h00;      memory[14722] <=  8'h00;      memory[14723] <=  8'h00;      memory[14724] <=  8'h00;      memory[14725] <=  8'h00;      memory[14726] <=  8'h00;      memory[14727] <=  8'h00;      memory[14728] <=  8'h00;      memory[14729] <=  8'h00;      memory[14730] <=  8'h00;      memory[14731] <=  8'h00;      memory[14732] <=  8'h00;      memory[14733] <=  8'h00;      memory[14734] <=  8'h00;      memory[14735] <=  8'h00;      memory[14736] <=  8'h00;      memory[14737] <=  8'h00;      memory[14738] <=  8'h00;      memory[14739] <=  8'h00;      memory[14740] <=  8'h00;      memory[14741] <=  8'h00;      memory[14742] <=  8'h00;      memory[14743] <=  8'h00;      memory[14744] <=  8'h00;      memory[14745] <=  8'h00;      memory[14746] <=  8'h00;      memory[14747] <=  8'h00;      memory[14748] <=  8'h00;      memory[14749] <=  8'h00;      memory[14750] <=  8'h00;      memory[14751] <=  8'h00;      memory[14752] <=  8'h00;      memory[14753] <=  8'h00;      memory[14754] <=  8'h00;      memory[14755] <=  8'h00;      memory[14756] <=  8'h00;      memory[14757] <=  8'h00;      memory[14758] <=  8'h00;      memory[14759] <=  8'h00;      memory[14760] <=  8'h00;      memory[14761] <=  8'h00;      memory[14762] <=  8'h00;      memory[14763] <=  8'h00;      memory[14764] <=  8'h00;      memory[14765] <=  8'h00;      memory[14766] <=  8'h00;      memory[14767] <=  8'h00;      memory[14768] <=  8'h00;      memory[14769] <=  8'h00;      memory[14770] <=  8'h00;      memory[14771] <=  8'h00;      memory[14772] <=  8'h00;      memory[14773] <=  8'h00;      memory[14774] <=  8'h00;      memory[14775] <=  8'h00;      memory[14776] <=  8'h00;      memory[14777] <=  8'h00;      memory[14778] <=  8'h00;      memory[14779] <=  8'h00;      memory[14780] <=  8'h00;      memory[14781] <=  8'h00;      memory[14782] <=  8'h00;      memory[14783] <=  8'h00;      memory[14784] <=  8'h00;      memory[14785] <=  8'h00;      memory[14786] <=  8'h00;      memory[14787] <=  8'h00;      memory[14788] <=  8'h00;      memory[14789] <=  8'h00;      memory[14790] <=  8'h00;      memory[14791] <=  8'h00;      memory[14792] <=  8'h00;      memory[14793] <=  8'h00;      memory[14794] <=  8'h00;      memory[14795] <=  8'h00;      memory[14796] <=  8'h00;      memory[14797] <=  8'h00;      memory[14798] <=  8'h00;      memory[14799] <=  8'h00;      memory[14800] <=  8'h00;      memory[14801] <=  8'h00;      memory[14802] <=  8'h00;      memory[14803] <=  8'h00;      memory[14804] <=  8'h00;      memory[14805] <=  8'h00;      memory[14806] <=  8'h00;      memory[14807] <=  8'h00;      memory[14808] <=  8'h00;      memory[14809] <=  8'h00;      memory[14810] <=  8'h00;      memory[14811] <=  8'h00;      memory[14812] <=  8'h00;      memory[14813] <=  8'h00;      memory[14814] <=  8'h00;      memory[14815] <=  8'h00;      memory[14816] <=  8'h00;      memory[14817] <=  8'h00;      memory[14818] <=  8'h00;      memory[14819] <=  8'h00;      memory[14820] <=  8'h00;      memory[14821] <=  8'h00;      memory[14822] <=  8'h00;      memory[14823] <=  8'h00;      memory[14824] <=  8'h00;      memory[14825] <=  8'h00;      memory[14826] <=  8'h00;      memory[14827] <=  8'h00;      memory[14828] <=  8'h00;      memory[14829] <=  8'h00;      memory[14830] <=  8'h00;      memory[14831] <=  8'h00;      memory[14832] <=  8'h00;      memory[14833] <=  8'h00;      memory[14834] <=  8'h00;      memory[14835] <=  8'h00;      memory[14836] <=  8'h00;      memory[14837] <=  8'h00;      memory[14838] <=  8'h00;      memory[14839] <=  8'h00;      memory[14840] <=  8'h00;      memory[14841] <=  8'h00;      memory[14842] <=  8'h00;      memory[14843] <=  8'h00;      memory[14844] <=  8'h00;      memory[14845] <=  8'h00;      memory[14846] <=  8'h00;      memory[14847] <=  8'h00;      memory[14848] <=  8'h00;      memory[14849] <=  8'h00;      memory[14850] <=  8'h00;      memory[14851] <=  8'h00;      memory[14852] <=  8'h00;      memory[14853] <=  8'h00;      memory[14854] <=  8'h00;      memory[14855] <=  8'h00;      memory[14856] <=  8'h00;      memory[14857] <=  8'h00;      memory[14858] <=  8'h00;      memory[14859] <=  8'h00;      memory[14860] <=  8'h00;      memory[14861] <=  8'h00;      memory[14862] <=  8'h00;      memory[14863] <=  8'h00;      memory[14864] <=  8'h00;      memory[14865] <=  8'h00;      memory[14866] <=  8'h00;      memory[14867] <=  8'h00;      memory[14868] <=  8'h00;      memory[14869] <=  8'h00;      memory[14870] <=  8'h00;      memory[14871] <=  8'h00;      memory[14872] <=  8'h00;      memory[14873] <=  8'h00;      memory[14874] <=  8'h00;      memory[14875] <=  8'h00;      memory[14876] <=  8'h00;      memory[14877] <=  8'h00;      memory[14878] <=  8'h00;      memory[14879] <=  8'h00;      memory[14880] <=  8'h00;      memory[14881] <=  8'h00;      memory[14882] <=  8'h00;      memory[14883] <=  8'h00;      memory[14884] <=  8'h00;      memory[14885] <=  8'h00;      memory[14886] <=  8'h00;      memory[14887] <=  8'h00;      memory[14888] <=  8'h00;      memory[14889] <=  8'h00;      memory[14890] <=  8'h00;      memory[14891] <=  8'h00;      memory[14892] <=  8'h00;      memory[14893] <=  8'h00;      memory[14894] <=  8'h00;      memory[14895] <=  8'h00;      memory[14896] <=  8'h00;      memory[14897] <=  8'h00;      memory[14898] <=  8'h00;      memory[14899] <=  8'h00;      memory[14900] <=  8'h00;      memory[14901] <=  8'h00;      memory[14902] <=  8'h00;      memory[14903] <=  8'h00;      memory[14904] <=  8'h00;      memory[14905] <=  8'h00;      memory[14906] <=  8'h00;      memory[14907] <=  8'h00;      memory[14908] <=  8'h00;      memory[14909] <=  8'h00;      memory[14910] <=  8'h00;      memory[14911] <=  8'h00;      memory[14912] <=  8'h00;      memory[14913] <=  8'h00;      memory[14914] <=  8'h00;      memory[14915] <=  8'h00;      memory[14916] <=  8'h00;      memory[14917] <=  8'h00;      memory[14918] <=  8'h00;      memory[14919] <=  8'h00;      memory[14920] <=  8'h00;      memory[14921] <=  8'h00;      memory[14922] <=  8'h00;      memory[14923] <=  8'h00;      memory[14924] <=  8'h00;      memory[14925] <=  8'h00;      memory[14926] <=  8'h00;      memory[14927] <=  8'h00;      memory[14928] <=  8'h00;      memory[14929] <=  8'h00;      memory[14930] <=  8'h00;      memory[14931] <=  8'h00;      memory[14932] <=  8'h00;      memory[14933] <=  8'h00;      memory[14934] <=  8'h00;      memory[14935] <=  8'h00;      memory[14936] <=  8'h00;      memory[14937] <=  8'h00;      memory[14938] <=  8'h00;      memory[14939] <=  8'h00;      memory[14940] <=  8'h00;      memory[14941] <=  8'h00;      memory[14942] <=  8'h00;      memory[14943] <=  8'h00;      memory[14944] <=  8'h00;      memory[14945] <=  8'h00;      memory[14946] <=  8'h00;      memory[14947] <=  8'h00;      memory[14948] <=  8'h00;      memory[14949] <=  8'h00;      memory[14950] <=  8'h00;      memory[14951] <=  8'h00;      memory[14952] <=  8'h00;      memory[14953] <=  8'h00;      memory[14954] <=  8'h00;      memory[14955] <=  8'h00;      memory[14956] <=  8'h00;      memory[14957] <=  8'h00;      memory[14958] <=  8'h00;      memory[14959] <=  8'h00;      memory[14960] <=  8'h00;      memory[14961] <=  8'h00;      memory[14962] <=  8'h00;      memory[14963] <=  8'h00;      memory[14964] <=  8'h00;      memory[14965] <=  8'h00;      memory[14966] <=  8'h00;      memory[14967] <=  8'h00;      memory[14968] <=  8'h00;      memory[14969] <=  8'h00;      memory[14970] <=  8'h00;      memory[14971] <=  8'h00;      memory[14972] <=  8'h00;      memory[14973] <=  8'h00;      memory[14974] <=  8'h00;      memory[14975] <=  8'h00;      memory[14976] <=  8'h00;      memory[14977] <=  8'h00;      memory[14978] <=  8'h00;      memory[14979] <=  8'h00;      memory[14980] <=  8'h00;      memory[14981] <=  8'h00;      memory[14982] <=  8'h00;      memory[14983] <=  8'h00;      memory[14984] <=  8'h00;      memory[14985] <=  8'h00;      memory[14986] <=  8'h00;      memory[14987] <=  8'h00;      memory[14988] <=  8'h00;      memory[14989] <=  8'h00;      memory[14990] <=  8'h00;      memory[14991] <=  8'h00;      memory[14992] <=  8'h00;      memory[14993] <=  8'h00;      memory[14994] <=  8'h00;      memory[14995] <=  8'h00;      memory[14996] <=  8'h00;      memory[14997] <=  8'h00;      memory[14998] <=  8'h00;      memory[14999] <=  8'h00;      memory[15000] <=  8'h00;      memory[15001] <=  8'h00;      memory[15002] <=  8'h00;      memory[15003] <=  8'h00;      memory[15004] <=  8'h00;      memory[15005] <=  8'h00;      memory[15006] <=  8'h00;      memory[15007] <=  8'h00;      memory[15008] <=  8'h00;      memory[15009] <=  8'h00;      memory[15010] <=  8'h00;      memory[15011] <=  8'h00;      memory[15012] <=  8'h00;      memory[15013] <=  8'h00;      memory[15014] <=  8'h00;      memory[15015] <=  8'h00;      memory[15016] <=  8'h00;      memory[15017] <=  8'h00;      memory[15018] <=  8'h00;      memory[15019] <=  8'h00;      memory[15020] <=  8'h00;      memory[15021] <=  8'h00;      memory[15022] <=  8'h00;      memory[15023] <=  8'h00;      memory[15024] <=  8'h00;      memory[15025] <=  8'h00;      memory[15026] <=  8'h00;      memory[15027] <=  8'h00;      memory[15028] <=  8'h00;      memory[15029] <=  8'h00;      memory[15030] <=  8'h00;      memory[15031] <=  8'h00;      memory[15032] <=  8'h00;      memory[15033] <=  8'h00;      memory[15034] <=  8'h00;      memory[15035] <=  8'h00;      memory[15036] <=  8'h00;      memory[15037] <=  8'h00;      memory[15038] <=  8'h00;      memory[15039] <=  8'h00;      memory[15040] <=  8'h00;      memory[15041] <=  8'h00;      memory[15042] <=  8'h00;      memory[15043] <=  8'h00;      memory[15044] <=  8'h00;      memory[15045] <=  8'h00;      memory[15046] <=  8'h00;      memory[15047] <=  8'h00;      memory[15048] <=  8'h00;      memory[15049] <=  8'h00;      memory[15050] <=  8'h00;      memory[15051] <=  8'h00;      memory[15052] <=  8'h00;      memory[15053] <=  8'h00;      memory[15054] <=  8'h00;      memory[15055] <=  8'h00;      memory[15056] <=  8'h00;      memory[15057] <=  8'h00;      memory[15058] <=  8'h00;      memory[15059] <=  8'h00;      memory[15060] <=  8'h00;      memory[15061] <=  8'h00;      memory[15062] <=  8'h00;      memory[15063] <=  8'h00;      memory[15064] <=  8'h00;      memory[15065] <=  8'h00;      memory[15066] <=  8'h00;      memory[15067] <=  8'h00;      memory[15068] <=  8'h00;      memory[15069] <=  8'h00;      memory[15070] <=  8'h00;      memory[15071] <=  8'h00;      memory[15072] <=  8'h00;      memory[15073] <=  8'h00;      memory[15074] <=  8'h00;      memory[15075] <=  8'h00;      memory[15076] <=  8'h00;      memory[15077] <=  8'h00;      memory[15078] <=  8'h00;      memory[15079] <=  8'h00;      memory[15080] <=  8'h00;      memory[15081] <=  8'h00;      memory[15082] <=  8'h00;      memory[15083] <=  8'h00;      memory[15084] <=  8'h00;      memory[15085] <=  8'h00;      memory[15086] <=  8'h00;      memory[15087] <=  8'h00;      memory[15088] <=  8'h00;      memory[15089] <=  8'h00;      memory[15090] <=  8'h00;      memory[15091] <=  8'h00;      memory[15092] <=  8'h00;      memory[15093] <=  8'h00;      memory[15094] <=  8'h00;      memory[15095] <=  8'h00;      memory[15096] <=  8'h00;      memory[15097] <=  8'h00;      memory[15098] <=  8'h00;      memory[15099] <=  8'h00;      memory[15100] <=  8'h00;      memory[15101] <=  8'h00;      memory[15102] <=  8'h00;      memory[15103] <=  8'h00;      memory[15104] <=  8'h00;      memory[15105] <=  8'h00;      memory[15106] <=  8'h00;      memory[15107] <=  8'h00;      memory[15108] <=  8'h00;      memory[15109] <=  8'h00;      memory[15110] <=  8'h00;      memory[15111] <=  8'h00;      memory[15112] <=  8'h00;      memory[15113] <=  8'h00;      memory[15114] <=  8'h00;      memory[15115] <=  8'h00;      memory[15116] <=  8'h00;      memory[15117] <=  8'h00;      memory[15118] <=  8'h00;      memory[15119] <=  8'h00;      memory[15120] <=  8'h00;      memory[15121] <=  8'h00;      memory[15122] <=  8'h00;      memory[15123] <=  8'h00;      memory[15124] <=  8'h00;      memory[15125] <=  8'h00;      memory[15126] <=  8'h00;      memory[15127] <=  8'h00;      memory[15128] <=  8'h00;      memory[15129] <=  8'h00;      memory[15130] <=  8'h00;      memory[15131] <=  8'h00;      memory[15132] <=  8'h00;      memory[15133] <=  8'h00;      memory[15134] <=  8'h00;      memory[15135] <=  8'h00;      memory[15136] <=  8'h00;      memory[15137] <=  8'h00;      memory[15138] <=  8'h00;      memory[15139] <=  8'h00;      memory[15140] <=  8'h00;      memory[15141] <=  8'h00;      memory[15142] <=  8'h00;      memory[15143] <=  8'h00;      memory[15144] <=  8'h00;      memory[15145] <=  8'h00;      memory[15146] <=  8'h00;      memory[15147] <=  8'h00;      memory[15148] <=  8'h00;      memory[15149] <=  8'h00;      memory[15150] <=  8'h00;      memory[15151] <=  8'h00;      memory[15152] <=  8'h00;      memory[15153] <=  8'h00;      memory[15154] <=  8'h00;      memory[15155] <=  8'h00;      memory[15156] <=  8'h00;      memory[15157] <=  8'h00;      memory[15158] <=  8'h00;      memory[15159] <=  8'h00;      memory[15160] <=  8'h00;      memory[15161] <=  8'h00;      memory[15162] <=  8'h00;      memory[15163] <=  8'h00;      memory[15164] <=  8'h00;      memory[15165] <=  8'h00;      memory[15166] <=  8'h00;      memory[15167] <=  8'h00;      memory[15168] <=  8'h00;      memory[15169] <=  8'h00;      memory[15170] <=  8'h00;      memory[15171] <=  8'h00;      memory[15172] <=  8'h00;      memory[15173] <=  8'h00;      memory[15174] <=  8'h00;      memory[15175] <=  8'h00;      memory[15176] <=  8'h00;      memory[15177] <=  8'h00;      memory[15178] <=  8'h00;      memory[15179] <=  8'h00;      memory[15180] <=  8'h00;      memory[15181] <=  8'h00;      memory[15182] <=  8'h00;      memory[15183] <=  8'h00;      memory[15184] <=  8'h00;      memory[15185] <=  8'h00;      memory[15186] <=  8'h00;      memory[15187] <=  8'h00;      memory[15188] <=  8'h00;      memory[15189] <=  8'h00;      memory[15190] <=  8'h00;      memory[15191] <=  8'h00;      memory[15192] <=  8'h00;      memory[15193] <=  8'h00;      memory[15194] <=  8'h00;      memory[15195] <=  8'h00;      memory[15196] <=  8'h00;      memory[15197] <=  8'h00;      memory[15198] <=  8'h00;      memory[15199] <=  8'h00;      memory[15200] <=  8'h00;      memory[15201] <=  8'h00;      memory[15202] <=  8'h00;      memory[15203] <=  8'h00;      memory[15204] <=  8'h00;      memory[15205] <=  8'h00;      memory[15206] <=  8'h00;      memory[15207] <=  8'h00;      memory[15208] <=  8'h00;      memory[15209] <=  8'h00;      memory[15210] <=  8'h00;      memory[15211] <=  8'h00;      memory[15212] <=  8'h00;      memory[15213] <=  8'h00;      memory[15214] <=  8'h00;      memory[15215] <=  8'h00;      memory[15216] <=  8'h00;      memory[15217] <=  8'h00;      memory[15218] <=  8'h00;      memory[15219] <=  8'h00;      memory[15220] <=  8'h00;      memory[15221] <=  8'h00;      memory[15222] <=  8'h00;      memory[15223] <=  8'h00;      memory[15224] <=  8'h00;      memory[15225] <=  8'h00;      memory[15226] <=  8'h00;      memory[15227] <=  8'h00;      memory[15228] <=  8'h00;      memory[15229] <=  8'h00;      memory[15230] <=  8'h00;      memory[15231] <=  8'h00;      memory[15232] <=  8'h00;      memory[15233] <=  8'h00;      memory[15234] <=  8'h00;      memory[15235] <=  8'h00;      memory[15236] <=  8'h00;      memory[15237] <=  8'h00;      memory[15238] <=  8'h00;      memory[15239] <=  8'h00;      memory[15240] <=  8'h00;      memory[15241] <=  8'h00;      memory[15242] <=  8'h00;      memory[15243] <=  8'h00;      memory[15244] <=  8'h00;      memory[15245] <=  8'h00;      memory[15246] <=  8'h00;      memory[15247] <=  8'h00;      memory[15248] <=  8'h00;      memory[15249] <=  8'h00;      memory[15250] <=  8'h00;      memory[15251] <=  8'h00;      memory[15252] <=  8'h00;      memory[15253] <=  8'h00;      memory[15254] <=  8'h00;      memory[15255] <=  8'h00;      memory[15256] <=  8'h00;      memory[15257] <=  8'h00;      memory[15258] <=  8'h00;      memory[15259] <=  8'h00;      memory[15260] <=  8'h00;      memory[15261] <=  8'h00;      memory[15262] <=  8'h00;      memory[15263] <=  8'h00;      memory[15264] <=  8'h00;      memory[15265] <=  8'h00;      memory[15266] <=  8'h00;      memory[15267] <=  8'h00;      memory[15268] <=  8'h00;      memory[15269] <=  8'h00;      memory[15270] <=  8'h00;      memory[15271] <=  8'h00;      memory[15272] <=  8'h00;      memory[15273] <=  8'h00;      memory[15274] <=  8'h00;      memory[15275] <=  8'h00;      memory[15276] <=  8'h00;      memory[15277] <=  8'h00;      memory[15278] <=  8'h00;      memory[15279] <=  8'h00;      memory[15280] <=  8'h00;      memory[15281] <=  8'h00;      memory[15282] <=  8'h00;      memory[15283] <=  8'h00;      memory[15284] <=  8'h00;      memory[15285] <=  8'h00;      memory[15286] <=  8'h00;      memory[15287] <=  8'h00;      memory[15288] <=  8'h00;      memory[15289] <=  8'h00;      memory[15290] <=  8'h00;      memory[15291] <=  8'h00;      memory[15292] <=  8'h00;      memory[15293] <=  8'h00;      memory[15294] <=  8'h00;      memory[15295] <=  8'h00;      memory[15296] <=  8'h00;      memory[15297] <=  8'h00;      memory[15298] <=  8'h00;      memory[15299] <=  8'h00;      memory[15300] <=  8'h00;      memory[15301] <=  8'h00;      memory[15302] <=  8'h00;      memory[15303] <=  8'h00;      memory[15304] <=  8'h00;      memory[15305] <=  8'h00;      memory[15306] <=  8'h00;      memory[15307] <=  8'h00;      memory[15308] <=  8'h00;      memory[15309] <=  8'h00;      memory[15310] <=  8'h00;      memory[15311] <=  8'h00;      memory[15312] <=  8'h00;      memory[15313] <=  8'h00;      memory[15314] <=  8'h00;      memory[15315] <=  8'h00;      memory[15316] <=  8'h00;      memory[15317] <=  8'h00;      memory[15318] <=  8'h00;      memory[15319] <=  8'h00;      memory[15320] <=  8'h00;      memory[15321] <=  8'h00;      memory[15322] <=  8'h00;      memory[15323] <=  8'h00;      memory[15324] <=  8'h00;      memory[15325] <=  8'h00;      memory[15326] <=  8'h00;      memory[15327] <=  8'h00;      memory[15328] <=  8'h00;      memory[15329] <=  8'h00;      memory[15330] <=  8'h00;      memory[15331] <=  8'h00;      memory[15332] <=  8'h00;      memory[15333] <=  8'h00;      memory[15334] <=  8'h00;      memory[15335] <=  8'h00;      memory[15336] <=  8'h00;      memory[15337] <=  8'h00;      memory[15338] <=  8'h00;      memory[15339] <=  8'h00;      memory[15340] <=  8'h00;      memory[15341] <=  8'h00;      memory[15342] <=  8'h00;      memory[15343] <=  8'h00;      memory[15344] <=  8'h00;      memory[15345] <=  8'h00;      memory[15346] <=  8'h00;      memory[15347] <=  8'h00;      memory[15348] <=  8'h00;      memory[15349] <=  8'h00;      memory[15350] <=  8'h00;      memory[15351] <=  8'h00;      memory[15352] <=  8'h00;      memory[15353] <=  8'h00;      memory[15354] <=  8'h00;      memory[15355] <=  8'h00;      memory[15356] <=  8'h00;      memory[15357] <=  8'h00;      memory[15358] <=  8'h00;      memory[15359] <=  8'h00;      memory[15360] <=  8'h00;      memory[15361] <=  8'h00;      memory[15362] <=  8'h00;      memory[15363] <=  8'h00;      memory[15364] <=  8'h00;      memory[15365] <=  8'h00;      memory[15366] <=  8'h00;      memory[15367] <=  8'h00;      memory[15368] <=  8'h00;      memory[15369] <=  8'h00;      memory[15370] <=  8'h00;      memory[15371] <=  8'h00;      memory[15372] <=  8'h00;      memory[15373] <=  8'h00;      memory[15374] <=  8'h00;      memory[15375] <=  8'h00;      memory[15376] <=  8'h00;      memory[15377] <=  8'h00;      memory[15378] <=  8'h00;      memory[15379] <=  8'h00;      memory[15380] <=  8'h00;      memory[15381] <=  8'h00;      memory[15382] <=  8'h00;      memory[15383] <=  8'h00;      memory[15384] <=  8'h00;      memory[15385] <=  8'h00;      memory[15386] <=  8'h00;      memory[15387] <=  8'h00;      memory[15388] <=  8'h00;      memory[15389] <=  8'h00;      memory[15390] <=  8'h00;      memory[15391] <=  8'h00;      memory[15392] <=  8'h00;      memory[15393] <=  8'h00;      memory[15394] <=  8'h00;      memory[15395] <=  8'h00;      memory[15396] <=  8'h00;      memory[15397] <=  8'h00;      memory[15398] <=  8'h00;      memory[15399] <=  8'h00;      memory[15400] <=  8'h00;      memory[15401] <=  8'h00;      memory[15402] <=  8'h00;      memory[15403] <=  8'h00;      memory[15404] <=  8'h00;      memory[15405] <=  8'h00;      memory[15406] <=  8'h00;      memory[15407] <=  8'h00;      memory[15408] <=  8'h00;      memory[15409] <=  8'h00;      memory[15410] <=  8'h00;      memory[15411] <=  8'h00;      memory[15412] <=  8'h00;      memory[15413] <=  8'h00;      memory[15414] <=  8'h00;      memory[15415] <=  8'h00;      memory[15416] <=  8'h00;      memory[15417] <=  8'h00;      memory[15418] <=  8'h00;      memory[15419] <=  8'h00;      memory[15420] <=  8'h00;      memory[15421] <=  8'h00;      memory[15422] <=  8'h00;      memory[15423] <=  8'h00;      memory[15424] <=  8'h00;      memory[15425] <=  8'h00;      memory[15426] <=  8'h00;      memory[15427] <=  8'h00;      memory[15428] <=  8'h00;      memory[15429] <=  8'h00;      memory[15430] <=  8'h00;      memory[15431] <=  8'h00;      memory[15432] <=  8'h00;      memory[15433] <=  8'h00;      memory[15434] <=  8'h00;      memory[15435] <=  8'h00;      memory[15436] <=  8'h00;      memory[15437] <=  8'h00;      memory[15438] <=  8'h00;      memory[15439] <=  8'h00;      memory[15440] <=  8'h00;      memory[15441] <=  8'h00;      memory[15442] <=  8'h00;      memory[15443] <=  8'h00;      memory[15444] <=  8'h00;      memory[15445] <=  8'h00;      memory[15446] <=  8'h00;      memory[15447] <=  8'h00;      memory[15448] <=  8'h00;      memory[15449] <=  8'h00;      memory[15450] <=  8'h00;      memory[15451] <=  8'h00;      memory[15452] <=  8'h00;      memory[15453] <=  8'h00;      memory[15454] <=  8'h00;      memory[15455] <=  8'h00;      memory[15456] <=  8'h00;      memory[15457] <=  8'h00;      memory[15458] <=  8'h00;      memory[15459] <=  8'h00;      memory[15460] <=  8'h00;      memory[15461] <=  8'h00;      memory[15462] <=  8'h00;      memory[15463] <=  8'h00;      memory[15464] <=  8'h00;      memory[15465] <=  8'h00;      memory[15466] <=  8'h00;      memory[15467] <=  8'h00;      memory[15468] <=  8'h00;      memory[15469] <=  8'h00;      memory[15470] <=  8'h00;      memory[15471] <=  8'h00;      memory[15472] <=  8'h00;      memory[15473] <=  8'h00;      memory[15474] <=  8'h00;      memory[15475] <=  8'h00;      memory[15476] <=  8'h00;      memory[15477] <=  8'h00;      memory[15478] <=  8'h00;      memory[15479] <=  8'h00;      memory[15480] <=  8'h00;      memory[15481] <=  8'h00;      memory[15482] <=  8'h00;      memory[15483] <=  8'h00;      memory[15484] <=  8'h00;      memory[15485] <=  8'h00;      memory[15486] <=  8'h00;      memory[15487] <=  8'h00;      memory[15488] <=  8'h00;      memory[15489] <=  8'h00;      memory[15490] <=  8'h00;      memory[15491] <=  8'h00;      memory[15492] <=  8'h00;      memory[15493] <=  8'h00;      memory[15494] <=  8'h00;      memory[15495] <=  8'h00;      memory[15496] <=  8'h00;      memory[15497] <=  8'h00;      memory[15498] <=  8'h00;      memory[15499] <=  8'h00;      memory[15500] <=  8'h00;      memory[15501] <=  8'h00;      memory[15502] <=  8'h00;      memory[15503] <=  8'h00;      memory[15504] <=  8'h00;      memory[15505] <=  8'h00;      memory[15506] <=  8'h00;      memory[15507] <=  8'h00;      memory[15508] <=  8'h00;      memory[15509] <=  8'h00;      memory[15510] <=  8'h00;      memory[15511] <=  8'h00;      memory[15512] <=  8'h00;      memory[15513] <=  8'h00;      memory[15514] <=  8'h00;      memory[15515] <=  8'h00;      memory[15516] <=  8'h00;      memory[15517] <=  8'h00;      memory[15518] <=  8'h00;      memory[15519] <=  8'h00;      memory[15520] <=  8'h00;      memory[15521] <=  8'h00;      memory[15522] <=  8'h00;      memory[15523] <=  8'h00;      memory[15524] <=  8'h00;      memory[15525] <=  8'h00;      memory[15526] <=  8'h00;      memory[15527] <=  8'h00;      memory[15528] <=  8'h00;      memory[15529] <=  8'h00;      memory[15530] <=  8'h00;      memory[15531] <=  8'h00;      memory[15532] <=  8'h00;      memory[15533] <=  8'h00;      memory[15534] <=  8'h00;      memory[15535] <=  8'h00;      memory[15536] <=  8'h00;      memory[15537] <=  8'h00;      memory[15538] <=  8'h00;      memory[15539] <=  8'h00;      memory[15540] <=  8'h00;      memory[15541] <=  8'h00;      memory[15542] <=  8'h00;      memory[15543] <=  8'h00;      memory[15544] <=  8'h00;      memory[15545] <=  8'h00;      memory[15546] <=  8'h00;      memory[15547] <=  8'h00;      memory[15548] <=  8'h00;      memory[15549] <=  8'h00;      memory[15550] <=  8'h00;      memory[15551] <=  8'h00;      memory[15552] <=  8'h00;      memory[15553] <=  8'h00;      memory[15554] <=  8'h00;      memory[15555] <=  8'h00;      memory[15556] <=  8'h00;      memory[15557] <=  8'h00;      memory[15558] <=  8'h00;      memory[15559] <=  8'h00;      memory[15560] <=  8'h00;      memory[15561] <=  8'h00;      memory[15562] <=  8'h00;      memory[15563] <=  8'h00;      memory[15564] <=  8'h00;      memory[15565] <=  8'h00;      memory[15566] <=  8'h00;      memory[15567] <=  8'h00;      memory[15568] <=  8'h00;      memory[15569] <=  8'h00;      memory[15570] <=  8'h00;      memory[15571] <=  8'h00;      memory[15572] <=  8'h00;      memory[15573] <=  8'h00;      memory[15574] <=  8'h00;      memory[15575] <=  8'h00;      memory[15576] <=  8'h00;      memory[15577] <=  8'h00;      memory[15578] <=  8'h00;      memory[15579] <=  8'h00;      memory[15580] <=  8'h00;      memory[15581] <=  8'h00;      memory[15582] <=  8'h00;      memory[15583] <=  8'h00;      memory[15584] <=  8'h00;      memory[15585] <=  8'h00;      memory[15586] <=  8'h00;      memory[15587] <=  8'h00;      memory[15588] <=  8'h00;      memory[15589] <=  8'h00;      memory[15590] <=  8'h00;      memory[15591] <=  8'h00;      memory[15592] <=  8'h00;      memory[15593] <=  8'h00;      memory[15594] <=  8'h00;      memory[15595] <=  8'h00;      memory[15596] <=  8'h00;      memory[15597] <=  8'h00;      memory[15598] <=  8'h00;      memory[15599] <=  8'h00;      memory[15600] <=  8'h00;      memory[15601] <=  8'h00;      memory[15602] <=  8'h00;      memory[15603] <=  8'h00;      memory[15604] <=  8'h00;      memory[15605] <=  8'h00;      memory[15606] <=  8'h00;      memory[15607] <=  8'h00;      memory[15608] <=  8'h00;      memory[15609] <=  8'h00;      memory[15610] <=  8'h00;      memory[15611] <=  8'h00;      memory[15612] <=  8'h00;      memory[15613] <=  8'h00;      memory[15614] <=  8'h00;      memory[15615] <=  8'h00;      memory[15616] <=  8'h00;      memory[15617] <=  8'h00;      memory[15618] <=  8'h00;      memory[15619] <=  8'h00;      memory[15620] <=  8'h00;      memory[15621] <=  8'h00;      memory[15622] <=  8'h00;      memory[15623] <=  8'h00;      memory[15624] <=  8'h00;      memory[15625] <=  8'h00;      memory[15626] <=  8'h00;      memory[15627] <=  8'h00;      memory[15628] <=  8'h00;      memory[15629] <=  8'h00;      memory[15630] <=  8'h00;      memory[15631] <=  8'h00;      memory[15632] <=  8'h00;      memory[15633] <=  8'h00;      memory[15634] <=  8'h00;      memory[15635] <=  8'h00;      memory[15636] <=  8'h00;      memory[15637] <=  8'h00;      memory[15638] <=  8'h00;      memory[15639] <=  8'h00;      memory[15640] <=  8'h00;      memory[15641] <=  8'h00;      memory[15642] <=  8'h00;      memory[15643] <=  8'h00;      memory[15644] <=  8'h00;      memory[15645] <=  8'h00;      memory[15646] <=  8'h00;      memory[15647] <=  8'h00;      memory[15648] <=  8'h00;      memory[15649] <=  8'h00;      memory[15650] <=  8'h00;      memory[15651] <=  8'h00;      memory[15652] <=  8'h00;      memory[15653] <=  8'h00;      memory[15654] <=  8'h00;      memory[15655] <=  8'h00;      memory[15656] <=  8'h00;      memory[15657] <=  8'h00;      memory[15658] <=  8'h00;      memory[15659] <=  8'h00;      memory[15660] <=  8'h00;      memory[15661] <=  8'h00;      memory[15662] <=  8'h00;      memory[15663] <=  8'h00;      memory[15664] <=  8'h00;      memory[15665] <=  8'h00;      memory[15666] <=  8'h00;      memory[15667] <=  8'h00;      memory[15668] <=  8'h00;      memory[15669] <=  8'h00;      memory[15670] <=  8'h00;      memory[15671] <=  8'h00;      memory[15672] <=  8'h00;      memory[15673] <=  8'h00;      memory[15674] <=  8'h00;      memory[15675] <=  8'h00;      memory[15676] <=  8'h00;      memory[15677] <=  8'h00;      memory[15678] <=  8'h00;      memory[15679] <=  8'h00;      memory[15680] <=  8'h00;      memory[15681] <=  8'h00;      memory[15682] <=  8'h00;      memory[15683] <=  8'h00;      memory[15684] <=  8'h00;      memory[15685] <=  8'h00;      memory[15686] <=  8'h00;      memory[15687] <=  8'h00;      memory[15688] <=  8'h00;      memory[15689] <=  8'h00;      memory[15690] <=  8'h00;      memory[15691] <=  8'h00;      memory[15692] <=  8'h00;      memory[15693] <=  8'h00;      memory[15694] <=  8'h00;      memory[15695] <=  8'h00;      memory[15696] <=  8'h00;      memory[15697] <=  8'h00;      memory[15698] <=  8'h00;      memory[15699] <=  8'h00;      memory[15700] <=  8'h00;      memory[15701] <=  8'h00;      memory[15702] <=  8'h00;      memory[15703] <=  8'h00;      memory[15704] <=  8'h00;      memory[15705] <=  8'h00;      memory[15706] <=  8'h00;      memory[15707] <=  8'h00;      memory[15708] <=  8'h00;      memory[15709] <=  8'h00;      memory[15710] <=  8'h00;      memory[15711] <=  8'h00;      memory[15712] <=  8'h00;      memory[15713] <=  8'h00;      memory[15714] <=  8'h00;      memory[15715] <=  8'h00;      memory[15716] <=  8'h00;      memory[15717] <=  8'h00;      memory[15718] <=  8'h00;      memory[15719] <=  8'h00;      memory[15720] <=  8'h00;      memory[15721] <=  8'h00;      memory[15722] <=  8'h00;      memory[15723] <=  8'h00;      memory[15724] <=  8'h00;      memory[15725] <=  8'h00;      memory[15726] <=  8'h00;      memory[15727] <=  8'h00;      memory[15728] <=  8'h00;      memory[15729] <=  8'h00;      memory[15730] <=  8'h00;      memory[15731] <=  8'h00;      memory[15732] <=  8'h00;      memory[15733] <=  8'h00;      memory[15734] <=  8'h00;      memory[15735] <=  8'h00;      memory[15736] <=  8'h00;      memory[15737] <=  8'h00;      memory[15738] <=  8'h00;      memory[15739] <=  8'h00;      memory[15740] <=  8'h00;      memory[15741] <=  8'h00;      memory[15742] <=  8'h00;      memory[15743] <=  8'h00;      memory[15744] <=  8'h00;      memory[15745] <=  8'h00;      memory[15746] <=  8'h00;      memory[15747] <=  8'h00;      memory[15748] <=  8'h00;      memory[15749] <=  8'h00;      memory[15750] <=  8'h00;      memory[15751] <=  8'h00;      memory[15752] <=  8'h00;      memory[15753] <=  8'h00;      memory[15754] <=  8'h00;      memory[15755] <=  8'h00;      memory[15756] <=  8'h00;      memory[15757] <=  8'h00;      memory[15758] <=  8'h00;      memory[15759] <=  8'h00;      memory[15760] <=  8'h00;      memory[15761] <=  8'h00;      memory[15762] <=  8'h00;      memory[15763] <=  8'h00;      memory[15764] <=  8'h00;      memory[15765] <=  8'h00;      memory[15766] <=  8'h00;      memory[15767] <=  8'h00;      memory[15768] <=  8'h00;      memory[15769] <=  8'h00;      memory[15770] <=  8'h00;      memory[15771] <=  8'h00;      memory[15772] <=  8'h00;      memory[15773] <=  8'h00;      memory[15774] <=  8'h00;      memory[15775] <=  8'h00;      memory[15776] <=  8'h00;      memory[15777] <=  8'h00;      memory[15778] <=  8'h00;      memory[15779] <=  8'h00;      memory[15780] <=  8'h00;      memory[15781] <=  8'h00;      memory[15782] <=  8'h00;      memory[15783] <=  8'h00;      memory[15784] <=  8'h00;      memory[15785] <=  8'h00;      memory[15786] <=  8'h00;      memory[15787] <=  8'h00;      memory[15788] <=  8'h00;      memory[15789] <=  8'h00;      memory[15790] <=  8'h00;      memory[15791] <=  8'h00;      memory[15792] <=  8'h00;      memory[15793] <=  8'h00;      memory[15794] <=  8'h00;      memory[15795] <=  8'h00;      memory[15796] <=  8'h00;      memory[15797] <=  8'h00;      memory[15798] <=  8'h00;      memory[15799] <=  8'h00;      memory[15800] <=  8'h00;      memory[15801] <=  8'h00;      memory[15802] <=  8'h00;      memory[15803] <=  8'h00;      memory[15804] <=  8'h00;      memory[15805] <=  8'h00;      memory[15806] <=  8'h00;      memory[15807] <=  8'h00;      memory[15808] <=  8'h00;      memory[15809] <=  8'h00;      memory[15810] <=  8'h00;      memory[15811] <=  8'h00;      memory[15812] <=  8'h00;      memory[15813] <=  8'h00;      memory[15814] <=  8'h00;      memory[15815] <=  8'h00;      memory[15816] <=  8'h00;      memory[15817] <=  8'h00;      memory[15818] <=  8'h00;      memory[15819] <=  8'h00;      memory[15820] <=  8'h00;      memory[15821] <=  8'h00;      memory[15822] <=  8'h00;      memory[15823] <=  8'h00;      memory[15824] <=  8'h00;      memory[15825] <=  8'h00;      memory[15826] <=  8'h00;      memory[15827] <=  8'h00;      memory[15828] <=  8'h00;      memory[15829] <=  8'h00;      memory[15830] <=  8'h00;      memory[15831] <=  8'h00;      memory[15832] <=  8'h00;      memory[15833] <=  8'h00;      memory[15834] <=  8'h00;      memory[15835] <=  8'h00;      memory[15836] <=  8'h00;      memory[15837] <=  8'h00;      memory[15838] <=  8'h00;      memory[15839] <=  8'h00;      memory[15840] <=  8'h00;      memory[15841] <=  8'h00;      memory[15842] <=  8'h00;      memory[15843] <=  8'h00;      memory[15844] <=  8'h00;      memory[15845] <=  8'h00;      memory[15846] <=  8'h00;      memory[15847] <=  8'h00;      memory[15848] <=  8'h00;      memory[15849] <=  8'h00;      memory[15850] <=  8'h00;      memory[15851] <=  8'h00;      memory[15852] <=  8'h00;      memory[15853] <=  8'h00;      memory[15854] <=  8'h00;      memory[15855] <=  8'h00;      memory[15856] <=  8'h00;      memory[15857] <=  8'h00;      memory[15858] <=  8'h00;      memory[15859] <=  8'h00;      memory[15860] <=  8'h00;      memory[15861] <=  8'h00;      memory[15862] <=  8'h00;      memory[15863] <=  8'h00;      memory[15864] <=  8'h00;      memory[15865] <=  8'h00;      memory[15866] <=  8'h00;      memory[15867] <=  8'h00;      memory[15868] <=  8'h00;      memory[15869] <=  8'h00;      memory[15870] <=  8'h00;      memory[15871] <=  8'h00;      memory[15872] <=  8'h00;      memory[15873] <=  8'h00;      memory[15874] <=  8'h00;      memory[15875] <=  8'h00;      memory[15876] <=  8'h00;      memory[15877] <=  8'h00;      memory[15878] <=  8'h00;      memory[15879] <=  8'h00;      memory[15880] <=  8'h00;      memory[15881] <=  8'h00;      memory[15882] <=  8'h00;      memory[15883] <=  8'h00;      memory[15884] <=  8'h00;      memory[15885] <=  8'h00;      memory[15886] <=  8'h00;      memory[15887] <=  8'h00;      memory[15888] <=  8'h00;      memory[15889] <=  8'h00;      memory[15890] <=  8'h00;      memory[15891] <=  8'h00;      memory[15892] <=  8'h00;      memory[15893] <=  8'h00;      memory[15894] <=  8'h00;      memory[15895] <=  8'h00;      memory[15896] <=  8'h00;      memory[15897] <=  8'h00;      memory[15898] <=  8'h00;      memory[15899] <=  8'h00;      memory[15900] <=  8'h00;      memory[15901] <=  8'h00;      memory[15902] <=  8'h00;      memory[15903] <=  8'h00;      memory[15904] <=  8'h00;      memory[15905] <=  8'h00;      memory[15906] <=  8'h00;      memory[15907] <=  8'h00;      memory[15908] <=  8'h00;      memory[15909] <=  8'h00;      memory[15910] <=  8'h00;      memory[15911] <=  8'h00;      memory[15912] <=  8'h00;      memory[15913] <=  8'h00;      memory[15914] <=  8'h00;      memory[15915] <=  8'h00;      memory[15916] <=  8'h00;      memory[15917] <=  8'h00;      memory[15918] <=  8'h00;      memory[15919] <=  8'h00;      memory[15920] <=  8'h00;      memory[15921] <=  8'h00;      memory[15922] <=  8'h00;      memory[15923] <=  8'h00;      memory[15924] <=  8'h00;      memory[15925] <=  8'h00;      memory[15926] <=  8'h00;      memory[15927] <=  8'h00;      memory[15928] <=  8'h00;      memory[15929] <=  8'h00;      memory[15930] <=  8'h00;      memory[15931] <=  8'h00;      memory[15932] <=  8'h00;      memory[15933] <=  8'h00;      memory[15934] <=  8'h00;      memory[15935] <=  8'h00;      memory[15936] <=  8'h00;      memory[15937] <=  8'h00;      memory[15938] <=  8'h00;      memory[15939] <=  8'h00;      memory[15940] <=  8'h00;      memory[15941] <=  8'h00;      memory[15942] <=  8'h00;      memory[15943] <=  8'h00;      memory[15944] <=  8'h00;      memory[15945] <=  8'h00;      memory[15946] <=  8'h00;      memory[15947] <=  8'h00;      memory[15948] <=  8'h00;      memory[15949] <=  8'h00;      memory[15950] <=  8'h00;      memory[15951] <=  8'h00;      memory[15952] <=  8'h00;      memory[15953] <=  8'h00;      memory[15954] <=  8'h00;      memory[15955] <=  8'h00;      memory[15956] <=  8'h00;      memory[15957] <=  8'h00;      memory[15958] <=  8'h00;      memory[15959] <=  8'h00;      memory[15960] <=  8'h00;      memory[15961] <=  8'h00;      memory[15962] <=  8'h00;      memory[15963] <=  8'h00;      memory[15964] <=  8'h00;      memory[15965] <=  8'h00;      memory[15966] <=  8'h00;      memory[15967] <=  8'h00;      memory[15968] <=  8'h00;      memory[15969] <=  8'h00;      memory[15970] <=  8'h00;      memory[15971] <=  8'h00;      memory[15972] <=  8'h00;      memory[15973] <=  8'h00;      memory[15974] <=  8'h00;      memory[15975] <=  8'h00;      memory[15976] <=  8'h00;      memory[15977] <=  8'h00;      memory[15978] <=  8'h00;      memory[15979] <=  8'h00;      memory[15980] <=  8'h00;      memory[15981] <=  8'h00;      memory[15982] <=  8'h00;      memory[15983] <=  8'h00;      memory[15984] <=  8'h00;      memory[15985] <=  8'h00;      memory[15986] <=  8'h00;      memory[15987] <=  8'h00;      memory[15988] <=  8'h00;      memory[15989] <=  8'h00;      memory[15990] <=  8'h00;      memory[15991] <=  8'h00;      memory[15992] <=  8'h00;      memory[15993] <=  8'h00;      memory[15994] <=  8'h00;      memory[15995] <=  8'h00;      memory[15996] <=  8'h00;      memory[15997] <=  8'h00;      memory[15998] <=  8'h00;      memory[15999] <=  8'h00;      memory[16000] <=  8'h00;      memory[16001] <=  8'h00;      memory[16002] <=  8'h00;      memory[16003] <=  8'h00;      memory[16004] <=  8'h00;      memory[16005] <=  8'h00;      memory[16006] <=  8'h00;      memory[16007] <=  8'h00;      memory[16008] <=  8'h00;      memory[16009] <=  8'h00;      memory[16010] <=  8'h00;      memory[16011] <=  8'h00;      memory[16012] <=  8'h00;      memory[16013] <=  8'h00;      memory[16014] <=  8'h00;      memory[16015] <=  8'h00;      memory[16016] <=  8'h00;      memory[16017] <=  8'h00;      memory[16018] <=  8'h00;      memory[16019] <=  8'h00;      memory[16020] <=  8'h00;      memory[16021] <=  8'h00;      memory[16022] <=  8'h00;      memory[16023] <=  8'h00;      memory[16024] <=  8'h00;      memory[16025] <=  8'h00;      memory[16026] <=  8'h00;      memory[16027] <=  8'h00;      memory[16028] <=  8'h00;      memory[16029] <=  8'h00;      memory[16030] <=  8'h00;      memory[16031] <=  8'h00;      memory[16032] <=  8'h00;      memory[16033] <=  8'h00;      memory[16034] <=  8'h00;      memory[16035] <=  8'h00;      memory[16036] <=  8'h00;      memory[16037] <=  8'h00;      memory[16038] <=  8'h00;      memory[16039] <=  8'h00;      memory[16040] <=  8'h00;      memory[16041] <=  8'h00;      memory[16042] <=  8'h00;      memory[16043] <=  8'h00;      memory[16044] <=  8'h00;      memory[16045] <=  8'h00;      memory[16046] <=  8'h00;      memory[16047] <=  8'h00;      memory[16048] <=  8'h00;      memory[16049] <=  8'h00;      memory[16050] <=  8'h00;      memory[16051] <=  8'h00;      memory[16052] <=  8'h00;      memory[16053] <=  8'h00;      memory[16054] <=  8'h00;      memory[16055] <=  8'h00;      memory[16056] <=  8'h00;      memory[16057] <=  8'h00;      memory[16058] <=  8'h00;      memory[16059] <=  8'h00;      memory[16060] <=  8'h00;      memory[16061] <=  8'h00;      memory[16062] <=  8'h00;      memory[16063] <=  8'h00;      memory[16064] <=  8'h00;      memory[16065] <=  8'h00;      memory[16066] <=  8'h00;      memory[16067] <=  8'h00;      memory[16068] <=  8'h00;      memory[16069] <=  8'h00;      memory[16070] <=  8'h00;      memory[16071] <=  8'h00;      memory[16072] <=  8'h00;      memory[16073] <=  8'h00;      memory[16074] <=  8'h00;      memory[16075] <=  8'h00;      memory[16076] <=  8'h00;      memory[16077] <=  8'h00;      memory[16078] <=  8'h00;      memory[16079] <=  8'h00;      memory[16080] <=  8'h00;      memory[16081] <=  8'h00;      memory[16082] <=  8'h00;      memory[16083] <=  8'h00;      memory[16084] <=  8'h00;      memory[16085] <=  8'h00;      memory[16086] <=  8'h00;      memory[16087] <=  8'h00;      memory[16088] <=  8'h00;      memory[16089] <=  8'h00;      memory[16090] <=  8'h00;      memory[16091] <=  8'h00;      memory[16092] <=  8'h00;      memory[16093] <=  8'h00;      memory[16094] <=  8'h00;      memory[16095] <=  8'h00;      memory[16096] <=  8'h00;      memory[16097] <=  8'h00;      memory[16098] <=  8'h00;      memory[16099] <=  8'h00;      memory[16100] <=  8'h00;      memory[16101] <=  8'h00;      memory[16102] <=  8'h00;      memory[16103] <=  8'h00;      memory[16104] <=  8'h00;      memory[16105] <=  8'h00;      memory[16106] <=  8'h00;      memory[16107] <=  8'h00;      memory[16108] <=  8'h00;      memory[16109] <=  8'h00;      memory[16110] <=  8'h00;      memory[16111] <=  8'h00;      memory[16112] <=  8'h00;      memory[16113] <=  8'h00;      memory[16114] <=  8'h00;      memory[16115] <=  8'h00;      memory[16116] <=  8'h00;      memory[16117] <=  8'h00;      memory[16118] <=  8'h00;      memory[16119] <=  8'h00;      memory[16120] <=  8'h00;      memory[16121] <=  8'h00;      memory[16122] <=  8'h00;      memory[16123] <=  8'h00;      memory[16124] <=  8'h00;      memory[16125] <=  8'h00;      memory[16126] <=  8'h00;      memory[16127] <=  8'h00;      memory[16128] <=  8'h00;      memory[16129] <=  8'h00;      memory[16130] <=  8'h00;      memory[16131] <=  8'h00;      memory[16132] <=  8'h00;      memory[16133] <=  8'h00;      memory[16134] <=  8'h00;      memory[16135] <=  8'h00;      memory[16136] <=  8'h00;      memory[16137] <=  8'h00;      memory[16138] <=  8'h00;      memory[16139] <=  8'h00;      memory[16140] <=  8'h00;      memory[16141] <=  8'h00;      memory[16142] <=  8'h00;      memory[16143] <=  8'h00;      memory[16144] <=  8'h00;      memory[16145] <=  8'h00;      memory[16146] <=  8'h00;      memory[16147] <=  8'h00;      memory[16148] <=  8'h00;      memory[16149] <=  8'h00;      memory[16150] <=  8'h00;      memory[16151] <=  8'h00;      memory[16152] <=  8'h00;      memory[16153] <=  8'h00;      memory[16154] <=  8'h00;      memory[16155] <=  8'h00;      memory[16156] <=  8'h00;      memory[16157] <=  8'h00;      memory[16158] <=  8'h00;      memory[16159] <=  8'h00;      memory[16160] <=  8'h00;      memory[16161] <=  8'h00;      memory[16162] <=  8'h00;      memory[16163] <=  8'h00;      memory[16164] <=  8'h00;      memory[16165] <=  8'h00;      memory[16166] <=  8'h00;      memory[16167] <=  8'h00;      memory[16168] <=  8'h00;      memory[16169] <=  8'h00;      memory[16170] <=  8'h00;      memory[16171] <=  8'h00;      memory[16172] <=  8'h00;      memory[16173] <=  8'h00;      memory[16174] <=  8'h00;      memory[16175] <=  8'h00;      memory[16176] <=  8'h00;      memory[16177] <=  8'h00;      memory[16178] <=  8'h00;      memory[16179] <=  8'h00;      memory[16180] <=  8'h00;      memory[16181] <=  8'h00;      memory[16182] <=  8'h00;      memory[16183] <=  8'h00;      memory[16184] <=  8'h00;      memory[16185] <=  8'h00;      memory[16186] <=  8'h00;      memory[16187] <=  8'h00;      memory[16188] <=  8'h00;      memory[16189] <=  8'h00;      memory[16190] <=  8'h00;      memory[16191] <=  8'h00;      memory[16192] <=  8'h00;      memory[16193] <=  8'h00;      memory[16194] <=  8'h00;      memory[16195] <=  8'h00;      memory[16196] <=  8'h00;      memory[16197] <=  8'h00;      memory[16198] <=  8'h00;      memory[16199] <=  8'h00;      memory[16200] <=  8'h00;      memory[16201] <=  8'h00;      memory[16202] <=  8'h00;      memory[16203] <=  8'h00;      memory[16204] <=  8'h00;      memory[16205] <=  8'h00;      memory[16206] <=  8'h00;      memory[16207] <=  8'h00;      memory[16208] <=  8'h00;      memory[16209] <=  8'h00;      memory[16210] <=  8'h00;      memory[16211] <=  8'h00;      memory[16212] <=  8'h00;      memory[16213] <=  8'h00;      memory[16214] <=  8'h00;      memory[16215] <=  8'h00;      memory[16216] <=  8'h00;      memory[16217] <=  8'h00;      memory[16218] <=  8'h00;      memory[16219] <=  8'h00;      memory[16220] <=  8'h00;      memory[16221] <=  8'h00;      memory[16222] <=  8'h00;      memory[16223] <=  8'h00;      memory[16224] <=  8'h00;      memory[16225] <=  8'h00;      memory[16226] <=  8'h00;      memory[16227] <=  8'h00;      memory[16228] <=  8'h00;      memory[16229] <=  8'h00;      memory[16230] <=  8'h00;      memory[16231] <=  8'h00;      memory[16232] <=  8'h00;      memory[16233] <=  8'h00;      memory[16234] <=  8'h00;      memory[16235] <=  8'h00;      memory[16236] <=  8'h00;      memory[16237] <=  8'h00;      memory[16238] <=  8'h00;      memory[16239] <=  8'h00;      memory[16240] <=  8'h00;      memory[16241] <=  8'h00;      memory[16242] <=  8'h00;      memory[16243] <=  8'h00;      memory[16244] <=  8'h00;      memory[16245] <=  8'h00;      memory[16246] <=  8'h00;      memory[16247] <=  8'h00;      memory[16248] <=  8'h00;      memory[16249] <=  8'h00;      memory[16250] <=  8'h00;      memory[16251] <=  8'h00;      memory[16252] <=  8'h00;      memory[16253] <=  8'h00;      memory[16254] <=  8'h00;      memory[16255] <=  8'h00;      memory[16256] <=  8'h00;      memory[16257] <=  8'h00;      memory[16258] <=  8'h00;      memory[16259] <=  8'h00;      memory[16260] <=  8'h00;      memory[16261] <=  8'h00;      memory[16262] <=  8'h00;      memory[16263] <=  8'h00;      memory[16264] <=  8'h00;      memory[16265] <=  8'h00;      memory[16266] <=  8'h00;      memory[16267] <=  8'h00;      memory[16268] <=  8'h00;      memory[16269] <=  8'h00;      memory[16270] <=  8'h00;      memory[16271] <=  8'h00;      memory[16272] <=  8'h00;      memory[16273] <=  8'h00;      memory[16274] <=  8'h00;      memory[16275] <=  8'h00;      memory[16276] <=  8'h00;      memory[16277] <=  8'h00;      memory[16278] <=  8'h00;      memory[16279] <=  8'h00;      memory[16280] <=  8'h00;      memory[16281] <=  8'h00;      memory[16282] <=  8'h00;      memory[16283] <=  8'h00;      memory[16284] <=  8'h00;      memory[16285] <=  8'h00;      memory[16286] <=  8'h00;      memory[16287] <=  8'h00;      memory[16288] <=  8'h00;      memory[16289] <=  8'h00;      memory[16290] <=  8'h00;      memory[16291] <=  8'h00;      memory[16292] <=  8'h00;      memory[16293] <=  8'h00;      memory[16294] <=  8'h00;      memory[16295] <=  8'h00;      memory[16296] <=  8'h00;      memory[16297] <=  8'h00;      memory[16298] <=  8'h00;      memory[16299] <=  8'h00;      memory[16300] <=  8'h00;      memory[16301] <=  8'h00;      memory[16302] <=  8'h00;      memory[16303] <=  8'h00;      memory[16304] <=  8'h00;      memory[16305] <=  8'h00;      memory[16306] <=  8'h00;      memory[16307] <=  8'h00;      memory[16308] <=  8'h00;      memory[16309] <=  8'h00;      memory[16310] <=  8'h00;      memory[16311] <=  8'h00;      memory[16312] <=  8'h00;      memory[16313] <=  8'h00;      memory[16314] <=  8'h00;      memory[16315] <=  8'h00;      memory[16316] <=  8'h00;      memory[16317] <=  8'h00;      memory[16318] <=  8'h00;      memory[16319] <=  8'h00;      memory[16320] <=  8'h00;      memory[16321] <=  8'h00;      memory[16322] <=  8'h00;      memory[16323] <=  8'h00;      memory[16324] <=  8'h00;      memory[16325] <=  8'h00;      memory[16326] <=  8'h00;      memory[16327] <=  8'h00;      memory[16328] <=  8'h00;      memory[16329] <=  8'h00;      memory[16330] <=  8'h00;      memory[16331] <=  8'h00;      memory[16332] <=  8'h00;      memory[16333] <=  8'h00;      memory[16334] <=  8'h00;      memory[16335] <=  8'h00;      memory[16336] <=  8'h00;      memory[16337] <=  8'h00;      memory[16338] <=  8'h00;      memory[16339] <=  8'h00;      memory[16340] <=  8'h00;      memory[16341] <=  8'h00;      memory[16342] <=  8'h00;      memory[16343] <=  8'h00;      memory[16344] <=  8'h00;      memory[16345] <=  8'h00;      memory[16346] <=  8'h00;      memory[16347] <=  8'h00;      memory[16348] <=  8'h00;      memory[16349] <=  8'h00;      memory[16350] <=  8'h00;      memory[16351] <=  8'h00;      memory[16352] <=  8'h00;      memory[16353] <=  8'h00;      memory[16354] <=  8'h00;      memory[16355] <=  8'h00;      memory[16356] <=  8'h00;      memory[16357] <=  8'h00;      memory[16358] <=  8'h00;      memory[16359] <=  8'h00;      memory[16360] <=  8'h00;      memory[16361] <=  8'h00;      memory[16362] <=  8'h00;      memory[16363] <=  8'h00;      memory[16364] <=  8'h00;      memory[16365] <=  8'h00;      memory[16366] <=  8'h00;      memory[16367] <=  8'h00;      memory[16368] <=  8'h00;      memory[16369] <=  8'h00;      memory[16370] <=  8'h00;      memory[16371] <=  8'h00;      memory[16372] <=  8'h00;      memory[16373] <=  8'h00;      memory[16374] <=  8'h00;      memory[16375] <=  8'h00;      memory[16376] <=  8'h00;      memory[16377] <=  8'h00;      memory[16378] <=  8'h00;      memory[16379] <=  8'h00;      memory[16380] <=  8'h00;      memory[16381] <=  8'h00;      memory[16382] <=  8'h00;      memory[16383] <=  8'h00;      memory[16384] <=  8'h00;      memory[16385] <=  8'h00;      memory[16386] <=  8'h00;      memory[16387] <=  8'h00;      memory[16388] <=  8'h00;      memory[16389] <=  8'h00;      memory[16390] <=  8'h00;      memory[16391] <=  8'h00;      memory[16392] <=  8'h00;      memory[16393] <=  8'h00;      memory[16394] <=  8'h00;      memory[16395] <=  8'h00;      memory[16396] <=  8'h00;      memory[16397] <=  8'h00;      memory[16398] <=  8'h00;      memory[16399] <=  8'h00;      memory[16400] <=  8'h00;      memory[16401] <=  8'h00;      memory[16402] <=  8'h00;      memory[16403] <=  8'h00;      memory[16404] <=  8'h00;      memory[16405] <=  8'h00;      memory[16406] <=  8'h00;      memory[16407] <=  8'h00;      memory[16408] <=  8'h00;      memory[16409] <=  8'h00;      memory[16410] <=  8'h00;      memory[16411] <=  8'h00;      memory[16412] <=  8'h00;      memory[16413] <=  8'h00;      memory[16414] <=  8'h00;      memory[16415] <=  8'h00;      memory[16416] <=  8'h00;      memory[16417] <=  8'h00;      memory[16418] <=  8'h00;      memory[16419] <=  8'h00;      memory[16420] <=  8'h00;      memory[16421] <=  8'h00;      memory[16422] <=  8'h00;      memory[16423] <=  8'h00;      memory[16424] <=  8'h00;      memory[16425] <=  8'h00;      memory[16426] <=  8'h00;      memory[16427] <=  8'h00;      memory[16428] <=  8'h00;      memory[16429] <=  8'h00;      memory[16430] <=  8'h00;      memory[16431] <=  8'h00;      memory[16432] <=  8'h00;      memory[16433] <=  8'h00;      memory[16434] <=  8'h00;      memory[16435] <=  8'h00;      memory[16436] <=  8'h00;      memory[16437] <=  8'h00;      memory[16438] <=  8'h00;      memory[16439] <=  8'h00;      memory[16440] <=  8'h00;      memory[16441] <=  8'h00;      memory[16442] <=  8'h00;      memory[16443] <=  8'h00;      memory[16444] <=  8'h00;      memory[16445] <=  8'h00;      memory[16446] <=  8'h00;      memory[16447] <=  8'h00;      memory[16448] <=  8'h00;      memory[16449] <=  8'h00;      memory[16450] <=  8'h00;      memory[16451] <=  8'h00;      memory[16452] <=  8'h00;      memory[16453] <=  8'h00;      memory[16454] <=  8'h00;      memory[16455] <=  8'h00;      memory[16456] <=  8'h00;      memory[16457] <=  8'h00;      memory[16458] <=  8'h00;      memory[16459] <=  8'h00;      memory[16460] <=  8'h00;      memory[16461] <=  8'h00;      memory[16462] <=  8'h00;      memory[16463] <=  8'h00;      memory[16464] <=  8'h00;      memory[16465] <=  8'h00;      memory[16466] <=  8'h00;      memory[16467] <=  8'h00;      memory[16468] <=  8'h00;      memory[16469] <=  8'h00;      memory[16470] <=  8'h00;      memory[16471] <=  8'h00;      memory[16472] <=  8'h00;      memory[16473] <=  8'h00;      memory[16474] <=  8'h00;      memory[16475] <=  8'h00;      memory[16476] <=  8'h00;      memory[16477] <=  8'h00;      memory[16478] <=  8'h00;      memory[16479] <=  8'h00;      memory[16480] <=  8'h00;      memory[16481] <=  8'h00;      memory[16482] <=  8'h00;      memory[16483] <=  8'h00;      memory[16484] <=  8'h00;      memory[16485] <=  8'h00;      memory[16486] <=  8'h00;      memory[16487] <=  8'h00;      memory[16488] <=  8'h00;      memory[16489] <=  8'h00;      memory[16490] <=  8'h00;      memory[16491] <=  8'h00;      memory[16492] <=  8'h00;      memory[16493] <=  8'h00;      memory[16494] <=  8'h00;      memory[16495] <=  8'h00;      memory[16496] <=  8'h00;      memory[16497] <=  8'h00;      memory[16498] <=  8'h00;      memory[16499] <=  8'h00;      memory[16500] <=  8'h00;      memory[16501] <=  8'h00;      memory[16502] <=  8'h00;      memory[16503] <=  8'h00;      memory[16504] <=  8'h00;      memory[16505] <=  8'h00;      memory[16506] <=  8'h00;      memory[16507] <=  8'h00;      memory[16508] <=  8'h00;      memory[16509] <=  8'h00;      memory[16510] <=  8'h00;      memory[16511] <=  8'h00;      memory[16512] <=  8'h00;      memory[16513] <=  8'h00;      memory[16514] <=  8'h00;      memory[16515] <=  8'h00;      memory[16516] <=  8'h00;      memory[16517] <=  8'h00;      memory[16518] <=  8'h00;      memory[16519] <=  8'h00;      memory[16520] <=  8'h00;      memory[16521] <=  8'h00;      memory[16522] <=  8'h00;      memory[16523] <=  8'h00;      memory[16524] <=  8'h00;      memory[16525] <=  8'h00;      memory[16526] <=  8'h00;      memory[16527] <=  8'h00;      memory[16528] <=  8'h00;      memory[16529] <=  8'h00;      memory[16530] <=  8'h00;      memory[16531] <=  8'h00;      memory[16532] <=  8'h00;      memory[16533] <=  8'h00;      memory[16534] <=  8'h00;      memory[16535] <=  8'h00;      memory[16536] <=  8'h00;      memory[16537] <=  8'h00;      memory[16538] <=  8'h00;      memory[16539] <=  8'h00;      memory[16540] <=  8'h00;      memory[16541] <=  8'h00;      memory[16542] <=  8'h00;      memory[16543] <=  8'h00;      memory[16544] <=  8'h00;      memory[16545] <=  8'h00;      memory[16546] <=  8'h00;      memory[16547] <=  8'h00;      memory[16548] <=  8'h00;      memory[16549] <=  8'h00;      memory[16550] <=  8'h00;      memory[16551] <=  8'h00;      memory[16552] <=  8'h00;      memory[16553] <=  8'h00;      memory[16554] <=  8'h00;      memory[16555] <=  8'h00;      memory[16556] <=  8'h00;      memory[16557] <=  8'h00;      memory[16558] <=  8'h00;      memory[16559] <=  8'h00;      memory[16560] <=  8'h00;      memory[16561] <=  8'h00;      memory[16562] <=  8'h00;      memory[16563] <=  8'h00;      memory[16564] <=  8'h00;      memory[16565] <=  8'h00;      memory[16566] <=  8'h00;      memory[16567] <=  8'h00;      memory[16568] <=  8'h00;      memory[16569] <=  8'h00;      memory[16570] <=  8'h00;      memory[16571] <=  8'h00;      memory[16572] <=  8'h00;      memory[16573] <=  8'h00;      memory[16574] <=  8'h00;      memory[16575] <=  8'h00;      memory[16576] <=  8'h00;      memory[16577] <=  8'h00;      memory[16578] <=  8'h00;      memory[16579] <=  8'h00;      memory[16580] <=  8'h00;      memory[16581] <=  8'h00;      memory[16582] <=  8'h00;      memory[16583] <=  8'h00;      memory[16584] <=  8'h00;      memory[16585] <=  8'h00;      memory[16586] <=  8'h00;      memory[16587] <=  8'h00;      memory[16588] <=  8'h00;      memory[16589] <=  8'h00;      memory[16590] <=  8'h00;      memory[16591] <=  8'h00;      memory[16592] <=  8'h00;      memory[16593] <=  8'h00;      memory[16594] <=  8'h00;      memory[16595] <=  8'h00;      memory[16596] <=  8'h00;      memory[16597] <=  8'h00;      memory[16598] <=  8'h00;      memory[16599] <=  8'h00;      memory[16600] <=  8'h00;      memory[16601] <=  8'h00;      memory[16602] <=  8'h00;      memory[16603] <=  8'h00;      memory[16604] <=  8'h00;      memory[16605] <=  8'h00;      memory[16606] <=  8'h00;      memory[16607] <=  8'h00;      memory[16608] <=  8'h00;      memory[16609] <=  8'h00;      memory[16610] <=  8'h00;      memory[16611] <=  8'h00;      memory[16612] <=  8'h00;      memory[16613] <=  8'h00;      memory[16614] <=  8'h00;      memory[16615] <=  8'h00;      memory[16616] <=  8'h00;      memory[16617] <=  8'h00;      memory[16618] <=  8'h00;      memory[16619] <=  8'h00;      memory[16620] <=  8'h00;      memory[16621] <=  8'h00;      memory[16622] <=  8'h00;      memory[16623] <=  8'h00;      memory[16624] <=  8'h00;      memory[16625] <=  8'h00;      memory[16626] <=  8'h00;      memory[16627] <=  8'h00;      memory[16628] <=  8'h00;      memory[16629] <=  8'h00;      memory[16630] <=  8'h00;      memory[16631] <=  8'h00;      memory[16632] <=  8'h00;      memory[16633] <=  8'h00;      memory[16634] <=  8'h00;      memory[16635] <=  8'h00;      memory[16636] <=  8'h00;      memory[16637] <=  8'h00;      memory[16638] <=  8'h00;      memory[16639] <=  8'h00;      memory[16640] <=  8'h00;      memory[16641] <=  8'h00;      memory[16642] <=  8'h00;      memory[16643] <=  8'h00;      memory[16644] <=  8'h00;      memory[16645] <=  8'h00;      memory[16646] <=  8'h00;      memory[16647] <=  8'h00;      memory[16648] <=  8'h00;      memory[16649] <=  8'h00;      memory[16650] <=  8'h00;      memory[16651] <=  8'h00;      memory[16652] <=  8'h00;      memory[16653] <=  8'h00;      memory[16654] <=  8'h00;      memory[16655] <=  8'h00;      memory[16656] <=  8'h00;      memory[16657] <=  8'h00;      memory[16658] <=  8'h00;      memory[16659] <=  8'h00;      memory[16660] <=  8'h00;      memory[16661] <=  8'h00;      memory[16662] <=  8'h00;      memory[16663] <=  8'h00;      memory[16664] <=  8'h00;      memory[16665] <=  8'h00;      memory[16666] <=  8'h00;      memory[16667] <=  8'h00;      memory[16668] <=  8'h00;      memory[16669] <=  8'h00;      memory[16670] <=  8'h00;      memory[16671] <=  8'h00;      memory[16672] <=  8'h00;      memory[16673] <=  8'h00;      memory[16674] <=  8'h00;      memory[16675] <=  8'h00;      memory[16676] <=  8'h00;      memory[16677] <=  8'h00;      memory[16678] <=  8'h00;      memory[16679] <=  8'h00;      memory[16680] <=  8'h00;      memory[16681] <=  8'h00;      memory[16682] <=  8'h00;      memory[16683] <=  8'h00;      memory[16684] <=  8'h00;      memory[16685] <=  8'h00;      memory[16686] <=  8'h00;      memory[16687] <=  8'h00;      memory[16688] <=  8'h00;      memory[16689] <=  8'h00;      memory[16690] <=  8'h00;      memory[16691] <=  8'h00;      memory[16692] <=  8'h00;      memory[16693] <=  8'h00;      memory[16694] <=  8'h00;      memory[16695] <=  8'h00;      memory[16696] <=  8'h00;      memory[16697] <=  8'h00;      memory[16698] <=  8'h00;      memory[16699] <=  8'h00;      memory[16700] <=  8'h00;      memory[16701] <=  8'h00;      memory[16702] <=  8'h00;      memory[16703] <=  8'h00;      memory[16704] <=  8'h00;      memory[16705] <=  8'h00;      memory[16706] <=  8'h00;      memory[16707] <=  8'h00;      memory[16708] <=  8'h00;      memory[16709] <=  8'h00;      memory[16710] <=  8'h00;      memory[16711] <=  8'h00;      memory[16712] <=  8'h00;      memory[16713] <=  8'h00;      memory[16714] <=  8'h00;      memory[16715] <=  8'h00;      memory[16716] <=  8'h00;      memory[16717] <=  8'h00;      memory[16718] <=  8'h00;      memory[16719] <=  8'h00;      memory[16720] <=  8'h00;      memory[16721] <=  8'h00;      memory[16722] <=  8'h00;      memory[16723] <=  8'h00;      memory[16724] <=  8'h00;      memory[16725] <=  8'h00;      memory[16726] <=  8'h00;      memory[16727] <=  8'h00;      memory[16728] <=  8'h00;      memory[16729] <=  8'h00;      memory[16730] <=  8'h00;      memory[16731] <=  8'h00;      memory[16732] <=  8'h00;      memory[16733] <=  8'h00;      memory[16734] <=  8'h00;      memory[16735] <=  8'h00;      memory[16736] <=  8'h00;      memory[16737] <=  8'h00;      memory[16738] <=  8'h00;      memory[16739] <=  8'h00;      memory[16740] <=  8'h00;      memory[16741] <=  8'h00;      memory[16742] <=  8'h00;      memory[16743] <=  8'h00;      memory[16744] <=  8'h00;      memory[16745] <=  8'h00;      memory[16746] <=  8'h00;      memory[16747] <=  8'h00;      memory[16748] <=  8'h00;      memory[16749] <=  8'h00;      memory[16750] <=  8'h00;      memory[16751] <=  8'h00;      memory[16752] <=  8'h00;      memory[16753] <=  8'h00;      memory[16754] <=  8'h00;      memory[16755] <=  8'h00;      memory[16756] <=  8'h00;      memory[16757] <=  8'h00;      memory[16758] <=  8'h00;      memory[16759] <=  8'h00;      memory[16760] <=  8'h00;      memory[16761] <=  8'h00;      memory[16762] <=  8'h00;      memory[16763] <=  8'h00;      memory[16764] <=  8'h00;      memory[16765] <=  8'h00;      memory[16766] <=  8'h00;      memory[16767] <=  8'h00;      memory[16768] <=  8'h00;      memory[16769] <=  8'h00;      memory[16770] <=  8'h00;      memory[16771] <=  8'h00;      memory[16772] <=  8'h00;      memory[16773] <=  8'h00;      memory[16774] <=  8'h00;      memory[16775] <=  8'h00;      memory[16776] <=  8'h00;      memory[16777] <=  8'h00;      memory[16778] <=  8'h00;      memory[16779] <=  8'h00;      memory[16780] <=  8'h00;      memory[16781] <=  8'h00;      memory[16782] <=  8'h00;      memory[16783] <=  8'h00;      memory[16784] <=  8'h00;      memory[16785] <=  8'h00;      memory[16786] <=  8'h00;      memory[16787] <=  8'h00;      memory[16788] <=  8'h00;      memory[16789] <=  8'h00;      memory[16790] <=  8'h00;      memory[16791] <=  8'h00;      memory[16792] <=  8'h00;      memory[16793] <=  8'h00;      memory[16794] <=  8'h00;      memory[16795] <=  8'h00;      memory[16796] <=  8'h00;      memory[16797] <=  8'h00;      memory[16798] <=  8'h00;      memory[16799] <=  8'h00;      memory[16800] <=  8'h00;      memory[16801] <=  8'h00;      memory[16802] <=  8'h00;      memory[16803] <=  8'h00;      memory[16804] <=  8'h00;      memory[16805] <=  8'h00;      memory[16806] <=  8'h00;      memory[16807] <=  8'h00;      memory[16808] <=  8'h00;      memory[16809] <=  8'h00;      memory[16810] <=  8'h00;      memory[16811] <=  8'h00;      memory[16812] <=  8'h00;      memory[16813] <=  8'h00;      memory[16814] <=  8'h00;      memory[16815] <=  8'h00;      memory[16816] <=  8'h00;      memory[16817] <=  8'h00;      memory[16818] <=  8'h00;      memory[16819] <=  8'h00;      memory[16820] <=  8'h00;      memory[16821] <=  8'h00;      memory[16822] <=  8'h00;      memory[16823] <=  8'h00;      memory[16824] <=  8'h00;      memory[16825] <=  8'h00;      memory[16826] <=  8'h00;      memory[16827] <=  8'h00;      memory[16828] <=  8'h00;      memory[16829] <=  8'h00;      memory[16830] <=  8'h00;      memory[16831] <=  8'h00;      memory[16832] <=  8'h00;      memory[16833] <=  8'h00;      memory[16834] <=  8'h00;      memory[16835] <=  8'h00;      memory[16836] <=  8'h00;      memory[16837] <=  8'h00;      memory[16838] <=  8'h00;      memory[16839] <=  8'h00;      memory[16840] <=  8'h00;      memory[16841] <=  8'h00;      memory[16842] <=  8'h00;      memory[16843] <=  8'h00;      memory[16844] <=  8'h00;      memory[16845] <=  8'h00;      memory[16846] <=  8'h00;      memory[16847] <=  8'h00;      memory[16848] <=  8'h00;      memory[16849] <=  8'h00;      memory[16850] <=  8'h00;      memory[16851] <=  8'h00;      memory[16852] <=  8'h00;      memory[16853] <=  8'h00;      memory[16854] <=  8'h00;      memory[16855] <=  8'h00;      memory[16856] <=  8'h00;      memory[16857] <=  8'h00;      memory[16858] <=  8'h00;      memory[16859] <=  8'h00;      memory[16860] <=  8'h00;      memory[16861] <=  8'h00;      memory[16862] <=  8'h00;      memory[16863] <=  8'h00;      memory[16864] <=  8'h00;      memory[16865] <=  8'h00;      memory[16866] <=  8'h00;      memory[16867] <=  8'h00;      memory[16868] <=  8'h00;      memory[16869] <=  8'h00;      memory[16870] <=  8'h00;      memory[16871] <=  8'h00;      memory[16872] <=  8'h00;      memory[16873] <=  8'h00;      memory[16874] <=  8'h00;      memory[16875] <=  8'h00;      memory[16876] <=  8'h00;      memory[16877] <=  8'h00;      memory[16878] <=  8'h00;      memory[16879] <=  8'h00;      memory[16880] <=  8'h00;      memory[16881] <=  8'h00;      memory[16882] <=  8'h00;      memory[16883] <=  8'h00;      memory[16884] <=  8'h00;      memory[16885] <=  8'h00;      memory[16886] <=  8'h00;      memory[16887] <=  8'h00;      memory[16888] <=  8'h00;      memory[16889] <=  8'h00;      memory[16890] <=  8'h00;      memory[16891] <=  8'h00;      memory[16892] <=  8'h00;      memory[16893] <=  8'h00;      memory[16894] <=  8'h00;      memory[16895] <=  8'h00;      memory[16896] <=  8'h00;      memory[16897] <=  8'h00;      memory[16898] <=  8'h00;      memory[16899] <=  8'h00;      memory[16900] <=  8'h00;      memory[16901] <=  8'h00;      memory[16902] <=  8'h00;      memory[16903] <=  8'h00;      memory[16904] <=  8'h00;      memory[16905] <=  8'h00;      memory[16906] <=  8'h00;      memory[16907] <=  8'h00;      memory[16908] <=  8'h00;      memory[16909] <=  8'h00;      memory[16910] <=  8'h00;      memory[16911] <=  8'h00;      memory[16912] <=  8'h00;      memory[16913] <=  8'h00;      memory[16914] <=  8'h00;      memory[16915] <=  8'h00;      memory[16916] <=  8'h00;      memory[16917] <=  8'h00;      memory[16918] <=  8'h00;      memory[16919] <=  8'h00;      memory[16920] <=  8'h00;      memory[16921] <=  8'h00;      memory[16922] <=  8'h00;      memory[16923] <=  8'h00;      memory[16924] <=  8'h00;      memory[16925] <=  8'h00;      memory[16926] <=  8'h00;      memory[16927] <=  8'h00;      memory[16928] <=  8'h00;      memory[16929] <=  8'h00;      memory[16930] <=  8'h00;      memory[16931] <=  8'h00;      memory[16932] <=  8'h00;      memory[16933] <=  8'h00;      memory[16934] <=  8'h00;      memory[16935] <=  8'h00;      memory[16936] <=  8'h00;      memory[16937] <=  8'h00;      memory[16938] <=  8'h00;      memory[16939] <=  8'h00;      memory[16940] <=  8'h00;      memory[16941] <=  8'h00;      memory[16942] <=  8'h00;      memory[16943] <=  8'h00;      memory[16944] <=  8'h00;      memory[16945] <=  8'h00;      memory[16946] <=  8'h00;      memory[16947] <=  8'h00;      memory[16948] <=  8'h00;      memory[16949] <=  8'h00;      memory[16950] <=  8'h00;      memory[16951] <=  8'h00;      memory[16952] <=  8'h00;      memory[16953] <=  8'h00;      memory[16954] <=  8'h00;      memory[16955] <=  8'h00;      memory[16956] <=  8'h00;      memory[16957] <=  8'h00;      memory[16958] <=  8'h00;      memory[16959] <=  8'h00;      memory[16960] <=  8'h00;      memory[16961] <=  8'h00;      memory[16962] <=  8'h00;      memory[16963] <=  8'h00;      memory[16964] <=  8'h00;      memory[16965] <=  8'h00;      memory[16966] <=  8'h00;      memory[16967] <=  8'h00;      memory[16968] <=  8'h00;      memory[16969] <=  8'h00;      memory[16970] <=  8'h00;      memory[16971] <=  8'h00;      memory[16972] <=  8'h00;      memory[16973] <=  8'h00;      memory[16974] <=  8'h00;      memory[16975] <=  8'h00;      memory[16976] <=  8'h00;      memory[16977] <=  8'h00;      memory[16978] <=  8'h00;      memory[16979] <=  8'h00;      memory[16980] <=  8'h00;      memory[16981] <=  8'h00;      memory[16982] <=  8'h00;      memory[16983] <=  8'h00;      memory[16984] <=  8'h00;      memory[16985] <=  8'h00;      memory[16986] <=  8'h00;      memory[16987] <=  8'h00;      memory[16988] <=  8'h00;      memory[16989] <=  8'h00;      memory[16990] <=  8'h00;      memory[16991] <=  8'h00;      memory[16992] <=  8'h00;      memory[16993] <=  8'h00;      memory[16994] <=  8'h00;      memory[16995] <=  8'h00;      memory[16996] <=  8'h00;      memory[16997] <=  8'h00;      memory[16998] <=  8'h00;      memory[16999] <=  8'h00;      memory[17000] <=  8'h00;      memory[17001] <=  8'h00;      memory[17002] <=  8'h00;      memory[17003] <=  8'h00;      memory[17004] <=  8'h00;      memory[17005] <=  8'h00;      memory[17006] <=  8'h00;      memory[17007] <=  8'h00;      memory[17008] <=  8'h00;      memory[17009] <=  8'h00;      memory[17010] <=  8'h00;      memory[17011] <=  8'h00;      memory[17012] <=  8'h00;      memory[17013] <=  8'h00;      memory[17014] <=  8'h00;      memory[17015] <=  8'h00;      memory[17016] <=  8'h00;      memory[17017] <=  8'h00;      memory[17018] <=  8'h00;      memory[17019] <=  8'h00;      memory[17020] <=  8'h00;      memory[17021] <=  8'h00;      memory[17022] <=  8'h00;      memory[17023] <=  8'h00;      memory[17024] <=  8'h00;      memory[17025] <=  8'h00;      memory[17026] <=  8'h00;      memory[17027] <=  8'h00;      memory[17028] <=  8'h00;      memory[17029] <=  8'h00;      memory[17030] <=  8'h00;      memory[17031] <=  8'h00;      memory[17032] <=  8'h00;      memory[17033] <=  8'h00;      memory[17034] <=  8'h00;      memory[17035] <=  8'h00;      memory[17036] <=  8'h00;      memory[17037] <=  8'h00;      memory[17038] <=  8'h00;      memory[17039] <=  8'h00;      memory[17040] <=  8'h00;      memory[17041] <=  8'h00;      memory[17042] <=  8'h00;      memory[17043] <=  8'h00;      memory[17044] <=  8'h00;      memory[17045] <=  8'h00;      memory[17046] <=  8'h00;      memory[17047] <=  8'h00;      memory[17048] <=  8'h00;      memory[17049] <=  8'h00;      memory[17050] <=  8'h00;      memory[17051] <=  8'h00;      memory[17052] <=  8'h00;      memory[17053] <=  8'h00;      memory[17054] <=  8'h00;      memory[17055] <=  8'h00;      memory[17056] <=  8'h00;      memory[17057] <=  8'h00;      memory[17058] <=  8'h00;      memory[17059] <=  8'h00;      memory[17060] <=  8'h00;      memory[17061] <=  8'h00;      memory[17062] <=  8'h00;      memory[17063] <=  8'h00;      memory[17064] <=  8'h00;      memory[17065] <=  8'h00;      memory[17066] <=  8'h00;      memory[17067] <=  8'h00;      memory[17068] <=  8'h00;      memory[17069] <=  8'h00;      memory[17070] <=  8'h00;      memory[17071] <=  8'h00;      memory[17072] <=  8'h00;      memory[17073] <=  8'h00;      memory[17074] <=  8'h00;      memory[17075] <=  8'h00;      memory[17076] <=  8'h00;      memory[17077] <=  8'h00;      memory[17078] <=  8'h00;      memory[17079] <=  8'h00;      memory[17080] <=  8'h00;      memory[17081] <=  8'h00;      memory[17082] <=  8'h00;      memory[17083] <=  8'h00;      memory[17084] <=  8'h00;      memory[17085] <=  8'h00;      memory[17086] <=  8'h00;      memory[17087] <=  8'h00;      memory[17088] <=  8'h00;      memory[17089] <=  8'h00;      memory[17090] <=  8'h00;      memory[17091] <=  8'h00;      memory[17092] <=  8'h00;      memory[17093] <=  8'h00;      memory[17094] <=  8'h00;      memory[17095] <=  8'h00;      memory[17096] <=  8'h00;      memory[17097] <=  8'h00;      memory[17098] <=  8'h00;      memory[17099] <=  8'h00;      memory[17100] <=  8'h00;      memory[17101] <=  8'h00;      memory[17102] <=  8'h00;      memory[17103] <=  8'h00;      memory[17104] <=  8'h00;      memory[17105] <=  8'h00;      memory[17106] <=  8'h00;      memory[17107] <=  8'h00;      memory[17108] <=  8'h00;      memory[17109] <=  8'h00;      memory[17110] <=  8'h00;      memory[17111] <=  8'h00;      memory[17112] <=  8'h00;      memory[17113] <=  8'h00;      memory[17114] <=  8'h00;      memory[17115] <=  8'h00;      memory[17116] <=  8'h00;      memory[17117] <=  8'h00;      memory[17118] <=  8'h00;      memory[17119] <=  8'h00;      memory[17120] <=  8'h00;      memory[17121] <=  8'h00;      memory[17122] <=  8'h00;      memory[17123] <=  8'h00;      memory[17124] <=  8'h00;      memory[17125] <=  8'h00;      memory[17126] <=  8'h00;      memory[17127] <=  8'h00;      memory[17128] <=  8'h00;      memory[17129] <=  8'h00;      memory[17130] <=  8'h00;      memory[17131] <=  8'h00;      memory[17132] <=  8'h00;      memory[17133] <=  8'h00;      memory[17134] <=  8'h00;      memory[17135] <=  8'h00;      memory[17136] <=  8'h00;      memory[17137] <=  8'h00;      memory[17138] <=  8'h00;      memory[17139] <=  8'h00;      memory[17140] <=  8'h00;      memory[17141] <=  8'h00;      memory[17142] <=  8'h00;      memory[17143] <=  8'h00;      memory[17144] <=  8'h00;      memory[17145] <=  8'h00;      memory[17146] <=  8'h00;      memory[17147] <=  8'h00;      memory[17148] <=  8'h00;      memory[17149] <=  8'h00;      memory[17150] <=  8'h00;      memory[17151] <=  8'h00;      memory[17152] <=  8'h00;      memory[17153] <=  8'h00;      memory[17154] <=  8'h00;      memory[17155] <=  8'h00;      memory[17156] <=  8'h00;      memory[17157] <=  8'h00;      memory[17158] <=  8'h00;      memory[17159] <=  8'h00;      memory[17160] <=  8'h00;      memory[17161] <=  8'h00;      memory[17162] <=  8'h00;      memory[17163] <=  8'h00;      memory[17164] <=  8'h00;      memory[17165] <=  8'h00;      memory[17166] <=  8'h00;      memory[17167] <=  8'h00;      memory[17168] <=  8'h00;      memory[17169] <=  8'h00;      memory[17170] <=  8'h00;      memory[17171] <=  8'h00;      memory[17172] <=  8'h00;      memory[17173] <=  8'h00;      memory[17174] <=  8'h00;      memory[17175] <=  8'h00;      memory[17176] <=  8'h00;      memory[17177] <=  8'h00;      memory[17178] <=  8'h00;      memory[17179] <=  8'h00;      memory[17180] <=  8'h00;      memory[17181] <=  8'h00;      memory[17182] <=  8'h00;      memory[17183] <=  8'h00;      memory[17184] <=  8'h00;      memory[17185] <=  8'h00;      memory[17186] <=  8'h00;      memory[17187] <=  8'h00;      memory[17188] <=  8'h00;      memory[17189] <=  8'h00;      memory[17190] <=  8'h00;      memory[17191] <=  8'h00;      memory[17192] <=  8'h00;      memory[17193] <=  8'h00;      memory[17194] <=  8'h00;      memory[17195] <=  8'h00;      memory[17196] <=  8'h00;      memory[17197] <=  8'h00;      memory[17198] <=  8'h00;      memory[17199] <=  8'h00;      memory[17200] <=  8'h00;      memory[17201] <=  8'h00;      memory[17202] <=  8'h00;      memory[17203] <=  8'h00;      memory[17204] <=  8'h00;      memory[17205] <=  8'h00;      memory[17206] <=  8'h00;      memory[17207] <=  8'h00;      memory[17208] <=  8'h00;      memory[17209] <=  8'h00;      memory[17210] <=  8'h00;      memory[17211] <=  8'h00;      memory[17212] <=  8'h00;      memory[17213] <=  8'h00;      memory[17214] <=  8'h00;      memory[17215] <=  8'h00;      memory[17216] <=  8'h00;      memory[17217] <=  8'h00;      memory[17218] <=  8'h00;      memory[17219] <=  8'h00;      memory[17220] <=  8'h00;      memory[17221] <=  8'h00;      memory[17222] <=  8'h00;      memory[17223] <=  8'h00;      memory[17224] <=  8'h00;      memory[17225] <=  8'h00;      memory[17226] <=  8'h00;      memory[17227] <=  8'h00;      memory[17228] <=  8'h00;      memory[17229] <=  8'h00;      memory[17230] <=  8'h00;      memory[17231] <=  8'h00;      memory[17232] <=  8'h00;      memory[17233] <=  8'h00;      memory[17234] <=  8'h00;      memory[17235] <=  8'h00;      memory[17236] <=  8'h00;      memory[17237] <=  8'h00;      memory[17238] <=  8'h00;      memory[17239] <=  8'h00;      memory[17240] <=  8'h00;      memory[17241] <=  8'h00;      memory[17242] <=  8'h00;      memory[17243] <=  8'h00;      memory[17244] <=  8'h00;      memory[17245] <=  8'h00;      memory[17246] <=  8'h00;      memory[17247] <=  8'h00;      memory[17248] <=  8'h00;      memory[17249] <=  8'h00;      memory[17250] <=  8'h00;      memory[17251] <=  8'h00;      memory[17252] <=  8'h00;      memory[17253] <=  8'h00;      memory[17254] <=  8'h00;      memory[17255] <=  8'h00;      memory[17256] <=  8'h00;      memory[17257] <=  8'h00;      memory[17258] <=  8'h00;      memory[17259] <=  8'h00;      memory[17260] <=  8'h00;      memory[17261] <=  8'h00;      memory[17262] <=  8'h00;      memory[17263] <=  8'h00;      memory[17264] <=  8'h00;      memory[17265] <=  8'h00;      memory[17266] <=  8'h00;      memory[17267] <=  8'h00;      memory[17268] <=  8'h00;      memory[17269] <=  8'h00;      memory[17270] <=  8'h00;      memory[17271] <=  8'h00;      memory[17272] <=  8'h00;      memory[17273] <=  8'h00;      memory[17274] <=  8'h00;      memory[17275] <=  8'h00;      memory[17276] <=  8'h00;      memory[17277] <=  8'h00;      memory[17278] <=  8'h00;      memory[17279] <=  8'h00;      memory[17280] <=  8'h00;      memory[17281] <=  8'h00;      memory[17282] <=  8'h00;      memory[17283] <=  8'h00;      memory[17284] <=  8'h00;      memory[17285] <=  8'h00;      memory[17286] <=  8'h00;      memory[17287] <=  8'h00;      memory[17288] <=  8'h00;      memory[17289] <=  8'h00;      memory[17290] <=  8'h00;      memory[17291] <=  8'h00;      memory[17292] <=  8'h00;      memory[17293] <=  8'h00;      memory[17294] <=  8'h00;      memory[17295] <=  8'h00;      memory[17296] <=  8'h00;      memory[17297] <=  8'h00;      memory[17298] <=  8'h00;      memory[17299] <=  8'h00;      memory[17300] <=  8'h00;      memory[17301] <=  8'h00;      memory[17302] <=  8'h00;      memory[17303] <=  8'h00;      memory[17304] <=  8'h00;      memory[17305] <=  8'h00;      memory[17306] <=  8'h00;      memory[17307] <=  8'h00;      memory[17308] <=  8'h00;      memory[17309] <=  8'h00;      memory[17310] <=  8'h00;      memory[17311] <=  8'h00;      memory[17312] <=  8'h00;      memory[17313] <=  8'h00;      memory[17314] <=  8'h00;      memory[17315] <=  8'h00;      memory[17316] <=  8'h00;      memory[17317] <=  8'h00;      memory[17318] <=  8'h00;      memory[17319] <=  8'h00;      memory[17320] <=  8'h00;      memory[17321] <=  8'h00;      memory[17322] <=  8'h00;      memory[17323] <=  8'h00;      memory[17324] <=  8'h00;      memory[17325] <=  8'h00;      memory[17326] <=  8'h00;      memory[17327] <=  8'h00;      memory[17328] <=  8'h00;      memory[17329] <=  8'h00;      memory[17330] <=  8'h00;      memory[17331] <=  8'h00;      memory[17332] <=  8'h00;      memory[17333] <=  8'h00;      memory[17334] <=  8'h00;      memory[17335] <=  8'h00;      memory[17336] <=  8'h00;      memory[17337] <=  8'h00;      memory[17338] <=  8'h00;      memory[17339] <=  8'h00;      memory[17340] <=  8'h00;      memory[17341] <=  8'h00;      memory[17342] <=  8'h00;      memory[17343] <=  8'h00;      memory[17344] <=  8'h00;      memory[17345] <=  8'h00;      memory[17346] <=  8'h00;      memory[17347] <=  8'h00;      memory[17348] <=  8'h00;      memory[17349] <=  8'h00;      memory[17350] <=  8'h00;      memory[17351] <=  8'h00;      memory[17352] <=  8'h00;      memory[17353] <=  8'h00;      memory[17354] <=  8'h00;      memory[17355] <=  8'h00;      memory[17356] <=  8'h00;      memory[17357] <=  8'h00;      memory[17358] <=  8'h00;      memory[17359] <=  8'h00;      memory[17360] <=  8'h00;      memory[17361] <=  8'h00;      memory[17362] <=  8'h00;      memory[17363] <=  8'h00;      memory[17364] <=  8'h00;      memory[17365] <=  8'h00;      memory[17366] <=  8'h00;      memory[17367] <=  8'h00;      memory[17368] <=  8'h00;      memory[17369] <=  8'h00;      memory[17370] <=  8'h00;      memory[17371] <=  8'h00;      memory[17372] <=  8'h00;      memory[17373] <=  8'h00;      memory[17374] <=  8'h00;      memory[17375] <=  8'h00;      memory[17376] <=  8'h00;      memory[17377] <=  8'h00;      memory[17378] <=  8'h00;      memory[17379] <=  8'h00;      memory[17380] <=  8'h00;      memory[17381] <=  8'h00;      memory[17382] <=  8'h00;      memory[17383] <=  8'h00;      memory[17384] <=  8'h00;      memory[17385] <=  8'h00;      memory[17386] <=  8'h00;      memory[17387] <=  8'h00;      memory[17388] <=  8'h00;      memory[17389] <=  8'h00;      memory[17390] <=  8'h00;      memory[17391] <=  8'h00;      memory[17392] <=  8'h00;      memory[17393] <=  8'h00;      memory[17394] <=  8'h00;      memory[17395] <=  8'h00;      memory[17396] <=  8'h00;      memory[17397] <=  8'h00;      memory[17398] <=  8'h00;      memory[17399] <=  8'h00;      memory[17400] <=  8'h00;      memory[17401] <=  8'h00;      memory[17402] <=  8'h00;      memory[17403] <=  8'h00;      memory[17404] <=  8'h00;      memory[17405] <=  8'h00;      memory[17406] <=  8'h00;      memory[17407] <=  8'h00;      memory[17408] <=  8'h00;      memory[17409] <=  8'h00;      memory[17410] <=  8'h00;      memory[17411] <=  8'h00;      memory[17412] <=  8'h00;      memory[17413] <=  8'h00;      memory[17414] <=  8'h00;      memory[17415] <=  8'h00;      memory[17416] <=  8'h00;      memory[17417] <=  8'h00;      memory[17418] <=  8'h00;      memory[17419] <=  8'h00;      memory[17420] <=  8'h00;      memory[17421] <=  8'h00;      memory[17422] <=  8'h00;      memory[17423] <=  8'h00;      memory[17424] <=  8'h00;      memory[17425] <=  8'h00;      memory[17426] <=  8'h00;      memory[17427] <=  8'h00;      memory[17428] <=  8'h00;      memory[17429] <=  8'h00;      memory[17430] <=  8'h00;      memory[17431] <=  8'h00;      memory[17432] <=  8'h00;      memory[17433] <=  8'h00;      memory[17434] <=  8'h00;      memory[17435] <=  8'h00;      memory[17436] <=  8'h00;      memory[17437] <=  8'h00;      memory[17438] <=  8'h00;      memory[17439] <=  8'h00;      memory[17440] <=  8'h00;      memory[17441] <=  8'h00;      memory[17442] <=  8'h00;      memory[17443] <=  8'h00;      memory[17444] <=  8'h00;      memory[17445] <=  8'h00;      memory[17446] <=  8'h00;      memory[17447] <=  8'h00;      memory[17448] <=  8'h00;      memory[17449] <=  8'h00;      memory[17450] <=  8'h00;      memory[17451] <=  8'h00;      memory[17452] <=  8'h00;      memory[17453] <=  8'h00;      memory[17454] <=  8'h00;      memory[17455] <=  8'h00;      memory[17456] <=  8'h00;      memory[17457] <=  8'h00;      memory[17458] <=  8'h00;      memory[17459] <=  8'h00;      memory[17460] <=  8'h00;      memory[17461] <=  8'h00;      memory[17462] <=  8'h00;      memory[17463] <=  8'h00;      memory[17464] <=  8'h00;      memory[17465] <=  8'h00;      memory[17466] <=  8'h00;      memory[17467] <=  8'h00;      memory[17468] <=  8'h00;      memory[17469] <=  8'h00;      memory[17470] <=  8'h00;      memory[17471] <=  8'h00;      memory[17472] <=  8'h00;      memory[17473] <=  8'h00;      memory[17474] <=  8'h00;      memory[17475] <=  8'h00;      memory[17476] <=  8'h00;      memory[17477] <=  8'h00;      memory[17478] <=  8'h00;      memory[17479] <=  8'h00;      memory[17480] <=  8'h00;      memory[17481] <=  8'h00;      memory[17482] <=  8'h00;      memory[17483] <=  8'h00;      memory[17484] <=  8'h00;      memory[17485] <=  8'h00;      memory[17486] <=  8'h00;      memory[17487] <=  8'h00;      memory[17488] <=  8'h00;      memory[17489] <=  8'h00;      memory[17490] <=  8'h00;      memory[17491] <=  8'h00;      memory[17492] <=  8'h00;      memory[17493] <=  8'h00;      memory[17494] <=  8'h00;      memory[17495] <=  8'h00;      memory[17496] <=  8'h00;      memory[17497] <=  8'h00;      memory[17498] <=  8'h00;      memory[17499] <=  8'h00;      memory[17500] <=  8'h00;      memory[17501] <=  8'h00;      memory[17502] <=  8'h00;      memory[17503] <=  8'h00;      memory[17504] <=  8'h00;      memory[17505] <=  8'h00;      memory[17506] <=  8'h00;      memory[17507] <=  8'h00;      memory[17508] <=  8'h00;      memory[17509] <=  8'h00;      memory[17510] <=  8'h00;      memory[17511] <=  8'h00;      memory[17512] <=  8'h00;      memory[17513] <=  8'h00;      memory[17514] <=  8'h00;      memory[17515] <=  8'h00;      memory[17516] <=  8'h00;      memory[17517] <=  8'h00;      memory[17518] <=  8'h00;      memory[17519] <=  8'h00;      memory[17520] <=  8'h00;      memory[17521] <=  8'h00;      memory[17522] <=  8'h00;      memory[17523] <=  8'h00;      memory[17524] <=  8'h00;      memory[17525] <=  8'h00;      memory[17526] <=  8'h00;      memory[17527] <=  8'h00;      memory[17528] <=  8'h00;      memory[17529] <=  8'h00;      memory[17530] <=  8'h00;      memory[17531] <=  8'h00;      memory[17532] <=  8'h00;      memory[17533] <=  8'h00;      memory[17534] <=  8'h00;      memory[17535] <=  8'h00;      memory[17536] <=  8'h00;      memory[17537] <=  8'h00;      memory[17538] <=  8'h00;      memory[17539] <=  8'h00;      memory[17540] <=  8'h00;      memory[17541] <=  8'h00;      memory[17542] <=  8'h00;      memory[17543] <=  8'h00;      memory[17544] <=  8'h00;      memory[17545] <=  8'h00;      memory[17546] <=  8'h00;      memory[17547] <=  8'h00;      memory[17548] <=  8'h00;      memory[17549] <=  8'h00;      memory[17550] <=  8'h00;      memory[17551] <=  8'h00;      memory[17552] <=  8'h00;      memory[17553] <=  8'h00;      memory[17554] <=  8'h00;      memory[17555] <=  8'h00;      memory[17556] <=  8'h00;      memory[17557] <=  8'h00;      memory[17558] <=  8'h00;      memory[17559] <=  8'h00;      memory[17560] <=  8'h00;      memory[17561] <=  8'h00;      memory[17562] <=  8'h00;      memory[17563] <=  8'h00;      memory[17564] <=  8'h00;      memory[17565] <=  8'h00;      memory[17566] <=  8'h00;      memory[17567] <=  8'h00;      memory[17568] <=  8'h00;      memory[17569] <=  8'h00;      memory[17570] <=  8'h00;      memory[17571] <=  8'h00;      memory[17572] <=  8'h00;      memory[17573] <=  8'h00;      memory[17574] <=  8'h00;      memory[17575] <=  8'h00;      memory[17576] <=  8'h00;      memory[17577] <=  8'h00;      memory[17578] <=  8'h00;      memory[17579] <=  8'h00;      memory[17580] <=  8'h00;      memory[17581] <=  8'h00;      memory[17582] <=  8'h00;      memory[17583] <=  8'h00;      memory[17584] <=  8'h00;      memory[17585] <=  8'h00;      memory[17586] <=  8'h00;      memory[17587] <=  8'h00;      memory[17588] <=  8'h00;      memory[17589] <=  8'h00;      memory[17590] <=  8'h00;      memory[17591] <=  8'h00;      memory[17592] <=  8'h00;      memory[17593] <=  8'h00;      memory[17594] <=  8'h00;      memory[17595] <=  8'h00;      memory[17596] <=  8'h00;      memory[17597] <=  8'h00;      memory[17598] <=  8'h00;      memory[17599] <=  8'h00;      memory[17600] <=  8'h00;      memory[17601] <=  8'h00;      memory[17602] <=  8'h00;      memory[17603] <=  8'h00;      memory[17604] <=  8'h00;      memory[17605] <=  8'h00;      memory[17606] <=  8'h00;      memory[17607] <=  8'h00;      memory[17608] <=  8'h00;      memory[17609] <=  8'h00;      memory[17610] <=  8'h00;      memory[17611] <=  8'h00;      memory[17612] <=  8'h00;      memory[17613] <=  8'h00;      memory[17614] <=  8'h00;      memory[17615] <=  8'h00;      memory[17616] <=  8'h00;      memory[17617] <=  8'h00;      memory[17618] <=  8'h00;      memory[17619] <=  8'h00;      memory[17620] <=  8'h00;      memory[17621] <=  8'h00;      memory[17622] <=  8'h00;      memory[17623] <=  8'h00;      memory[17624] <=  8'h00;      memory[17625] <=  8'h00;      memory[17626] <=  8'h00;      memory[17627] <=  8'h00;      memory[17628] <=  8'h00;      memory[17629] <=  8'h00;      memory[17630] <=  8'h00;      memory[17631] <=  8'h00;      memory[17632] <=  8'h00;      memory[17633] <=  8'h00;      memory[17634] <=  8'h00;      memory[17635] <=  8'h00;      memory[17636] <=  8'h00;      memory[17637] <=  8'h00;      memory[17638] <=  8'h00;      memory[17639] <=  8'h00;      memory[17640] <=  8'h00;      memory[17641] <=  8'h00;      memory[17642] <=  8'h00;      memory[17643] <=  8'h00;      memory[17644] <=  8'h00;      memory[17645] <=  8'h00;      memory[17646] <=  8'h00;      memory[17647] <=  8'h00;      memory[17648] <=  8'h00;      memory[17649] <=  8'h00;      memory[17650] <=  8'h00;      memory[17651] <=  8'h00;      memory[17652] <=  8'h00;      memory[17653] <=  8'h00;      memory[17654] <=  8'h00;      memory[17655] <=  8'h00;      memory[17656] <=  8'h00;      memory[17657] <=  8'h00;      memory[17658] <=  8'h00;      memory[17659] <=  8'h00;      memory[17660] <=  8'h00;      memory[17661] <=  8'h00;      memory[17662] <=  8'h00;      memory[17663] <=  8'h00;      memory[17664] <=  8'h00;      memory[17665] <=  8'h00;      memory[17666] <=  8'h00;      memory[17667] <=  8'h00;      memory[17668] <=  8'h00;      memory[17669] <=  8'h00;      memory[17670] <=  8'h00;      memory[17671] <=  8'h00;      memory[17672] <=  8'h00;      memory[17673] <=  8'h00;      memory[17674] <=  8'h00;      memory[17675] <=  8'h00;      memory[17676] <=  8'h00;      memory[17677] <=  8'h00;      memory[17678] <=  8'h00;      memory[17679] <=  8'h00;      memory[17680] <=  8'h00;      memory[17681] <=  8'h00;      memory[17682] <=  8'h00;      memory[17683] <=  8'h00;      memory[17684] <=  8'h00;      memory[17685] <=  8'h00;      memory[17686] <=  8'h00;      memory[17687] <=  8'h00;      memory[17688] <=  8'h00;      memory[17689] <=  8'h00;      memory[17690] <=  8'h00;      memory[17691] <=  8'h00;      memory[17692] <=  8'h00;      memory[17693] <=  8'h00;      memory[17694] <=  8'h00;      memory[17695] <=  8'h00;      memory[17696] <=  8'h00;      memory[17697] <=  8'h00;      memory[17698] <=  8'h00;      memory[17699] <=  8'h00;      memory[17700] <=  8'h00;      memory[17701] <=  8'h00;      memory[17702] <=  8'h00;      memory[17703] <=  8'h00;      memory[17704] <=  8'h00;      memory[17705] <=  8'h00;      memory[17706] <=  8'h00;      memory[17707] <=  8'h00;      memory[17708] <=  8'h00;      memory[17709] <=  8'h00;      memory[17710] <=  8'h00;      memory[17711] <=  8'h00;      memory[17712] <=  8'h00;      memory[17713] <=  8'h00;      memory[17714] <=  8'h00;      memory[17715] <=  8'h00;      memory[17716] <=  8'h00;      memory[17717] <=  8'h00;      memory[17718] <=  8'h00;      memory[17719] <=  8'h00;      memory[17720] <=  8'h00;      memory[17721] <=  8'h00;      memory[17722] <=  8'h00;      memory[17723] <=  8'h00;      memory[17724] <=  8'h00;      memory[17725] <=  8'h00;      memory[17726] <=  8'h00;      memory[17727] <=  8'h00;      memory[17728] <=  8'h00;      memory[17729] <=  8'h00;      memory[17730] <=  8'h00;      memory[17731] <=  8'h00;      memory[17732] <=  8'h00;      memory[17733] <=  8'h00;      memory[17734] <=  8'h00;      memory[17735] <=  8'h00;      memory[17736] <=  8'h00;      memory[17737] <=  8'h00;      memory[17738] <=  8'h00;      memory[17739] <=  8'h00;      memory[17740] <=  8'h00;      memory[17741] <=  8'h00;      memory[17742] <=  8'h00;      memory[17743] <=  8'h00;      memory[17744] <=  8'h00;      memory[17745] <=  8'h00;      memory[17746] <=  8'h00;      memory[17747] <=  8'h00;      memory[17748] <=  8'h00;      memory[17749] <=  8'h00;      memory[17750] <=  8'h00;      memory[17751] <=  8'h00;      memory[17752] <=  8'h00;      memory[17753] <=  8'h00;      memory[17754] <=  8'h00;      memory[17755] <=  8'h00;      memory[17756] <=  8'h00;      memory[17757] <=  8'h00;      memory[17758] <=  8'h00;      memory[17759] <=  8'h00;      memory[17760] <=  8'h00;      memory[17761] <=  8'h00;      memory[17762] <=  8'h00;      memory[17763] <=  8'h00;      memory[17764] <=  8'h00;      memory[17765] <=  8'h00;      memory[17766] <=  8'h00;      memory[17767] <=  8'h00;      memory[17768] <=  8'h00;      memory[17769] <=  8'h00;      memory[17770] <=  8'h00;      memory[17771] <=  8'h00;      memory[17772] <=  8'h00;      memory[17773] <=  8'h00;      memory[17774] <=  8'h00;      memory[17775] <=  8'h00;      memory[17776] <=  8'h00;      memory[17777] <=  8'h00;      memory[17778] <=  8'h00;      memory[17779] <=  8'h00;      memory[17780] <=  8'h00;      memory[17781] <=  8'h00;      memory[17782] <=  8'h00;      memory[17783] <=  8'h00;      memory[17784] <=  8'h00;      memory[17785] <=  8'h00;      memory[17786] <=  8'h00;      memory[17787] <=  8'h00;      memory[17788] <=  8'h00;      memory[17789] <=  8'h00;      memory[17790] <=  8'h00;      memory[17791] <=  8'h00;      memory[17792] <=  8'h00;      memory[17793] <=  8'h00;      memory[17794] <=  8'h00;      memory[17795] <=  8'h00;      memory[17796] <=  8'h00;      memory[17797] <=  8'h00;      memory[17798] <=  8'h00;      memory[17799] <=  8'h00;      memory[17800] <=  8'h00;      memory[17801] <=  8'h00;      memory[17802] <=  8'h00;      memory[17803] <=  8'h00;      memory[17804] <=  8'h00;      memory[17805] <=  8'h00;      memory[17806] <=  8'h00;      memory[17807] <=  8'h00;      memory[17808] <=  8'h00;      memory[17809] <=  8'h00;      memory[17810] <=  8'h00;      memory[17811] <=  8'h00;      memory[17812] <=  8'h00;      memory[17813] <=  8'h00;      memory[17814] <=  8'h00;      memory[17815] <=  8'h00;      memory[17816] <=  8'h00;      memory[17817] <=  8'h00;      memory[17818] <=  8'h00;      memory[17819] <=  8'h00;      memory[17820] <=  8'h00;      memory[17821] <=  8'h00;      memory[17822] <=  8'h00;      memory[17823] <=  8'h00;      memory[17824] <=  8'h00;      memory[17825] <=  8'h00;      memory[17826] <=  8'h00;      memory[17827] <=  8'h00;      memory[17828] <=  8'h00;      memory[17829] <=  8'h00;      memory[17830] <=  8'h00;      memory[17831] <=  8'h00;      memory[17832] <=  8'h00;      memory[17833] <=  8'h00;      memory[17834] <=  8'h00;      memory[17835] <=  8'h00;      memory[17836] <=  8'h00;      memory[17837] <=  8'h00;      memory[17838] <=  8'h00;      memory[17839] <=  8'h00;      memory[17840] <=  8'h00;      memory[17841] <=  8'h00;      memory[17842] <=  8'h00;      memory[17843] <=  8'h00;      memory[17844] <=  8'h00;      memory[17845] <=  8'h00;      memory[17846] <=  8'h00;      memory[17847] <=  8'h00;      memory[17848] <=  8'h00;      memory[17849] <=  8'h00;      memory[17850] <=  8'h00;      memory[17851] <=  8'h00;      memory[17852] <=  8'h00;      memory[17853] <=  8'h00;      memory[17854] <=  8'h00;      memory[17855] <=  8'h00;      memory[17856] <=  8'h00;      memory[17857] <=  8'h00;      memory[17858] <=  8'h00;      memory[17859] <=  8'h00;      memory[17860] <=  8'h00;      memory[17861] <=  8'h00;      memory[17862] <=  8'h00;      memory[17863] <=  8'h00;      memory[17864] <=  8'h00;      memory[17865] <=  8'h00;      memory[17866] <=  8'h00;      memory[17867] <=  8'h00;      memory[17868] <=  8'h00;      memory[17869] <=  8'h00;      memory[17870] <=  8'h00;      memory[17871] <=  8'h00;      memory[17872] <=  8'h00;      memory[17873] <=  8'h00;      memory[17874] <=  8'h00;      memory[17875] <=  8'h00;      memory[17876] <=  8'h00;      memory[17877] <=  8'h00;      memory[17878] <=  8'h00;      memory[17879] <=  8'h00;      memory[17880] <=  8'h00;      memory[17881] <=  8'h00;      memory[17882] <=  8'h00;      memory[17883] <=  8'h00;      memory[17884] <=  8'h00;      memory[17885] <=  8'h00;      memory[17886] <=  8'h00;      memory[17887] <=  8'h00;      memory[17888] <=  8'h00;      memory[17889] <=  8'h00;      memory[17890] <=  8'h00;      memory[17891] <=  8'h00;      memory[17892] <=  8'h00;      memory[17893] <=  8'h00;      memory[17894] <=  8'h00;      memory[17895] <=  8'h00;      memory[17896] <=  8'h00;      memory[17897] <=  8'h00;      memory[17898] <=  8'h00;      memory[17899] <=  8'h00;      memory[17900] <=  8'h00;      memory[17901] <=  8'h00;      memory[17902] <=  8'h00;      memory[17903] <=  8'h00;      memory[17904] <=  8'h00;      memory[17905] <=  8'h00;      memory[17906] <=  8'h00;      memory[17907] <=  8'h00;      memory[17908] <=  8'h00;      memory[17909] <=  8'h00;      memory[17910] <=  8'h00;      memory[17911] <=  8'h00;      memory[17912] <=  8'h00;      memory[17913] <=  8'h00;      memory[17914] <=  8'h00;      memory[17915] <=  8'h00;      memory[17916] <=  8'h00;      memory[17917] <=  8'h00;      memory[17918] <=  8'h00;      memory[17919] <=  8'h00;      memory[17920] <=  8'h00;      memory[17921] <=  8'h00;      memory[17922] <=  8'h00;      memory[17923] <=  8'h00;      memory[17924] <=  8'h00;      memory[17925] <=  8'h00;      memory[17926] <=  8'h00;      memory[17927] <=  8'h00;      memory[17928] <=  8'h00;      memory[17929] <=  8'h00;      memory[17930] <=  8'h00;      memory[17931] <=  8'h00;      memory[17932] <=  8'h00;      memory[17933] <=  8'h00;      memory[17934] <=  8'h00;      memory[17935] <=  8'h00;      memory[17936] <=  8'h00;      memory[17937] <=  8'h00;      memory[17938] <=  8'h00;      memory[17939] <=  8'h00;      memory[17940] <=  8'h00;      memory[17941] <=  8'h00;      memory[17942] <=  8'h00;      memory[17943] <=  8'h00;      memory[17944] <=  8'h00;      memory[17945] <=  8'h00;      memory[17946] <=  8'h00;      memory[17947] <=  8'h00;      memory[17948] <=  8'h00;      memory[17949] <=  8'h00;      memory[17950] <=  8'h00;      memory[17951] <=  8'h00;      memory[17952] <=  8'h00;      memory[17953] <=  8'h00;      memory[17954] <=  8'h00;      memory[17955] <=  8'h00;      memory[17956] <=  8'h00;      memory[17957] <=  8'h00;      memory[17958] <=  8'h00;      memory[17959] <=  8'h00;      memory[17960] <=  8'h00;      memory[17961] <=  8'h00;      memory[17962] <=  8'h00;      memory[17963] <=  8'h00;      memory[17964] <=  8'h00;      memory[17965] <=  8'h00;      memory[17966] <=  8'h00;      memory[17967] <=  8'h00;      memory[17968] <=  8'h00;      memory[17969] <=  8'h00;      memory[17970] <=  8'h00;      memory[17971] <=  8'h00;      memory[17972] <=  8'h00;      memory[17973] <=  8'h00;      memory[17974] <=  8'h00;      memory[17975] <=  8'h00;      memory[17976] <=  8'h00;      memory[17977] <=  8'h00;      memory[17978] <=  8'h00;      memory[17979] <=  8'h00;      memory[17980] <=  8'h00;      memory[17981] <=  8'h00;      memory[17982] <=  8'h00;      memory[17983] <=  8'h00;      memory[17984] <=  8'h00;      memory[17985] <=  8'h00;      memory[17986] <=  8'h00;      memory[17987] <=  8'h00;      memory[17988] <=  8'h00;      memory[17989] <=  8'h00;      memory[17990] <=  8'h00;      memory[17991] <=  8'h00;      memory[17992] <=  8'h00;      memory[17993] <=  8'h00;      memory[17994] <=  8'h00;      memory[17995] <=  8'h00;      memory[17996] <=  8'h00;      memory[17997] <=  8'h00;      memory[17998] <=  8'h00;      memory[17999] <=  8'h00;      memory[18000] <=  8'h00;      memory[18001] <=  8'h00;      memory[18002] <=  8'h00;      memory[18003] <=  8'h00;      memory[18004] <=  8'h00;      memory[18005] <=  8'h00;      memory[18006] <=  8'h00;      memory[18007] <=  8'h00;      memory[18008] <=  8'h00;      memory[18009] <=  8'h00;      memory[18010] <=  8'h00;      memory[18011] <=  8'h00;      memory[18012] <=  8'h00;      memory[18013] <=  8'h00;      memory[18014] <=  8'h00;      memory[18015] <=  8'h00;      memory[18016] <=  8'h00;      memory[18017] <=  8'h00;      memory[18018] <=  8'h00;      memory[18019] <=  8'h00;      memory[18020] <=  8'h00;      memory[18021] <=  8'h00;      memory[18022] <=  8'h00;      memory[18023] <=  8'h00;      memory[18024] <=  8'h00;      memory[18025] <=  8'h00;      memory[18026] <=  8'h00;      memory[18027] <=  8'h00;      memory[18028] <=  8'h00;      memory[18029] <=  8'h00;      memory[18030] <=  8'h00;      memory[18031] <=  8'h00;      memory[18032] <=  8'h00;      memory[18033] <=  8'h00;      memory[18034] <=  8'h00;      memory[18035] <=  8'h00;      memory[18036] <=  8'h00;      memory[18037] <=  8'h00;      memory[18038] <=  8'h00;      memory[18039] <=  8'h00;      memory[18040] <=  8'h00;      memory[18041] <=  8'h00;      memory[18042] <=  8'h00;      memory[18043] <=  8'h00;      memory[18044] <=  8'h00;      memory[18045] <=  8'h00;      memory[18046] <=  8'h00;      memory[18047] <=  8'h00;      memory[18048] <=  8'h00;      memory[18049] <=  8'h00;      memory[18050] <=  8'h00;      memory[18051] <=  8'h00;      memory[18052] <=  8'h00;      memory[18053] <=  8'h00;      memory[18054] <=  8'h00;      memory[18055] <=  8'h00;      memory[18056] <=  8'h00;      memory[18057] <=  8'h00;      memory[18058] <=  8'h00;      memory[18059] <=  8'h00;      memory[18060] <=  8'h00;      memory[18061] <=  8'h00;      memory[18062] <=  8'h00;      memory[18063] <=  8'h00;      memory[18064] <=  8'h00;      memory[18065] <=  8'h00;      memory[18066] <=  8'h00;      memory[18067] <=  8'h00;      memory[18068] <=  8'h00;      memory[18069] <=  8'h00;      memory[18070] <=  8'h00;      memory[18071] <=  8'h00;      memory[18072] <=  8'h00;      memory[18073] <=  8'h00;      memory[18074] <=  8'h00;      memory[18075] <=  8'h00;      memory[18076] <=  8'h00;      memory[18077] <=  8'h00;      memory[18078] <=  8'h00;      memory[18079] <=  8'h00;      memory[18080] <=  8'h00;      memory[18081] <=  8'h00;      memory[18082] <=  8'h00;      memory[18083] <=  8'h00;      memory[18084] <=  8'h00;      memory[18085] <=  8'h00;      memory[18086] <=  8'h00;      memory[18087] <=  8'h00;      memory[18088] <=  8'h00;      memory[18089] <=  8'h00;      memory[18090] <=  8'h00;      memory[18091] <=  8'h00;      memory[18092] <=  8'h00;      memory[18093] <=  8'h00;      memory[18094] <=  8'h00;      memory[18095] <=  8'h00;      memory[18096] <=  8'h00;      memory[18097] <=  8'h00;      memory[18098] <=  8'h00;      memory[18099] <=  8'h00;      memory[18100] <=  8'h00;      memory[18101] <=  8'h00;      memory[18102] <=  8'h00;      memory[18103] <=  8'h00;      memory[18104] <=  8'h00;      memory[18105] <=  8'h00;      memory[18106] <=  8'h00;      memory[18107] <=  8'h00;      memory[18108] <=  8'h00;      memory[18109] <=  8'h00;      memory[18110] <=  8'h00;      memory[18111] <=  8'h00;      memory[18112] <=  8'h00;      memory[18113] <=  8'h00;      memory[18114] <=  8'h00;      memory[18115] <=  8'h00;      memory[18116] <=  8'h00;      memory[18117] <=  8'h00;      memory[18118] <=  8'h00;      memory[18119] <=  8'h00;      memory[18120] <=  8'h00;      memory[18121] <=  8'h00;      memory[18122] <=  8'h00;      memory[18123] <=  8'h00;      memory[18124] <=  8'h00;      memory[18125] <=  8'h00;      memory[18126] <=  8'h00;      memory[18127] <=  8'h00;      memory[18128] <=  8'h00;      memory[18129] <=  8'h00;      memory[18130] <=  8'h00;      memory[18131] <=  8'h00;      memory[18132] <=  8'h00;      memory[18133] <=  8'h00;      memory[18134] <=  8'h00;      memory[18135] <=  8'h00;      memory[18136] <=  8'h00;      memory[18137] <=  8'h00;      memory[18138] <=  8'h00;      memory[18139] <=  8'h00;      memory[18140] <=  8'h00;      memory[18141] <=  8'h00;      memory[18142] <=  8'h00;      memory[18143] <=  8'h00;      memory[18144] <=  8'h00;      memory[18145] <=  8'h00;      memory[18146] <=  8'h00;      memory[18147] <=  8'h00;      memory[18148] <=  8'h00;      memory[18149] <=  8'h00;      memory[18150] <=  8'h00;      memory[18151] <=  8'h00;      memory[18152] <=  8'h00;      memory[18153] <=  8'h00;      memory[18154] <=  8'h00;      memory[18155] <=  8'h00;      memory[18156] <=  8'h00;      memory[18157] <=  8'h00;      memory[18158] <=  8'h00;      memory[18159] <=  8'h00;      memory[18160] <=  8'h00;      memory[18161] <=  8'h00;      memory[18162] <=  8'h00;      memory[18163] <=  8'h00;      memory[18164] <=  8'h00;      memory[18165] <=  8'h00;      memory[18166] <=  8'h00;      memory[18167] <=  8'h00;      memory[18168] <=  8'h00;      memory[18169] <=  8'h00;      memory[18170] <=  8'h00;      memory[18171] <=  8'h00;      memory[18172] <=  8'h00;      memory[18173] <=  8'h00;      memory[18174] <=  8'h00;      memory[18175] <=  8'h00;      memory[18176] <=  8'h00;      memory[18177] <=  8'h00;      memory[18178] <=  8'h00;      memory[18179] <=  8'h00;      memory[18180] <=  8'h00;      memory[18181] <=  8'h00;      memory[18182] <=  8'h00;      memory[18183] <=  8'h00;      memory[18184] <=  8'h00;      memory[18185] <=  8'h00;      memory[18186] <=  8'h00;      memory[18187] <=  8'h00;      memory[18188] <=  8'h00;      memory[18189] <=  8'h00;      memory[18190] <=  8'h00;      memory[18191] <=  8'h00;      memory[18192] <=  8'h00;      memory[18193] <=  8'h00;      memory[18194] <=  8'h00;      memory[18195] <=  8'h00;      memory[18196] <=  8'h00;      memory[18197] <=  8'h00;      memory[18198] <=  8'h00;      memory[18199] <=  8'h00;      memory[18200] <=  8'h00;      memory[18201] <=  8'h00;      memory[18202] <=  8'h00;      memory[18203] <=  8'h00;      memory[18204] <=  8'h00;      memory[18205] <=  8'h00;      memory[18206] <=  8'h00;      memory[18207] <=  8'h00;      memory[18208] <=  8'h00;      memory[18209] <=  8'h00;      memory[18210] <=  8'h00;      memory[18211] <=  8'h00;      memory[18212] <=  8'h00;      memory[18213] <=  8'h00;      memory[18214] <=  8'h00;      memory[18215] <=  8'h00;      memory[18216] <=  8'h00;      memory[18217] <=  8'h00;      memory[18218] <=  8'h00;      memory[18219] <=  8'h00;      memory[18220] <=  8'h00;      memory[18221] <=  8'h00;      memory[18222] <=  8'h00;      memory[18223] <=  8'h00;      memory[18224] <=  8'h00;      memory[18225] <=  8'h00;      memory[18226] <=  8'h00;      memory[18227] <=  8'h00;      memory[18228] <=  8'h00;      memory[18229] <=  8'h00;      memory[18230] <=  8'h00;      memory[18231] <=  8'h00;      memory[18232] <=  8'h00;      memory[18233] <=  8'h00;      memory[18234] <=  8'h00;      memory[18235] <=  8'h00;      memory[18236] <=  8'h00;      memory[18237] <=  8'h00;      memory[18238] <=  8'h00;      memory[18239] <=  8'h00;      memory[18240] <=  8'h00;      memory[18241] <=  8'h00;      memory[18242] <=  8'h00;      memory[18243] <=  8'h00;      memory[18244] <=  8'h00;      memory[18245] <=  8'h00;      memory[18246] <=  8'h00;      memory[18247] <=  8'h00;      memory[18248] <=  8'h00;      memory[18249] <=  8'h00;      memory[18250] <=  8'h00;      memory[18251] <=  8'h00;      memory[18252] <=  8'h00;      memory[18253] <=  8'h00;      memory[18254] <=  8'h00;      memory[18255] <=  8'h00;      memory[18256] <=  8'h00;      memory[18257] <=  8'h00;      memory[18258] <=  8'h00;      memory[18259] <=  8'h00;      memory[18260] <=  8'h00;      memory[18261] <=  8'h00;      memory[18262] <=  8'h00;      memory[18263] <=  8'h00;      memory[18264] <=  8'h00;      memory[18265] <=  8'h00;      memory[18266] <=  8'h00;      memory[18267] <=  8'h00;      memory[18268] <=  8'h00;      memory[18269] <=  8'h00;      memory[18270] <=  8'h00;      memory[18271] <=  8'h00;      memory[18272] <=  8'h00;      memory[18273] <=  8'h00;      memory[18274] <=  8'h00;      memory[18275] <=  8'h00;      memory[18276] <=  8'h00;      memory[18277] <=  8'h00;      memory[18278] <=  8'h00;      memory[18279] <=  8'h00;      memory[18280] <=  8'h00;      memory[18281] <=  8'h00;      memory[18282] <=  8'h00;      memory[18283] <=  8'h00;      memory[18284] <=  8'h00;      memory[18285] <=  8'h00;      memory[18286] <=  8'h00;      memory[18287] <=  8'h00;      memory[18288] <=  8'h00;      memory[18289] <=  8'h00;      memory[18290] <=  8'h00;      memory[18291] <=  8'h00;      memory[18292] <=  8'h00;      memory[18293] <=  8'h00;      memory[18294] <=  8'h00;      memory[18295] <=  8'h00;      memory[18296] <=  8'h00;      memory[18297] <=  8'h00;      memory[18298] <=  8'h00;      memory[18299] <=  8'h00;      memory[18300] <=  8'h00;      memory[18301] <=  8'h00;      memory[18302] <=  8'h00;      memory[18303] <=  8'h00;      memory[18304] <=  8'h00;      memory[18305] <=  8'h00;      memory[18306] <=  8'h00;      memory[18307] <=  8'h00;      memory[18308] <=  8'h00;      memory[18309] <=  8'h00;      memory[18310] <=  8'h00;      memory[18311] <=  8'h00;      memory[18312] <=  8'h00;      memory[18313] <=  8'h00;      memory[18314] <=  8'h00;      memory[18315] <=  8'h00;      memory[18316] <=  8'h00;      memory[18317] <=  8'h00;      memory[18318] <=  8'h00;      memory[18319] <=  8'h00;      memory[18320] <=  8'h00;      memory[18321] <=  8'h00;      memory[18322] <=  8'h00;      memory[18323] <=  8'h00;      memory[18324] <=  8'h00;      memory[18325] <=  8'h00;      memory[18326] <=  8'h00;      memory[18327] <=  8'h00;      memory[18328] <=  8'h00;      memory[18329] <=  8'h00;      memory[18330] <=  8'h00;      memory[18331] <=  8'h00;      memory[18332] <=  8'h00;      memory[18333] <=  8'h00;      memory[18334] <=  8'h00;      memory[18335] <=  8'h00;      memory[18336] <=  8'h00;      memory[18337] <=  8'h00;      memory[18338] <=  8'h00;      memory[18339] <=  8'h00;      memory[18340] <=  8'h00;      memory[18341] <=  8'h00;      memory[18342] <=  8'h00;      memory[18343] <=  8'h00;      memory[18344] <=  8'h00;      memory[18345] <=  8'h00;      memory[18346] <=  8'h00;      memory[18347] <=  8'h00;      memory[18348] <=  8'h00;      memory[18349] <=  8'h00;      memory[18350] <=  8'h00;      memory[18351] <=  8'h00;      memory[18352] <=  8'h00;      memory[18353] <=  8'h00;      memory[18354] <=  8'h00;      memory[18355] <=  8'h00;      memory[18356] <=  8'h00;      memory[18357] <=  8'h00;      memory[18358] <=  8'h00;      memory[18359] <=  8'h00;      memory[18360] <=  8'h00;      memory[18361] <=  8'h00;      memory[18362] <=  8'h00;      memory[18363] <=  8'h00;      memory[18364] <=  8'h00;      memory[18365] <=  8'h00;      memory[18366] <=  8'h00;      memory[18367] <=  8'h00;      memory[18368] <=  8'h00;      memory[18369] <=  8'h00;      memory[18370] <=  8'h00;      memory[18371] <=  8'h00;      memory[18372] <=  8'h00;      memory[18373] <=  8'h00;      memory[18374] <=  8'h00;      memory[18375] <=  8'h00;      memory[18376] <=  8'h00;      memory[18377] <=  8'h00;      memory[18378] <=  8'h00;      memory[18379] <=  8'h00;      memory[18380] <=  8'h00;      memory[18381] <=  8'h00;      memory[18382] <=  8'h00;      memory[18383] <=  8'h00;      memory[18384] <=  8'h00;      memory[18385] <=  8'h00;      memory[18386] <=  8'h00;      memory[18387] <=  8'h00;      memory[18388] <=  8'h00;      memory[18389] <=  8'h00;      memory[18390] <=  8'h00;      memory[18391] <=  8'h00;      memory[18392] <=  8'h00;      memory[18393] <=  8'h00;      memory[18394] <=  8'h00;      memory[18395] <=  8'h00;      memory[18396] <=  8'h00;      memory[18397] <=  8'h00;      memory[18398] <=  8'h00;      memory[18399] <=  8'h00;      memory[18400] <=  8'h00;      memory[18401] <=  8'h00;      memory[18402] <=  8'h00;      memory[18403] <=  8'h00;      memory[18404] <=  8'h00;      memory[18405] <=  8'h00;      memory[18406] <=  8'h00;      memory[18407] <=  8'h00;      memory[18408] <=  8'h00;      memory[18409] <=  8'h00;      memory[18410] <=  8'h00;      memory[18411] <=  8'h00;      memory[18412] <=  8'h00;      memory[18413] <=  8'h00;      memory[18414] <=  8'h00;      memory[18415] <=  8'h00;      memory[18416] <=  8'h00;      memory[18417] <=  8'h00;      memory[18418] <=  8'h00;      memory[18419] <=  8'h00;      memory[18420] <=  8'h00;      memory[18421] <=  8'h00;      memory[18422] <=  8'h00;      memory[18423] <=  8'h00;      memory[18424] <=  8'h00;      memory[18425] <=  8'h00;      memory[18426] <=  8'h00;      memory[18427] <=  8'h00;      memory[18428] <=  8'h00;      memory[18429] <=  8'h00;      memory[18430] <=  8'h00;      memory[18431] <=  8'h00;      memory[18432] <=  8'h00;      memory[18433] <=  8'h00;      memory[18434] <=  8'h00;      memory[18435] <=  8'h00;      memory[18436] <=  8'h00;      memory[18437] <=  8'h00;      memory[18438] <=  8'h00;      memory[18439] <=  8'h00;      memory[18440] <=  8'h00;      memory[18441] <=  8'h00;      memory[18442] <=  8'h00;      memory[18443] <=  8'h00;      memory[18444] <=  8'h00;      memory[18445] <=  8'h00;      memory[18446] <=  8'h00;      memory[18447] <=  8'h00;      memory[18448] <=  8'h00;      memory[18449] <=  8'h00;      memory[18450] <=  8'h00;      memory[18451] <=  8'h00;      memory[18452] <=  8'h00;      memory[18453] <=  8'h00;      memory[18454] <=  8'h00;      memory[18455] <=  8'h00;      memory[18456] <=  8'h00;      memory[18457] <=  8'h00;      memory[18458] <=  8'h00;      memory[18459] <=  8'h00;      memory[18460] <=  8'h00;      memory[18461] <=  8'h00;      memory[18462] <=  8'h00;      memory[18463] <=  8'h00;      memory[18464] <=  8'h00;      memory[18465] <=  8'h00;      memory[18466] <=  8'h00;      memory[18467] <=  8'h00;      memory[18468] <=  8'h00;      memory[18469] <=  8'h00;      memory[18470] <=  8'h00;      memory[18471] <=  8'h00;      memory[18472] <=  8'h00;      memory[18473] <=  8'h00;      memory[18474] <=  8'h00;      memory[18475] <=  8'h00;      memory[18476] <=  8'h00;      memory[18477] <=  8'h00;      memory[18478] <=  8'h00;      memory[18479] <=  8'h00;      memory[18480] <=  8'h00;      memory[18481] <=  8'h00;      memory[18482] <=  8'h00;      memory[18483] <=  8'h00;      memory[18484] <=  8'h00;      memory[18485] <=  8'h00;      memory[18486] <=  8'h00;      memory[18487] <=  8'h00;      memory[18488] <=  8'h00;      memory[18489] <=  8'h00;      memory[18490] <=  8'h00;      memory[18491] <=  8'h00;      memory[18492] <=  8'h00;      memory[18493] <=  8'h00;      memory[18494] <=  8'h00;      memory[18495] <=  8'h00;      memory[18496] <=  8'h00;      memory[18497] <=  8'h00;      memory[18498] <=  8'h00;      memory[18499] <=  8'h00;      memory[18500] <=  8'h00;      memory[18501] <=  8'h00;      memory[18502] <=  8'h00;      memory[18503] <=  8'h00;      memory[18504] <=  8'h00;      memory[18505] <=  8'h00;      memory[18506] <=  8'h00;      memory[18507] <=  8'h00;      memory[18508] <=  8'h00;      memory[18509] <=  8'h00;      memory[18510] <=  8'h00;      memory[18511] <=  8'h00;      memory[18512] <=  8'h00;      memory[18513] <=  8'h00;      memory[18514] <=  8'h00;      memory[18515] <=  8'h00;      memory[18516] <=  8'h00;      memory[18517] <=  8'h00;      memory[18518] <=  8'h00;      memory[18519] <=  8'h00;      memory[18520] <=  8'h00;      memory[18521] <=  8'h00;      memory[18522] <=  8'h00;      memory[18523] <=  8'h00;      memory[18524] <=  8'h00;      memory[18525] <=  8'h00;      memory[18526] <=  8'h00;      memory[18527] <=  8'h00;      memory[18528] <=  8'h00;      memory[18529] <=  8'h00;      memory[18530] <=  8'h00;      memory[18531] <=  8'h00;      memory[18532] <=  8'h00;      memory[18533] <=  8'h00;      memory[18534] <=  8'h00;      memory[18535] <=  8'h00;      memory[18536] <=  8'h00;      memory[18537] <=  8'h00;      memory[18538] <=  8'h00;      memory[18539] <=  8'h00;      memory[18540] <=  8'h00;      memory[18541] <=  8'h00;      memory[18542] <=  8'h00;      memory[18543] <=  8'h00;      memory[18544] <=  8'h00;      memory[18545] <=  8'h00;      memory[18546] <=  8'h00;      memory[18547] <=  8'h00;      memory[18548] <=  8'h00;      memory[18549] <=  8'h00;      memory[18550] <=  8'h00;      memory[18551] <=  8'h00;      memory[18552] <=  8'h00;      memory[18553] <=  8'h00;      memory[18554] <=  8'h00;      memory[18555] <=  8'h00;      memory[18556] <=  8'h00;      memory[18557] <=  8'h00;      memory[18558] <=  8'h00;      memory[18559] <=  8'h00;      memory[18560] <=  8'h00;      memory[18561] <=  8'h00;      memory[18562] <=  8'h00;      memory[18563] <=  8'h00;      memory[18564] <=  8'h00;      memory[18565] <=  8'h00;      memory[18566] <=  8'h00;      memory[18567] <=  8'h00;      memory[18568] <=  8'h00;      memory[18569] <=  8'h00;      memory[18570] <=  8'h00;      memory[18571] <=  8'h00;      memory[18572] <=  8'h00;      memory[18573] <=  8'h00;      memory[18574] <=  8'h00;      memory[18575] <=  8'h00;      memory[18576] <=  8'h00;      memory[18577] <=  8'h00;      memory[18578] <=  8'h00;      memory[18579] <=  8'h00;      memory[18580] <=  8'h00;      memory[18581] <=  8'h00;      memory[18582] <=  8'h00;      memory[18583] <=  8'h00;      memory[18584] <=  8'h00;      memory[18585] <=  8'h00;      memory[18586] <=  8'h00;      memory[18587] <=  8'h00;      memory[18588] <=  8'h00;      memory[18589] <=  8'h00;      memory[18590] <=  8'h00;      memory[18591] <=  8'h00;      memory[18592] <=  8'h00;      memory[18593] <=  8'h00;      memory[18594] <=  8'h00;      memory[18595] <=  8'h00;      memory[18596] <=  8'h00;      memory[18597] <=  8'h00;      memory[18598] <=  8'h00;      memory[18599] <=  8'h00;      memory[18600] <=  8'h00;      memory[18601] <=  8'h00;      memory[18602] <=  8'h00;      memory[18603] <=  8'h00;      memory[18604] <=  8'h00;      memory[18605] <=  8'h00;      memory[18606] <=  8'h00;      memory[18607] <=  8'h00;      memory[18608] <=  8'h00;      memory[18609] <=  8'h00;      memory[18610] <=  8'h00;      memory[18611] <=  8'h00;      memory[18612] <=  8'h00;      memory[18613] <=  8'h00;      memory[18614] <=  8'h00;      memory[18615] <=  8'h00;      memory[18616] <=  8'h00;      memory[18617] <=  8'h00;      memory[18618] <=  8'h00;      memory[18619] <=  8'h00;      memory[18620] <=  8'h00;      memory[18621] <=  8'h00;      memory[18622] <=  8'h00;      memory[18623] <=  8'h00;      memory[18624] <=  8'h00;      memory[18625] <=  8'h00;      memory[18626] <=  8'h00;      memory[18627] <=  8'h00;      memory[18628] <=  8'h00;      memory[18629] <=  8'h00;      memory[18630] <=  8'h00;      memory[18631] <=  8'h00;      memory[18632] <=  8'h00;      memory[18633] <=  8'h00;      memory[18634] <=  8'h00;      memory[18635] <=  8'h00;      memory[18636] <=  8'h00;      memory[18637] <=  8'h00;      memory[18638] <=  8'h00;      memory[18639] <=  8'h00;      memory[18640] <=  8'h00;      memory[18641] <=  8'h00;      memory[18642] <=  8'h00;      memory[18643] <=  8'h00;      memory[18644] <=  8'h00;      memory[18645] <=  8'h00;      memory[18646] <=  8'h00;      memory[18647] <=  8'h00;      memory[18648] <=  8'h00;      memory[18649] <=  8'h00;      memory[18650] <=  8'h00;      memory[18651] <=  8'h00;      memory[18652] <=  8'h00;      memory[18653] <=  8'h00;      memory[18654] <=  8'h00;      memory[18655] <=  8'h00;      memory[18656] <=  8'h00;      memory[18657] <=  8'h00;      memory[18658] <=  8'h00;      memory[18659] <=  8'h00;      memory[18660] <=  8'h00;      memory[18661] <=  8'h00;      memory[18662] <=  8'h00;      memory[18663] <=  8'h00;      memory[18664] <=  8'h00;      memory[18665] <=  8'h00;      memory[18666] <=  8'h00;      memory[18667] <=  8'h00;      memory[18668] <=  8'h00;      memory[18669] <=  8'h00;      memory[18670] <=  8'h00;      memory[18671] <=  8'h00;      memory[18672] <=  8'h00;      memory[18673] <=  8'h00;      memory[18674] <=  8'h00;      memory[18675] <=  8'h00;      memory[18676] <=  8'h00;      memory[18677] <=  8'h00;      memory[18678] <=  8'h00;      memory[18679] <=  8'h00;      memory[18680] <=  8'h00;      memory[18681] <=  8'h00;      memory[18682] <=  8'h00;      memory[18683] <=  8'h00;      memory[18684] <=  8'h00;      memory[18685] <=  8'h00;      memory[18686] <=  8'h00;      memory[18687] <=  8'h00;      memory[18688] <=  8'h00;      memory[18689] <=  8'h00;      memory[18690] <=  8'h00;      memory[18691] <=  8'h00;      memory[18692] <=  8'h00;      memory[18693] <=  8'h00;      memory[18694] <=  8'h00;      memory[18695] <=  8'h00;      memory[18696] <=  8'h00;      memory[18697] <=  8'h00;      memory[18698] <=  8'h00;      memory[18699] <=  8'h00;      memory[18700] <=  8'h00;      memory[18701] <=  8'h00;      memory[18702] <=  8'h00;      memory[18703] <=  8'h00;      memory[18704] <=  8'h00;      memory[18705] <=  8'h00;      memory[18706] <=  8'h00;      memory[18707] <=  8'h00;      memory[18708] <=  8'h00;      memory[18709] <=  8'h00;      memory[18710] <=  8'h00;      memory[18711] <=  8'h00;      memory[18712] <=  8'h00;      memory[18713] <=  8'h00;      memory[18714] <=  8'h00;      memory[18715] <=  8'h00;      memory[18716] <=  8'h00;      memory[18717] <=  8'h00;      memory[18718] <=  8'h00;      memory[18719] <=  8'h00;      memory[18720] <=  8'h00;      memory[18721] <=  8'h00;      memory[18722] <=  8'h00;      memory[18723] <=  8'h00;      memory[18724] <=  8'h00;      memory[18725] <=  8'h00;      memory[18726] <=  8'h00;      memory[18727] <=  8'h00;      memory[18728] <=  8'h00;      memory[18729] <=  8'h00;      memory[18730] <=  8'h00;      memory[18731] <=  8'h00;      memory[18732] <=  8'h00;      memory[18733] <=  8'h00;      memory[18734] <=  8'h00;      memory[18735] <=  8'h00;      memory[18736] <=  8'h00;      memory[18737] <=  8'h00;      memory[18738] <=  8'h00;      memory[18739] <=  8'h00;      memory[18740] <=  8'h00;      memory[18741] <=  8'h00;      memory[18742] <=  8'h00;      memory[18743] <=  8'h00;      memory[18744] <=  8'h00;      memory[18745] <=  8'h00;      memory[18746] <=  8'h00;      memory[18747] <=  8'h00;      memory[18748] <=  8'h00;      memory[18749] <=  8'h00;      memory[18750] <=  8'h00;      memory[18751] <=  8'h00;      memory[18752] <=  8'h00;      memory[18753] <=  8'h00;      memory[18754] <=  8'h00;      memory[18755] <=  8'h00;      memory[18756] <=  8'h00;      memory[18757] <=  8'h00;      memory[18758] <=  8'h00;      memory[18759] <=  8'h00;      memory[18760] <=  8'h00;      memory[18761] <=  8'h00;      memory[18762] <=  8'h00;      memory[18763] <=  8'h00;      memory[18764] <=  8'h00;      memory[18765] <=  8'h00;      memory[18766] <=  8'h00;      memory[18767] <=  8'h00;      memory[18768] <=  8'h00;      memory[18769] <=  8'h00;      memory[18770] <=  8'h00;      memory[18771] <=  8'h00;      memory[18772] <=  8'h00;      memory[18773] <=  8'h00;      memory[18774] <=  8'h00;      memory[18775] <=  8'h00;      memory[18776] <=  8'h00;      memory[18777] <=  8'h00;      memory[18778] <=  8'h00;      memory[18779] <=  8'h00;      memory[18780] <=  8'h00;      memory[18781] <=  8'h00;      memory[18782] <=  8'h00;      memory[18783] <=  8'h00;      memory[18784] <=  8'h00;      memory[18785] <=  8'h00;      memory[18786] <=  8'h00;      memory[18787] <=  8'h00;      memory[18788] <=  8'h00;      memory[18789] <=  8'h00;      memory[18790] <=  8'h00;      memory[18791] <=  8'h00;      memory[18792] <=  8'h00;      memory[18793] <=  8'h00;      memory[18794] <=  8'h00;      memory[18795] <=  8'h00;      memory[18796] <=  8'h00;      memory[18797] <=  8'h00;      memory[18798] <=  8'h00;      memory[18799] <=  8'h00;      memory[18800] <=  8'h00;      memory[18801] <=  8'h00;      memory[18802] <=  8'h00;      memory[18803] <=  8'h00;      memory[18804] <=  8'h00;      memory[18805] <=  8'h00;      memory[18806] <=  8'h00;      memory[18807] <=  8'h00;      memory[18808] <=  8'h00;      memory[18809] <=  8'h00;      memory[18810] <=  8'h00;      memory[18811] <=  8'h00;      memory[18812] <=  8'h00;      memory[18813] <=  8'h00;      memory[18814] <=  8'h00;      memory[18815] <=  8'h00;      memory[18816] <=  8'h00;      memory[18817] <=  8'h00;      memory[18818] <=  8'h00;      memory[18819] <=  8'h00;      memory[18820] <=  8'h00;      memory[18821] <=  8'h00;      memory[18822] <=  8'h00;      memory[18823] <=  8'h00;      memory[18824] <=  8'h00;      memory[18825] <=  8'h00;      memory[18826] <=  8'h00;      memory[18827] <=  8'h00;      memory[18828] <=  8'h00;      memory[18829] <=  8'h00;      memory[18830] <=  8'h00;      memory[18831] <=  8'h00;      memory[18832] <=  8'h00;      memory[18833] <=  8'h00;      memory[18834] <=  8'h00;      memory[18835] <=  8'h00;      memory[18836] <=  8'h00;      memory[18837] <=  8'h00;      memory[18838] <=  8'h00;      memory[18839] <=  8'h00;      memory[18840] <=  8'h00;      memory[18841] <=  8'h00;      memory[18842] <=  8'h00;      memory[18843] <=  8'h00;      memory[18844] <=  8'h00;      memory[18845] <=  8'h00;      memory[18846] <=  8'h00;      memory[18847] <=  8'h00;      memory[18848] <=  8'h00;      memory[18849] <=  8'h00;      memory[18850] <=  8'h00;      memory[18851] <=  8'h00;      memory[18852] <=  8'h00;      memory[18853] <=  8'h00;      memory[18854] <=  8'h00;      memory[18855] <=  8'h00;      memory[18856] <=  8'h00;      memory[18857] <=  8'h00;      memory[18858] <=  8'h00;      memory[18859] <=  8'h00;      memory[18860] <=  8'h00;      memory[18861] <=  8'h00;      memory[18862] <=  8'h00;      memory[18863] <=  8'h00;      memory[18864] <=  8'h00;      memory[18865] <=  8'h00;      memory[18866] <=  8'h00;      memory[18867] <=  8'h00;      memory[18868] <=  8'h00;      memory[18869] <=  8'h00;      memory[18870] <=  8'h00;      memory[18871] <=  8'h00;      memory[18872] <=  8'h00;      memory[18873] <=  8'h00;      memory[18874] <=  8'h00;      memory[18875] <=  8'h00;      memory[18876] <=  8'h00;      memory[18877] <=  8'h00;      memory[18878] <=  8'h00;      memory[18879] <=  8'h00;      memory[18880] <=  8'h00;      memory[18881] <=  8'h00;      memory[18882] <=  8'h00;      memory[18883] <=  8'h00;      memory[18884] <=  8'h00;      memory[18885] <=  8'h00;      memory[18886] <=  8'h00;      memory[18887] <=  8'h00;      memory[18888] <=  8'h00;      memory[18889] <=  8'h00;      memory[18890] <=  8'h00;      memory[18891] <=  8'h00;      memory[18892] <=  8'h00;      memory[18893] <=  8'h00;      memory[18894] <=  8'h00;      memory[18895] <=  8'h00;      memory[18896] <=  8'h00;      memory[18897] <=  8'h00;      memory[18898] <=  8'h00;      memory[18899] <=  8'h00;      memory[18900] <=  8'h00;      memory[18901] <=  8'h00;      memory[18902] <=  8'h00;      memory[18903] <=  8'h00;      memory[18904] <=  8'h00;      memory[18905] <=  8'h00;      memory[18906] <=  8'h00;      memory[18907] <=  8'h00;      memory[18908] <=  8'h00;      memory[18909] <=  8'h00;      memory[18910] <=  8'h00;      memory[18911] <=  8'h00;      memory[18912] <=  8'h00;      memory[18913] <=  8'h00;      memory[18914] <=  8'h00;      memory[18915] <=  8'h00;      memory[18916] <=  8'h00;      memory[18917] <=  8'h00;      memory[18918] <=  8'h00;      memory[18919] <=  8'h00;      memory[18920] <=  8'h00;      memory[18921] <=  8'h00;      memory[18922] <=  8'h00;      memory[18923] <=  8'h00;      memory[18924] <=  8'h00;      memory[18925] <=  8'h00;      memory[18926] <=  8'h00;      memory[18927] <=  8'h00;      memory[18928] <=  8'h00;      memory[18929] <=  8'h00;      memory[18930] <=  8'h00;      memory[18931] <=  8'h00;      memory[18932] <=  8'h00;      memory[18933] <=  8'h00;      memory[18934] <=  8'h00;      memory[18935] <=  8'h00;      memory[18936] <=  8'h00;      memory[18937] <=  8'h00;      memory[18938] <=  8'h00;      memory[18939] <=  8'h00;      memory[18940] <=  8'h00;      memory[18941] <=  8'h00;      memory[18942] <=  8'h00;      memory[18943] <=  8'h00;      memory[18944] <=  8'h00;      memory[18945] <=  8'h00;      memory[18946] <=  8'h00;      memory[18947] <=  8'h00;      memory[18948] <=  8'h00;      memory[18949] <=  8'h00;      memory[18950] <=  8'h00;      memory[18951] <=  8'h00;      memory[18952] <=  8'h00;      memory[18953] <=  8'h00;      memory[18954] <=  8'h00;      memory[18955] <=  8'h00;      memory[18956] <=  8'h00;      memory[18957] <=  8'h00;      memory[18958] <=  8'h00;      memory[18959] <=  8'h00;      memory[18960] <=  8'h00;      memory[18961] <=  8'h00;      memory[18962] <=  8'h00;      memory[18963] <=  8'h00;      memory[18964] <=  8'h00;      memory[18965] <=  8'h00;      memory[18966] <=  8'h00;      memory[18967] <=  8'h00;      memory[18968] <=  8'h00;      memory[18969] <=  8'h00;      memory[18970] <=  8'h00;      memory[18971] <=  8'h00;      memory[18972] <=  8'h00;      memory[18973] <=  8'h00;      memory[18974] <=  8'h00;      memory[18975] <=  8'h00;      memory[18976] <=  8'h00;      memory[18977] <=  8'h00;      memory[18978] <=  8'h00;      memory[18979] <=  8'h00;      memory[18980] <=  8'h00;      memory[18981] <=  8'h00;      memory[18982] <=  8'h00;      memory[18983] <=  8'h00;      memory[18984] <=  8'h00;      memory[18985] <=  8'h00;      memory[18986] <=  8'h00;      memory[18987] <=  8'h00;      memory[18988] <=  8'h00;      memory[18989] <=  8'h00;      memory[18990] <=  8'h00;      memory[18991] <=  8'h00;      memory[18992] <=  8'h00;      memory[18993] <=  8'h00;      memory[18994] <=  8'h00;      memory[18995] <=  8'h00;      memory[18996] <=  8'h00;      memory[18997] <=  8'h00;      memory[18998] <=  8'h00;      memory[18999] <=  8'h00;      memory[19000] <=  8'h00;      memory[19001] <=  8'h00;      memory[19002] <=  8'h00;      memory[19003] <=  8'h00;      memory[19004] <=  8'h00;      memory[19005] <=  8'h00;      memory[19006] <=  8'h00;      memory[19007] <=  8'h00;      memory[19008] <=  8'h00;      memory[19009] <=  8'h00;      memory[19010] <=  8'h00;      memory[19011] <=  8'h00;      memory[19012] <=  8'h00;      memory[19013] <=  8'h00;      memory[19014] <=  8'h00;      memory[19015] <=  8'h00;      memory[19016] <=  8'h00;      memory[19017] <=  8'h00;      memory[19018] <=  8'h00;      memory[19019] <=  8'h00;      memory[19020] <=  8'h00;      memory[19021] <=  8'h00;      memory[19022] <=  8'h00;      memory[19023] <=  8'h00;      memory[19024] <=  8'h00;      memory[19025] <=  8'h00;      memory[19026] <=  8'h00;      memory[19027] <=  8'h00;      memory[19028] <=  8'h00;      memory[19029] <=  8'h00;      memory[19030] <=  8'h00;      memory[19031] <=  8'h00;      memory[19032] <=  8'h00;      memory[19033] <=  8'h00;      memory[19034] <=  8'h00;      memory[19035] <=  8'h00;      memory[19036] <=  8'h00;      memory[19037] <=  8'h00;      memory[19038] <=  8'h00;      memory[19039] <=  8'h00;      memory[19040] <=  8'h00;      memory[19041] <=  8'h00;      memory[19042] <=  8'h00;      memory[19043] <=  8'h00;      memory[19044] <=  8'h00;      memory[19045] <=  8'h00;      memory[19046] <=  8'h00;      memory[19047] <=  8'h00;      memory[19048] <=  8'h00;      memory[19049] <=  8'h00;      memory[19050] <=  8'h00;      memory[19051] <=  8'h00;      memory[19052] <=  8'h00;      memory[19053] <=  8'h00;      memory[19054] <=  8'h00;      memory[19055] <=  8'h00;      memory[19056] <=  8'h00;      memory[19057] <=  8'h00;      memory[19058] <=  8'h00;      memory[19059] <=  8'h00;      memory[19060] <=  8'h00;      memory[19061] <=  8'h00;      memory[19062] <=  8'h00;      memory[19063] <=  8'h00;      memory[19064] <=  8'h00;      memory[19065] <=  8'h00;      memory[19066] <=  8'h00;      memory[19067] <=  8'h00;      memory[19068] <=  8'h00;      memory[19069] <=  8'h00;      memory[19070] <=  8'h00;      memory[19071] <=  8'h00;      memory[19072] <=  8'h00;      memory[19073] <=  8'h00;      memory[19074] <=  8'h00;      memory[19075] <=  8'h00;      memory[19076] <=  8'h00;      memory[19077] <=  8'h00;      memory[19078] <=  8'h00;      memory[19079] <=  8'h00;      memory[19080] <=  8'h00;      memory[19081] <=  8'h00;      memory[19082] <=  8'h00;      memory[19083] <=  8'h00;      memory[19084] <=  8'h00;      memory[19085] <=  8'h00;      memory[19086] <=  8'h00;      memory[19087] <=  8'h00;      memory[19088] <=  8'h00;      memory[19089] <=  8'h00;      memory[19090] <=  8'h00;      memory[19091] <=  8'h00;      memory[19092] <=  8'h00;      memory[19093] <=  8'h00;      memory[19094] <=  8'h00;      memory[19095] <=  8'h00;      memory[19096] <=  8'h00;      memory[19097] <=  8'h00;      memory[19098] <=  8'h00;      memory[19099] <=  8'h00;      memory[19100] <=  8'h00;      memory[19101] <=  8'h00;      memory[19102] <=  8'h00;      memory[19103] <=  8'h00;      memory[19104] <=  8'h00;      memory[19105] <=  8'h00;      memory[19106] <=  8'h00;      memory[19107] <=  8'h00;      memory[19108] <=  8'h00;      memory[19109] <=  8'h00;      memory[19110] <=  8'h00;      memory[19111] <=  8'h00;      memory[19112] <=  8'h00;      memory[19113] <=  8'h00;      memory[19114] <=  8'h00;      memory[19115] <=  8'h00;      memory[19116] <=  8'h00;      memory[19117] <=  8'h00;      memory[19118] <=  8'h00;      memory[19119] <=  8'h00;      memory[19120] <=  8'h00;      memory[19121] <=  8'h00;      memory[19122] <=  8'h00;      memory[19123] <=  8'h00;      memory[19124] <=  8'h00;      memory[19125] <=  8'h00;      memory[19126] <=  8'h00;      memory[19127] <=  8'h00;      memory[19128] <=  8'h00;      memory[19129] <=  8'h00;      memory[19130] <=  8'h00;      memory[19131] <=  8'h00;      memory[19132] <=  8'h00;      memory[19133] <=  8'h00;      memory[19134] <=  8'h00;      memory[19135] <=  8'h00;      memory[19136] <=  8'h00;      memory[19137] <=  8'h00;      memory[19138] <=  8'h00;      memory[19139] <=  8'h00;      memory[19140] <=  8'h00;      memory[19141] <=  8'h00;      memory[19142] <=  8'h00;      memory[19143] <=  8'h00;      memory[19144] <=  8'h00;      memory[19145] <=  8'h00;      memory[19146] <=  8'h00;      memory[19147] <=  8'h00;      memory[19148] <=  8'h00;      memory[19149] <=  8'h00;      memory[19150] <=  8'h00;      memory[19151] <=  8'h00;      memory[19152] <=  8'h00;      memory[19153] <=  8'h00;      memory[19154] <=  8'h00;      memory[19155] <=  8'h00;      memory[19156] <=  8'h00;      memory[19157] <=  8'h00;      memory[19158] <=  8'h00;      memory[19159] <=  8'h00;      memory[19160] <=  8'h00;      memory[19161] <=  8'h00;      memory[19162] <=  8'h00;      memory[19163] <=  8'h00;      memory[19164] <=  8'h00;      memory[19165] <=  8'h00;      memory[19166] <=  8'h00;      memory[19167] <=  8'h00;      memory[19168] <=  8'h00;      memory[19169] <=  8'h00;      memory[19170] <=  8'h00;      memory[19171] <=  8'h00;      memory[19172] <=  8'h00;      memory[19173] <=  8'h00;      memory[19174] <=  8'h00;      memory[19175] <=  8'h00;      memory[19176] <=  8'h00;      memory[19177] <=  8'h00;      memory[19178] <=  8'h00;      memory[19179] <=  8'h00;      memory[19180] <=  8'h00;      memory[19181] <=  8'h00;      memory[19182] <=  8'h00;      memory[19183] <=  8'h00;      memory[19184] <=  8'h00;      memory[19185] <=  8'h00;      memory[19186] <=  8'h00;      memory[19187] <=  8'h00;      memory[19188] <=  8'h00;      memory[19189] <=  8'h00;      memory[19190] <=  8'h00;      memory[19191] <=  8'h00;      memory[19192] <=  8'h00;      memory[19193] <=  8'h00;      memory[19194] <=  8'h00;      memory[19195] <=  8'h00;      memory[19196] <=  8'h00;      memory[19197] <=  8'h00;      memory[19198] <=  8'h00;      memory[19199] <=  8'h00;      memory[19200] <=  8'h00;      memory[19201] <=  8'h00;      memory[19202] <=  8'h00;      memory[19203] <=  8'h00;      memory[19204] <=  8'h00;      memory[19205] <=  8'h00;      memory[19206] <=  8'h00;      memory[19207] <=  8'h00;      memory[19208] <=  8'h00;      memory[19209] <=  8'h00;      memory[19210] <=  8'h00;      memory[19211] <=  8'h00;      memory[19212] <=  8'h00;      memory[19213] <=  8'h00;      memory[19214] <=  8'h00;      memory[19215] <=  8'h00;      memory[19216] <=  8'h00;      memory[19217] <=  8'h00;      memory[19218] <=  8'h00;      memory[19219] <=  8'h00;      memory[19220] <=  8'h00;      memory[19221] <=  8'h00;      memory[19222] <=  8'h00;      memory[19223] <=  8'h00;      memory[19224] <=  8'h00;      memory[19225] <=  8'h00;      memory[19226] <=  8'h00;      memory[19227] <=  8'h00;      memory[19228] <=  8'h00;      memory[19229] <=  8'h00;      memory[19230] <=  8'h00;      memory[19231] <=  8'h00;      memory[19232] <=  8'h00;      memory[19233] <=  8'h00;      memory[19234] <=  8'h00;      memory[19235] <=  8'h00;      memory[19236] <=  8'h00;      memory[19237] <=  8'h00;      memory[19238] <=  8'h00;      memory[19239] <=  8'h00;      memory[19240] <=  8'h00;      memory[19241] <=  8'h00;      memory[19242] <=  8'h00;      memory[19243] <=  8'h00;      memory[19244] <=  8'h00;      memory[19245] <=  8'h00;      memory[19246] <=  8'h00;      memory[19247] <=  8'h00;      memory[19248] <=  8'h00;      memory[19249] <=  8'h00;      memory[19250] <=  8'h00;      memory[19251] <=  8'h00;      memory[19252] <=  8'h00;      memory[19253] <=  8'h00;      memory[19254] <=  8'h00;      memory[19255] <=  8'h00;      memory[19256] <=  8'h00;      memory[19257] <=  8'h00;      memory[19258] <=  8'h00;      memory[19259] <=  8'h00;      memory[19260] <=  8'h00;      memory[19261] <=  8'h00;      memory[19262] <=  8'h00;      memory[19263] <=  8'h00;      memory[19264] <=  8'h00;      memory[19265] <=  8'h00;      memory[19266] <=  8'h00;      memory[19267] <=  8'h00;      memory[19268] <=  8'h00;      memory[19269] <=  8'h00;      memory[19270] <=  8'h00;      memory[19271] <=  8'h00;      memory[19272] <=  8'h00;      memory[19273] <=  8'h00;      memory[19274] <=  8'h00;      memory[19275] <=  8'h00;      memory[19276] <=  8'h00;      memory[19277] <=  8'h00;      memory[19278] <=  8'h00;      memory[19279] <=  8'h00;      memory[19280] <=  8'h00;      memory[19281] <=  8'h00;      memory[19282] <=  8'h00;      memory[19283] <=  8'h00;      memory[19284] <=  8'h00;      memory[19285] <=  8'h00;      memory[19286] <=  8'h00;      memory[19287] <=  8'h00;      memory[19288] <=  8'h00;      memory[19289] <=  8'h00;      memory[19290] <=  8'h00;      memory[19291] <=  8'h00;      memory[19292] <=  8'h00;      memory[19293] <=  8'h00;      memory[19294] <=  8'h00;      memory[19295] <=  8'h00;      memory[19296] <=  8'h00;      memory[19297] <=  8'h00;      memory[19298] <=  8'h00;      memory[19299] <=  8'h00;      memory[19300] <=  8'h00;      memory[19301] <=  8'h00;      memory[19302] <=  8'h00;      memory[19303] <=  8'h00;      memory[19304] <=  8'h00;      memory[19305] <=  8'h00;      memory[19306] <=  8'h00;      memory[19307] <=  8'h00;      memory[19308] <=  8'h00;      memory[19309] <=  8'h00;      memory[19310] <=  8'h00;      memory[19311] <=  8'h00;      memory[19312] <=  8'h00;      memory[19313] <=  8'h00;      memory[19314] <=  8'h00;      memory[19315] <=  8'h00;      memory[19316] <=  8'h00;      memory[19317] <=  8'h00;      memory[19318] <=  8'h00;      memory[19319] <=  8'h00;      memory[19320] <=  8'h00;      memory[19321] <=  8'h00;      memory[19322] <=  8'h00;      memory[19323] <=  8'h00;      memory[19324] <=  8'h00;      memory[19325] <=  8'h00;      memory[19326] <=  8'h00;      memory[19327] <=  8'h00;      memory[19328] <=  8'h00;      memory[19329] <=  8'h00;      memory[19330] <=  8'h00;      memory[19331] <=  8'h00;      memory[19332] <=  8'h00;      memory[19333] <=  8'h00;      memory[19334] <=  8'h00;      memory[19335] <=  8'h00;      memory[19336] <=  8'h00;      memory[19337] <=  8'h00;      memory[19338] <=  8'h00;      memory[19339] <=  8'h00;      memory[19340] <=  8'h00;      memory[19341] <=  8'h00;      memory[19342] <=  8'h00;      memory[19343] <=  8'h00;      memory[19344] <=  8'h00;      memory[19345] <=  8'h00;      memory[19346] <=  8'h00;      memory[19347] <=  8'h00;      memory[19348] <=  8'h00;      memory[19349] <=  8'h00;      memory[19350] <=  8'h00;      memory[19351] <=  8'h00;      memory[19352] <=  8'h00;      memory[19353] <=  8'h00;      memory[19354] <=  8'h00;      memory[19355] <=  8'h00;      memory[19356] <=  8'h00;      memory[19357] <=  8'h00;      memory[19358] <=  8'h00;      memory[19359] <=  8'h00;      memory[19360] <=  8'h00;      memory[19361] <=  8'h00;      memory[19362] <=  8'h00;      memory[19363] <=  8'h00;      memory[19364] <=  8'h00;      memory[19365] <=  8'h00;      memory[19366] <=  8'h00;      memory[19367] <=  8'h00;      memory[19368] <=  8'h00;      memory[19369] <=  8'h00;      memory[19370] <=  8'h00;      memory[19371] <=  8'h00;      memory[19372] <=  8'h00;      memory[19373] <=  8'h00;      memory[19374] <=  8'h00;      memory[19375] <=  8'h00;      memory[19376] <=  8'h00;      memory[19377] <=  8'h00;      memory[19378] <=  8'h00;      memory[19379] <=  8'h00;      memory[19380] <=  8'h00;      memory[19381] <=  8'h00;      memory[19382] <=  8'h00;      memory[19383] <=  8'h00;      memory[19384] <=  8'h00;      memory[19385] <=  8'h00;      memory[19386] <=  8'h00;      memory[19387] <=  8'h00;      memory[19388] <=  8'h00;      memory[19389] <=  8'h00;      memory[19390] <=  8'h00;      memory[19391] <=  8'h00;      memory[19392] <=  8'h00;      memory[19393] <=  8'h00;      memory[19394] <=  8'h00;      memory[19395] <=  8'h00;      memory[19396] <=  8'h00;      memory[19397] <=  8'h00;      memory[19398] <=  8'h00;      memory[19399] <=  8'h00;      memory[19400] <=  8'h00;      memory[19401] <=  8'h00;      memory[19402] <=  8'h00;      memory[19403] <=  8'h00;      memory[19404] <=  8'h00;      memory[19405] <=  8'h00;      memory[19406] <=  8'h00;      memory[19407] <=  8'h00;      memory[19408] <=  8'h00;      memory[19409] <=  8'h00;      memory[19410] <=  8'h00;      memory[19411] <=  8'h00;      memory[19412] <=  8'h00;      memory[19413] <=  8'h00;      memory[19414] <=  8'h00;      memory[19415] <=  8'h00;      memory[19416] <=  8'h00;      memory[19417] <=  8'h00;      memory[19418] <=  8'h00;      memory[19419] <=  8'h00;      memory[19420] <=  8'h00;      memory[19421] <=  8'h00;      memory[19422] <=  8'h00;      memory[19423] <=  8'h00;      memory[19424] <=  8'h00;      memory[19425] <=  8'h00;      memory[19426] <=  8'h00;      memory[19427] <=  8'h00;      memory[19428] <=  8'h00;      memory[19429] <=  8'h00;      memory[19430] <=  8'h00;      memory[19431] <=  8'h00;      memory[19432] <=  8'h00;      memory[19433] <=  8'h00;      memory[19434] <=  8'h00;      memory[19435] <=  8'h00;      memory[19436] <=  8'h00;      memory[19437] <=  8'h00;      memory[19438] <=  8'h00;      memory[19439] <=  8'h00;      memory[19440] <=  8'h00;      memory[19441] <=  8'h00;      memory[19442] <=  8'h00;      memory[19443] <=  8'h00;      memory[19444] <=  8'h00;      memory[19445] <=  8'h00;      memory[19446] <=  8'h00;      memory[19447] <=  8'h00;      memory[19448] <=  8'h00;      memory[19449] <=  8'h00;      memory[19450] <=  8'h00;      memory[19451] <=  8'h00;      memory[19452] <=  8'h00;      memory[19453] <=  8'h00;      memory[19454] <=  8'h00;      memory[19455] <=  8'h00;      memory[19456] <=  8'h00;      memory[19457] <=  8'h00;      memory[19458] <=  8'h00;      memory[19459] <=  8'h00;      memory[19460] <=  8'h00;      memory[19461] <=  8'h00;      memory[19462] <=  8'h00;      memory[19463] <=  8'h00;      memory[19464] <=  8'h00;      memory[19465] <=  8'h00;      memory[19466] <=  8'h00;      memory[19467] <=  8'h00;      memory[19468] <=  8'h00;      memory[19469] <=  8'h00;      memory[19470] <=  8'h00;      memory[19471] <=  8'h00;      memory[19472] <=  8'h00;      memory[19473] <=  8'h00;      memory[19474] <=  8'h00;      memory[19475] <=  8'h00;      memory[19476] <=  8'h00;      memory[19477] <=  8'h00;      memory[19478] <=  8'h00;      memory[19479] <=  8'h00;      memory[19480] <=  8'h00;      memory[19481] <=  8'h00;      memory[19482] <=  8'h00;      memory[19483] <=  8'h00;      memory[19484] <=  8'h00;      memory[19485] <=  8'h00;      memory[19486] <=  8'h00;      memory[19487] <=  8'h00;      memory[19488] <=  8'h00;      memory[19489] <=  8'h00;      memory[19490] <=  8'h00;      memory[19491] <=  8'h00;      memory[19492] <=  8'h00;      memory[19493] <=  8'h00;      memory[19494] <=  8'h00;      memory[19495] <=  8'h00;      memory[19496] <=  8'h00;      memory[19497] <=  8'h00;      memory[19498] <=  8'h00;      memory[19499] <=  8'h00;      memory[19500] <=  8'h00;      memory[19501] <=  8'h00;      memory[19502] <=  8'h00;      memory[19503] <=  8'h00;      memory[19504] <=  8'h00;      memory[19505] <=  8'h00;      memory[19506] <=  8'h00;      memory[19507] <=  8'h00;      memory[19508] <=  8'h00;      memory[19509] <=  8'h00;      memory[19510] <=  8'h00;      memory[19511] <=  8'h00;      memory[19512] <=  8'h00;      memory[19513] <=  8'h00;      memory[19514] <=  8'h00;      memory[19515] <=  8'h00;      memory[19516] <=  8'h00;      memory[19517] <=  8'h00;      memory[19518] <=  8'h00;      memory[19519] <=  8'h00;      memory[19520] <=  8'h00;      memory[19521] <=  8'h00;      memory[19522] <=  8'h00;      memory[19523] <=  8'h00;      memory[19524] <=  8'h00;      memory[19525] <=  8'h00;      memory[19526] <=  8'h00;      memory[19527] <=  8'h00;      memory[19528] <=  8'h00;      memory[19529] <=  8'h00;      memory[19530] <=  8'h00;      memory[19531] <=  8'h00;      memory[19532] <=  8'h00;      memory[19533] <=  8'h00;      memory[19534] <=  8'h00;      memory[19535] <=  8'h00;      memory[19536] <=  8'h00;      memory[19537] <=  8'h00;      memory[19538] <=  8'h00;      memory[19539] <=  8'h00;      memory[19540] <=  8'h00;      memory[19541] <=  8'h00;      memory[19542] <=  8'h00;      memory[19543] <=  8'h00;      memory[19544] <=  8'h00;      memory[19545] <=  8'h00;      memory[19546] <=  8'h00;      memory[19547] <=  8'h00;      memory[19548] <=  8'h00;      memory[19549] <=  8'h00;      memory[19550] <=  8'h00;      memory[19551] <=  8'h00;      memory[19552] <=  8'h00;      memory[19553] <=  8'h00;      memory[19554] <=  8'h00;      memory[19555] <=  8'h00;      memory[19556] <=  8'h00;      memory[19557] <=  8'h00;      memory[19558] <=  8'h00;      memory[19559] <=  8'h00;      memory[19560] <=  8'h00;      memory[19561] <=  8'h00;      memory[19562] <=  8'h00;      memory[19563] <=  8'h00;      memory[19564] <=  8'h00;      memory[19565] <=  8'h00;      memory[19566] <=  8'h00;      memory[19567] <=  8'h00;      memory[19568] <=  8'h00;      memory[19569] <=  8'h00;      memory[19570] <=  8'h00;      memory[19571] <=  8'h00;      memory[19572] <=  8'h00;      memory[19573] <=  8'h00;      memory[19574] <=  8'h00;      memory[19575] <=  8'h00;      memory[19576] <=  8'h00;      memory[19577] <=  8'h00;      memory[19578] <=  8'h00;      memory[19579] <=  8'h00;      memory[19580] <=  8'h00;      memory[19581] <=  8'h00;      memory[19582] <=  8'h00;      memory[19583] <=  8'h00;      memory[19584] <=  8'h00;      memory[19585] <=  8'h00;      memory[19586] <=  8'h00;      memory[19587] <=  8'h00;      memory[19588] <=  8'h00;      memory[19589] <=  8'h00;      memory[19590] <=  8'h00;      memory[19591] <=  8'h00;      memory[19592] <=  8'h00;      memory[19593] <=  8'h00;      memory[19594] <=  8'h00;      memory[19595] <=  8'h00;      memory[19596] <=  8'h00;      memory[19597] <=  8'h00;      memory[19598] <=  8'h00;      memory[19599] <=  8'h00;      memory[19600] <=  8'h00;      memory[19601] <=  8'h00;      memory[19602] <=  8'h00;      memory[19603] <=  8'h00;      memory[19604] <=  8'h00;      memory[19605] <=  8'h00;      memory[19606] <=  8'h00;      memory[19607] <=  8'h00;      memory[19608] <=  8'h00;      memory[19609] <=  8'h00;      memory[19610] <=  8'h00;      memory[19611] <=  8'h00;      memory[19612] <=  8'h00;      memory[19613] <=  8'h00;      memory[19614] <=  8'h00;      memory[19615] <=  8'h00;      memory[19616] <=  8'h00;      memory[19617] <=  8'h00;      memory[19618] <=  8'h00;      memory[19619] <=  8'h00;      memory[19620] <=  8'h00;      memory[19621] <=  8'h00;      memory[19622] <=  8'h00;      memory[19623] <=  8'h00;      memory[19624] <=  8'h00;      memory[19625] <=  8'h00;      memory[19626] <=  8'h00;      memory[19627] <=  8'h00;      memory[19628] <=  8'h00;      memory[19629] <=  8'h00;      memory[19630] <=  8'h00;      memory[19631] <=  8'h00;      memory[19632] <=  8'h00;      memory[19633] <=  8'h00;      memory[19634] <=  8'h00;      memory[19635] <=  8'h00;      memory[19636] <=  8'h00;      memory[19637] <=  8'h00;      memory[19638] <=  8'h00;      memory[19639] <=  8'h00;      memory[19640] <=  8'h00;      memory[19641] <=  8'h00;      memory[19642] <=  8'h00;      memory[19643] <=  8'h00;      memory[19644] <=  8'h00;      memory[19645] <=  8'h00;      memory[19646] <=  8'h00;      memory[19647] <=  8'h00;      memory[19648] <=  8'h00;      memory[19649] <=  8'h00;      memory[19650] <=  8'h00;      memory[19651] <=  8'h00;      memory[19652] <=  8'h00;      memory[19653] <=  8'h00;      memory[19654] <=  8'h00;      memory[19655] <=  8'h00;      memory[19656] <=  8'h00;      memory[19657] <=  8'h00;      memory[19658] <=  8'h00;      memory[19659] <=  8'h00;      memory[19660] <=  8'h00;      memory[19661] <=  8'h00;      memory[19662] <=  8'h00;      memory[19663] <=  8'h00;      memory[19664] <=  8'h00;      memory[19665] <=  8'h00;      memory[19666] <=  8'h00;      memory[19667] <=  8'h00;      memory[19668] <=  8'h00;      memory[19669] <=  8'h00;      memory[19670] <=  8'h00;      memory[19671] <=  8'h00;      memory[19672] <=  8'h00;      memory[19673] <=  8'h00;      memory[19674] <=  8'h00;      memory[19675] <=  8'h00;      memory[19676] <=  8'h00;      memory[19677] <=  8'h00;      memory[19678] <=  8'h00;      memory[19679] <=  8'h00;      memory[19680] <=  8'h00;      memory[19681] <=  8'h00;      memory[19682] <=  8'h00;      memory[19683] <=  8'h00;      memory[19684] <=  8'h00;      memory[19685] <=  8'h00;      memory[19686] <=  8'h00;      memory[19687] <=  8'h00;      memory[19688] <=  8'h00;      memory[19689] <=  8'h00;      memory[19690] <=  8'h00;      memory[19691] <=  8'h00;      memory[19692] <=  8'h00;      memory[19693] <=  8'h00;      memory[19694] <=  8'h00;      memory[19695] <=  8'h00;      memory[19696] <=  8'h00;      memory[19697] <=  8'h00;      memory[19698] <=  8'h00;      memory[19699] <=  8'h00;      memory[19700] <=  8'h00;      memory[19701] <=  8'h00;      memory[19702] <=  8'h00;      memory[19703] <=  8'h00;      memory[19704] <=  8'h00;      memory[19705] <=  8'h00;      memory[19706] <=  8'h00;      memory[19707] <=  8'h00;      memory[19708] <=  8'h00;      memory[19709] <=  8'h00;      memory[19710] <=  8'h00;      memory[19711] <=  8'h00;      memory[19712] <=  8'h00;      memory[19713] <=  8'h00;      memory[19714] <=  8'h00;      memory[19715] <=  8'h00;      memory[19716] <=  8'h00;      memory[19717] <=  8'h00;      memory[19718] <=  8'h00;      memory[19719] <=  8'h00;      memory[19720] <=  8'h00;      memory[19721] <=  8'h00;      memory[19722] <=  8'h00;      memory[19723] <=  8'h00;      memory[19724] <=  8'h00;      memory[19725] <=  8'h00;      memory[19726] <=  8'h00;      memory[19727] <=  8'h00;      memory[19728] <=  8'h00;      memory[19729] <=  8'h00;      memory[19730] <=  8'h00;      memory[19731] <=  8'h00;      memory[19732] <=  8'h00;      memory[19733] <=  8'h00;      memory[19734] <=  8'h00;      memory[19735] <=  8'h00;      memory[19736] <=  8'h00;      memory[19737] <=  8'h00;      memory[19738] <=  8'h00;      memory[19739] <=  8'h00;      memory[19740] <=  8'h00;      memory[19741] <=  8'h00;      memory[19742] <=  8'h00;      memory[19743] <=  8'h00;      memory[19744] <=  8'h00;      memory[19745] <=  8'h00;      memory[19746] <=  8'h00;      memory[19747] <=  8'h00;      memory[19748] <=  8'h00;      memory[19749] <=  8'h00;      memory[19750] <=  8'h00;      memory[19751] <=  8'h00;      memory[19752] <=  8'h00;      memory[19753] <=  8'h00;      memory[19754] <=  8'h00;      memory[19755] <=  8'h00;      memory[19756] <=  8'h00;      memory[19757] <=  8'h00;      memory[19758] <=  8'h00;      memory[19759] <=  8'h00;      memory[19760] <=  8'h00;      memory[19761] <=  8'h00;      memory[19762] <=  8'h00;      memory[19763] <=  8'h00;      memory[19764] <=  8'h00;      memory[19765] <=  8'h00;      memory[19766] <=  8'h00;      memory[19767] <=  8'h00;      memory[19768] <=  8'h00;      memory[19769] <=  8'h00;      memory[19770] <=  8'h00;      memory[19771] <=  8'h00;      memory[19772] <=  8'h00;      memory[19773] <=  8'h00;      memory[19774] <=  8'h00;      memory[19775] <=  8'h00;      memory[19776] <=  8'h00;      memory[19777] <=  8'h00;      memory[19778] <=  8'h00;      memory[19779] <=  8'h00;      memory[19780] <=  8'h00;      memory[19781] <=  8'h00;      memory[19782] <=  8'h00;      memory[19783] <=  8'h00;      memory[19784] <=  8'h00;      memory[19785] <=  8'h00;      memory[19786] <=  8'h00;      memory[19787] <=  8'h00;      memory[19788] <=  8'h00;      memory[19789] <=  8'h00;      memory[19790] <=  8'h00;      memory[19791] <=  8'h00;      memory[19792] <=  8'h00;      memory[19793] <=  8'h00;      memory[19794] <=  8'h00;      memory[19795] <=  8'h00;      memory[19796] <=  8'h00;      memory[19797] <=  8'h00;      memory[19798] <=  8'h00;      memory[19799] <=  8'h00;      memory[19800] <=  8'h00;      memory[19801] <=  8'h00;      memory[19802] <=  8'h00;      memory[19803] <=  8'h00;      memory[19804] <=  8'h00;      memory[19805] <=  8'h00;      memory[19806] <=  8'h00;      memory[19807] <=  8'h00;      memory[19808] <=  8'h00;      memory[19809] <=  8'h00;      memory[19810] <=  8'h00;      memory[19811] <=  8'h00;      memory[19812] <=  8'h00;      memory[19813] <=  8'h00;      memory[19814] <=  8'h00;      memory[19815] <=  8'h00;      memory[19816] <=  8'h00;      memory[19817] <=  8'h00;      memory[19818] <=  8'h00;      memory[19819] <=  8'h00;      memory[19820] <=  8'h00;      memory[19821] <=  8'h00;      memory[19822] <=  8'h00;      memory[19823] <=  8'h00;      memory[19824] <=  8'h00;      memory[19825] <=  8'h00;      memory[19826] <=  8'h00;      memory[19827] <=  8'h00;      memory[19828] <=  8'h00;      memory[19829] <=  8'h00;      memory[19830] <=  8'h00;      memory[19831] <=  8'h00;      memory[19832] <=  8'h00;      memory[19833] <=  8'h00;      memory[19834] <=  8'h00;      memory[19835] <=  8'h00;      memory[19836] <=  8'h00;      memory[19837] <=  8'h00;      memory[19838] <=  8'h00;      memory[19839] <=  8'h00;      memory[19840] <=  8'h00;      memory[19841] <=  8'h00;      memory[19842] <=  8'h00;      memory[19843] <=  8'h00;      memory[19844] <=  8'h00;      memory[19845] <=  8'h00;      memory[19846] <=  8'h00;      memory[19847] <=  8'h00;      memory[19848] <=  8'h00;      memory[19849] <=  8'h00;      memory[19850] <=  8'h00;      memory[19851] <=  8'h00;      memory[19852] <=  8'h00;      memory[19853] <=  8'h00;      memory[19854] <=  8'h00;      memory[19855] <=  8'h00;      memory[19856] <=  8'h00;      memory[19857] <=  8'h00;      memory[19858] <=  8'h00;      memory[19859] <=  8'h00;      memory[19860] <=  8'h00;      memory[19861] <=  8'h00;      memory[19862] <=  8'h00;      memory[19863] <=  8'h00;      memory[19864] <=  8'h00;      memory[19865] <=  8'h00;      memory[19866] <=  8'h00;      memory[19867] <=  8'h00;      memory[19868] <=  8'h00;      memory[19869] <=  8'h00;      memory[19870] <=  8'h00;      memory[19871] <=  8'h00;      memory[19872] <=  8'h00;      memory[19873] <=  8'h00;      memory[19874] <=  8'h00;      memory[19875] <=  8'h00;      memory[19876] <=  8'h00;      memory[19877] <=  8'h00;      memory[19878] <=  8'h00;      memory[19879] <=  8'h00;      memory[19880] <=  8'h00;      memory[19881] <=  8'h00;      memory[19882] <=  8'h00;      memory[19883] <=  8'h00;      memory[19884] <=  8'h00;      memory[19885] <=  8'h00;      memory[19886] <=  8'h00;      memory[19887] <=  8'h00;      memory[19888] <=  8'h00;      memory[19889] <=  8'h00;      memory[19890] <=  8'h00;      memory[19891] <=  8'h00;      memory[19892] <=  8'h00;      memory[19893] <=  8'h00;      memory[19894] <=  8'h00;      memory[19895] <=  8'h00;      memory[19896] <=  8'h00;      memory[19897] <=  8'h00;      memory[19898] <=  8'h00;      memory[19899] <=  8'h00;      memory[19900] <=  8'h00;      memory[19901] <=  8'h00;      memory[19902] <=  8'h00;      memory[19903] <=  8'h00;      memory[19904] <=  8'h00;      memory[19905] <=  8'h00;      memory[19906] <=  8'h00;      memory[19907] <=  8'h00;      memory[19908] <=  8'h00;      memory[19909] <=  8'h00;      memory[19910] <=  8'h00;      memory[19911] <=  8'h00;      memory[19912] <=  8'h00;      memory[19913] <=  8'h00;      memory[19914] <=  8'h00;      memory[19915] <=  8'h00;      memory[19916] <=  8'h00;      memory[19917] <=  8'h00;      memory[19918] <=  8'h00;      memory[19919] <=  8'h00;      memory[19920] <=  8'h00;      memory[19921] <=  8'h00;      memory[19922] <=  8'h00;      memory[19923] <=  8'h00;      memory[19924] <=  8'h00;      memory[19925] <=  8'h00;      memory[19926] <=  8'h00;      memory[19927] <=  8'h00;      memory[19928] <=  8'h00;      memory[19929] <=  8'h00;      memory[19930] <=  8'h00;      memory[19931] <=  8'h00;      memory[19932] <=  8'h00;      memory[19933] <=  8'h00;      memory[19934] <=  8'h00;      memory[19935] <=  8'h00;      memory[19936] <=  8'h00;      memory[19937] <=  8'h00;      memory[19938] <=  8'h00;      memory[19939] <=  8'h00;      memory[19940] <=  8'h00;      memory[19941] <=  8'h00;      memory[19942] <=  8'h00;      memory[19943] <=  8'h00;      memory[19944] <=  8'h00;      memory[19945] <=  8'h00;      memory[19946] <=  8'h00;      memory[19947] <=  8'h00;      memory[19948] <=  8'h00;      memory[19949] <=  8'h00;      memory[19950] <=  8'h00;      memory[19951] <=  8'h00;      memory[19952] <=  8'h00;      memory[19953] <=  8'h00;      memory[19954] <=  8'h00;      memory[19955] <=  8'h00;      memory[19956] <=  8'h00;      memory[19957] <=  8'h00;      memory[19958] <=  8'h00;      memory[19959] <=  8'h00;      memory[19960] <=  8'h00;      memory[19961] <=  8'h00;      memory[19962] <=  8'h00;      memory[19963] <=  8'h00;      memory[19964] <=  8'h00;      memory[19965] <=  8'h00;      memory[19966] <=  8'h00;      memory[19967] <=  8'h00;      memory[19968] <=  8'h00;      memory[19969] <=  8'h00;      memory[19970] <=  8'h00;      memory[19971] <=  8'h00;      memory[19972] <=  8'h00;      memory[19973] <=  8'h00;      memory[19974] <=  8'h00;      memory[19975] <=  8'h00;      memory[19976] <=  8'h00;      memory[19977] <=  8'h00;      memory[19978] <=  8'h00;      memory[19979] <=  8'h00;      memory[19980] <=  8'h00;      memory[19981] <=  8'h00;      memory[19982] <=  8'h00;      memory[19983] <=  8'h00;      memory[19984] <=  8'h00;      memory[19985] <=  8'h00;      memory[19986] <=  8'h00;      memory[19987] <=  8'h00;      memory[19988] <=  8'h00;      memory[19989] <=  8'h00;      memory[19990] <=  8'h00;      memory[19991] <=  8'h00;      memory[19992] <=  8'h00;      memory[19993] <=  8'h00;      memory[19994] <=  8'h00;      memory[19995] <=  8'h00;      memory[19996] <=  8'h00;      memory[19997] <=  8'h00;      memory[19998] <=  8'h00;      memory[19999] <=  8'h00;      memory[20000] <=  8'h00;      memory[20001] <=  8'h00;      memory[20002] <=  8'h00;      memory[20003] <=  8'h00;      memory[20004] <=  8'h00;      memory[20005] <=  8'h00;      memory[20006] <=  8'h00;      memory[20007] <=  8'h00;      memory[20008] <=  8'h00;      memory[20009] <=  8'h00;      memory[20010] <=  8'h00;      memory[20011] <=  8'h00;      memory[20012] <=  8'h00;      memory[20013] <=  8'h00;      memory[20014] <=  8'h00;      memory[20015] <=  8'h00;      memory[20016] <=  8'h00;      memory[20017] <=  8'h00;      memory[20018] <=  8'h00;      memory[20019] <=  8'h00;      memory[20020] <=  8'h00;      memory[20021] <=  8'h00;      memory[20022] <=  8'h00;      memory[20023] <=  8'h00;      memory[20024] <=  8'h00;      memory[20025] <=  8'h00;      memory[20026] <=  8'h00;      memory[20027] <=  8'h00;      memory[20028] <=  8'h00;      memory[20029] <=  8'h00;      memory[20030] <=  8'h00;      memory[20031] <=  8'h00;      memory[20032] <=  8'h00;      memory[20033] <=  8'h00;      memory[20034] <=  8'h00;      memory[20035] <=  8'h00;      memory[20036] <=  8'h00;      memory[20037] <=  8'h00;      memory[20038] <=  8'h00;      memory[20039] <=  8'h00;      memory[20040] <=  8'h00;      memory[20041] <=  8'h00;      memory[20042] <=  8'h00;      memory[20043] <=  8'h00;      memory[20044] <=  8'h00;      memory[20045] <=  8'h00;      memory[20046] <=  8'h00;      memory[20047] <=  8'h00;      memory[20048] <=  8'h00;      memory[20049] <=  8'h00;      memory[20050] <=  8'h00;      memory[20051] <=  8'h00;      memory[20052] <=  8'h00;      memory[20053] <=  8'h00;      memory[20054] <=  8'h00;      memory[20055] <=  8'h00;      memory[20056] <=  8'h00;      memory[20057] <=  8'h00;      memory[20058] <=  8'h00;      memory[20059] <=  8'h00;      memory[20060] <=  8'h00;      memory[20061] <=  8'h00;      memory[20062] <=  8'h00;      memory[20063] <=  8'h00;      memory[20064] <=  8'h00;      memory[20065] <=  8'h00;      memory[20066] <=  8'h00;      memory[20067] <=  8'h00;      memory[20068] <=  8'h00;      memory[20069] <=  8'h00;      memory[20070] <=  8'h00;      memory[20071] <=  8'h00;      memory[20072] <=  8'h00;      memory[20073] <=  8'h00;      memory[20074] <=  8'h00;      memory[20075] <=  8'h00;      memory[20076] <=  8'h00;      memory[20077] <=  8'h00;      memory[20078] <=  8'h00;      memory[20079] <=  8'h00;      memory[20080] <=  8'h00;      memory[20081] <=  8'h00;      memory[20082] <=  8'h00;      memory[20083] <=  8'h00;      memory[20084] <=  8'h00;      memory[20085] <=  8'h00;      memory[20086] <=  8'h00;      memory[20087] <=  8'h00;      memory[20088] <=  8'h00;      memory[20089] <=  8'h00;      memory[20090] <=  8'h00;      memory[20091] <=  8'h00;      memory[20092] <=  8'h00;      memory[20093] <=  8'h00;      memory[20094] <=  8'h00;      memory[20095] <=  8'h00;      memory[20096] <=  8'h00;      memory[20097] <=  8'h00;      memory[20098] <=  8'h00;      memory[20099] <=  8'h00;      memory[20100] <=  8'h00;      memory[20101] <=  8'h00;      memory[20102] <=  8'h00;      memory[20103] <=  8'h00;      memory[20104] <=  8'h00;      memory[20105] <=  8'h00;      memory[20106] <=  8'h00;      memory[20107] <=  8'h00;      memory[20108] <=  8'h00;      memory[20109] <=  8'h00;      memory[20110] <=  8'h00;      memory[20111] <=  8'h00;      memory[20112] <=  8'h00;      memory[20113] <=  8'h00;      memory[20114] <=  8'h00;      memory[20115] <=  8'h00;      memory[20116] <=  8'h00;      memory[20117] <=  8'h00;      memory[20118] <=  8'h00;      memory[20119] <=  8'h00;      memory[20120] <=  8'h00;      memory[20121] <=  8'h00;      memory[20122] <=  8'h00;      memory[20123] <=  8'h00;      memory[20124] <=  8'h00;      memory[20125] <=  8'h00;      memory[20126] <=  8'h00;      memory[20127] <=  8'h00;      memory[20128] <=  8'h00;      memory[20129] <=  8'h00;      memory[20130] <=  8'h00;      memory[20131] <=  8'h00;      memory[20132] <=  8'h00;      memory[20133] <=  8'h00;      memory[20134] <=  8'h00;      memory[20135] <=  8'h00;      memory[20136] <=  8'h00;      memory[20137] <=  8'h00;      memory[20138] <=  8'h00;      memory[20139] <=  8'h00;      memory[20140] <=  8'h00;      memory[20141] <=  8'h00;      memory[20142] <=  8'h00;      memory[20143] <=  8'h00;      memory[20144] <=  8'h00;      memory[20145] <=  8'h00;      memory[20146] <=  8'h00;      memory[20147] <=  8'h00;      memory[20148] <=  8'h00;      memory[20149] <=  8'h00;      memory[20150] <=  8'h00;      memory[20151] <=  8'h00;      memory[20152] <=  8'h00;      memory[20153] <=  8'h00;      memory[20154] <=  8'h00;      memory[20155] <=  8'h00;      memory[20156] <=  8'h00;      memory[20157] <=  8'h00;      memory[20158] <=  8'h00;      memory[20159] <=  8'h00;      memory[20160] <=  8'h00;      memory[20161] <=  8'h00;      memory[20162] <=  8'h00;      memory[20163] <=  8'h00;      memory[20164] <=  8'h00;      memory[20165] <=  8'h00;      memory[20166] <=  8'h00;      memory[20167] <=  8'h00;      memory[20168] <=  8'h00;      memory[20169] <=  8'h00;      memory[20170] <=  8'h00;      memory[20171] <=  8'h00;      memory[20172] <=  8'h00;      memory[20173] <=  8'h00;      memory[20174] <=  8'h00;      memory[20175] <=  8'h00;      memory[20176] <=  8'h00;      memory[20177] <=  8'h00;      memory[20178] <=  8'h00;      memory[20179] <=  8'h00;      memory[20180] <=  8'h00;      memory[20181] <=  8'h00;      memory[20182] <=  8'h00;      memory[20183] <=  8'h00;      memory[20184] <=  8'h00;      memory[20185] <=  8'h00;      memory[20186] <=  8'h00;      memory[20187] <=  8'h00;      memory[20188] <=  8'h00;      memory[20189] <=  8'h00;      memory[20190] <=  8'h00;      memory[20191] <=  8'h00;      memory[20192] <=  8'h00;      memory[20193] <=  8'h00;      memory[20194] <=  8'h00;      memory[20195] <=  8'h00;      memory[20196] <=  8'h00;      memory[20197] <=  8'h00;      memory[20198] <=  8'h00;      memory[20199] <=  8'h00;      memory[20200] <=  8'h00;      memory[20201] <=  8'h00;      memory[20202] <=  8'h00;      memory[20203] <=  8'h00;      memory[20204] <=  8'h00;      memory[20205] <=  8'h00;      memory[20206] <=  8'h00;      memory[20207] <=  8'h00;      memory[20208] <=  8'h00;      memory[20209] <=  8'h00;      memory[20210] <=  8'h00;      memory[20211] <=  8'h00;      memory[20212] <=  8'h00;      memory[20213] <=  8'h00;      memory[20214] <=  8'h00;      memory[20215] <=  8'h00;      memory[20216] <=  8'h00;      memory[20217] <=  8'h00;      memory[20218] <=  8'h00;      memory[20219] <=  8'h00;      memory[20220] <=  8'h00;      memory[20221] <=  8'h00;      memory[20222] <=  8'h00;      memory[20223] <=  8'h00;      memory[20224] <=  8'h00;      memory[20225] <=  8'h00;      memory[20226] <=  8'h00;      memory[20227] <=  8'h00;      memory[20228] <=  8'h00;      memory[20229] <=  8'h00;      memory[20230] <=  8'h00;      memory[20231] <=  8'h00;      memory[20232] <=  8'h00;      memory[20233] <=  8'h00;      memory[20234] <=  8'h00;      memory[20235] <=  8'h00;      memory[20236] <=  8'h00;      memory[20237] <=  8'h00;      memory[20238] <=  8'h00;      memory[20239] <=  8'h00;      memory[20240] <=  8'h00;      memory[20241] <=  8'h00;      memory[20242] <=  8'h00;      memory[20243] <=  8'h00;      memory[20244] <=  8'h00;      memory[20245] <=  8'h00;      memory[20246] <=  8'h00;      memory[20247] <=  8'h00;      memory[20248] <=  8'h00;      memory[20249] <=  8'h00;      memory[20250] <=  8'h00;      memory[20251] <=  8'h00;      memory[20252] <=  8'h00;      memory[20253] <=  8'h00;      memory[20254] <=  8'h00;      memory[20255] <=  8'h00;      memory[20256] <=  8'h00;      memory[20257] <=  8'h00;      memory[20258] <=  8'h00;      memory[20259] <=  8'h00;      memory[20260] <=  8'h00;      memory[20261] <=  8'h00;      memory[20262] <=  8'h00;      memory[20263] <=  8'h00;      memory[20264] <=  8'h00;      memory[20265] <=  8'h00;      memory[20266] <=  8'h00;      memory[20267] <=  8'h00;      memory[20268] <=  8'h00;      memory[20269] <=  8'h00;      memory[20270] <=  8'h00;      memory[20271] <=  8'h00;      memory[20272] <=  8'h00;      memory[20273] <=  8'h00;      memory[20274] <=  8'h00;      memory[20275] <=  8'h00;      memory[20276] <=  8'h00;      memory[20277] <=  8'h00;      memory[20278] <=  8'h00;      memory[20279] <=  8'h00;      memory[20280] <=  8'h00;      memory[20281] <=  8'h00;      memory[20282] <=  8'h00;      memory[20283] <=  8'h00;      memory[20284] <=  8'h00;      memory[20285] <=  8'h00;      memory[20286] <=  8'h00;      memory[20287] <=  8'h00;      memory[20288] <=  8'h00;      memory[20289] <=  8'h00;      memory[20290] <=  8'h00;      memory[20291] <=  8'h00;      memory[20292] <=  8'h00;      memory[20293] <=  8'h00;      memory[20294] <=  8'h00;      memory[20295] <=  8'h00;      memory[20296] <=  8'h00;      memory[20297] <=  8'h00;      memory[20298] <=  8'h00;      memory[20299] <=  8'h00;      memory[20300] <=  8'h00;      memory[20301] <=  8'h00;      memory[20302] <=  8'h00;      memory[20303] <=  8'h00;      memory[20304] <=  8'h00;      memory[20305] <=  8'h00;      memory[20306] <=  8'h00;      memory[20307] <=  8'h00;      memory[20308] <=  8'h00;      memory[20309] <=  8'h00;      memory[20310] <=  8'h00;      memory[20311] <=  8'h00;      memory[20312] <=  8'h00;      memory[20313] <=  8'h00;      memory[20314] <=  8'h00;      memory[20315] <=  8'h00;      memory[20316] <=  8'h00;      memory[20317] <=  8'h00;      memory[20318] <=  8'h00;      memory[20319] <=  8'h00;      memory[20320] <=  8'h00;      memory[20321] <=  8'h00;      memory[20322] <=  8'h00;      memory[20323] <=  8'h00;      memory[20324] <=  8'h00;      memory[20325] <=  8'h00;      memory[20326] <=  8'h00;      memory[20327] <=  8'h00;      memory[20328] <=  8'h00;      memory[20329] <=  8'h00;      memory[20330] <=  8'h00;      memory[20331] <=  8'h00;      memory[20332] <=  8'h00;      memory[20333] <=  8'h00;      memory[20334] <=  8'h00;      memory[20335] <=  8'h00;      memory[20336] <=  8'h00;      memory[20337] <=  8'h00;      memory[20338] <=  8'h00;      memory[20339] <=  8'h00;      memory[20340] <=  8'h00;      memory[20341] <=  8'h00;      memory[20342] <=  8'h00;      memory[20343] <=  8'h00;      memory[20344] <=  8'h00;      memory[20345] <=  8'h00;      memory[20346] <=  8'h00;      memory[20347] <=  8'h00;      memory[20348] <=  8'h00;      memory[20349] <=  8'h00;      memory[20350] <=  8'h00;      memory[20351] <=  8'h00;      memory[20352] <=  8'h00;      memory[20353] <=  8'h00;      memory[20354] <=  8'h00;      memory[20355] <=  8'h00;      memory[20356] <=  8'h00;      memory[20357] <=  8'h00;      memory[20358] <=  8'h00;      memory[20359] <=  8'h00;      memory[20360] <=  8'h00;      memory[20361] <=  8'h00;      memory[20362] <=  8'h00;      memory[20363] <=  8'h00;      memory[20364] <=  8'h00;      memory[20365] <=  8'h00;      memory[20366] <=  8'h00;      memory[20367] <=  8'h00;      memory[20368] <=  8'h00;      memory[20369] <=  8'h00;      memory[20370] <=  8'h00;      memory[20371] <=  8'h00;      memory[20372] <=  8'h00;      memory[20373] <=  8'h00;      memory[20374] <=  8'h00;      memory[20375] <=  8'h00;      memory[20376] <=  8'h00;      memory[20377] <=  8'h00;      memory[20378] <=  8'h00;      memory[20379] <=  8'h00;      memory[20380] <=  8'h00;      memory[20381] <=  8'h00;      memory[20382] <=  8'h00;      memory[20383] <=  8'h00;      memory[20384] <=  8'h00;      memory[20385] <=  8'h00;      memory[20386] <=  8'h00;      memory[20387] <=  8'h00;      memory[20388] <=  8'h00;      memory[20389] <=  8'h00;      memory[20390] <=  8'h00;      memory[20391] <=  8'h00;      memory[20392] <=  8'h00;      memory[20393] <=  8'h00;      memory[20394] <=  8'h00;      memory[20395] <=  8'h00;      memory[20396] <=  8'h00;      memory[20397] <=  8'h00;      memory[20398] <=  8'h00;      memory[20399] <=  8'h00;      memory[20400] <=  8'h00;      memory[20401] <=  8'h00;      memory[20402] <=  8'h00;      memory[20403] <=  8'h00;      memory[20404] <=  8'h00;      memory[20405] <=  8'h00;      memory[20406] <=  8'h00;      memory[20407] <=  8'h00;      memory[20408] <=  8'h00;      memory[20409] <=  8'h00;      memory[20410] <=  8'h00;      memory[20411] <=  8'h00;      memory[20412] <=  8'h00;      memory[20413] <=  8'h00;      memory[20414] <=  8'h00;      memory[20415] <=  8'h00;      memory[20416] <=  8'h00;      memory[20417] <=  8'h00;      memory[20418] <=  8'h00;      memory[20419] <=  8'h00;      memory[20420] <=  8'h00;      memory[20421] <=  8'h00;      memory[20422] <=  8'h00;      memory[20423] <=  8'h00;      memory[20424] <=  8'h00;      memory[20425] <=  8'h00;      memory[20426] <=  8'h00;      memory[20427] <=  8'h00;      memory[20428] <=  8'h00;      memory[20429] <=  8'h00;      memory[20430] <=  8'h00;      memory[20431] <=  8'h00;      memory[20432] <=  8'h00;      memory[20433] <=  8'h00;      memory[20434] <=  8'h00;      memory[20435] <=  8'h00;      memory[20436] <=  8'h00;      memory[20437] <=  8'h00;      memory[20438] <=  8'h00;      memory[20439] <=  8'h00;      memory[20440] <=  8'h00;      memory[20441] <=  8'h00;      memory[20442] <=  8'h00;      memory[20443] <=  8'h00;      memory[20444] <=  8'h00;      memory[20445] <=  8'h00;      memory[20446] <=  8'h00;      memory[20447] <=  8'h00;      memory[20448] <=  8'h00;      memory[20449] <=  8'h00;      memory[20450] <=  8'h00;      memory[20451] <=  8'h00;      memory[20452] <=  8'h00;      memory[20453] <=  8'h00;      memory[20454] <=  8'h00;      memory[20455] <=  8'h00;      memory[20456] <=  8'h00;      memory[20457] <=  8'h00;      memory[20458] <=  8'h00;      memory[20459] <=  8'h00;      memory[20460] <=  8'h00;      memory[20461] <=  8'h00;      memory[20462] <=  8'h00;      memory[20463] <=  8'h00;      memory[20464] <=  8'h00;      memory[20465] <=  8'h00;      memory[20466] <=  8'h00;      memory[20467] <=  8'h00;      memory[20468] <=  8'h00;      memory[20469] <=  8'h00;      memory[20470] <=  8'h00;      memory[20471] <=  8'h00;      memory[20472] <=  8'h00;      memory[20473] <=  8'h00;      memory[20474] <=  8'h00;      memory[20475] <=  8'h00;      memory[20476] <=  8'h00;      memory[20477] <=  8'h00;      memory[20478] <=  8'h00;      memory[20479] <=  8'h00;      memory[20480] <=  8'h00;      memory[20481] <=  8'h00;      memory[20482] <=  8'h00;      memory[20483] <=  8'h00;      memory[20484] <=  8'h00;      memory[20485] <=  8'h00;      memory[20486] <=  8'h00;      memory[20487] <=  8'h00;      memory[20488] <=  8'h00;      memory[20489] <=  8'h00;      memory[20490] <=  8'h00;      memory[20491] <=  8'h00;      memory[20492] <=  8'h00;      memory[20493] <=  8'h00;      memory[20494] <=  8'h00;      memory[20495] <=  8'h00;      memory[20496] <=  8'h00;      memory[20497] <=  8'h00;      memory[20498] <=  8'h00;      memory[20499] <=  8'h00;      memory[20500] <=  8'h00;      memory[20501] <=  8'h00;      memory[20502] <=  8'h00;      memory[20503] <=  8'h00;      memory[20504] <=  8'h00;      memory[20505] <=  8'h00;      memory[20506] <=  8'h00;      memory[20507] <=  8'h00;      memory[20508] <=  8'h00;      memory[20509] <=  8'h00;      memory[20510] <=  8'h00;      memory[20511] <=  8'h00;      memory[20512] <=  8'h00;      memory[20513] <=  8'h00;      memory[20514] <=  8'h00;      memory[20515] <=  8'h00;      memory[20516] <=  8'h00;      memory[20517] <=  8'h00;      memory[20518] <=  8'h00;      memory[20519] <=  8'h00;      memory[20520] <=  8'h00;      memory[20521] <=  8'h00;      memory[20522] <=  8'h00;      memory[20523] <=  8'h00;      memory[20524] <=  8'h00;      memory[20525] <=  8'h00;      memory[20526] <=  8'h00;      memory[20527] <=  8'h00;      memory[20528] <=  8'h00;      memory[20529] <=  8'h00;      memory[20530] <=  8'h00;      memory[20531] <=  8'h00;      memory[20532] <=  8'h00;      memory[20533] <=  8'h00;      memory[20534] <=  8'h00;      memory[20535] <=  8'h00;      memory[20536] <=  8'h00;      memory[20537] <=  8'h00;      memory[20538] <=  8'h00;      memory[20539] <=  8'h00;      memory[20540] <=  8'h00;      memory[20541] <=  8'h00;      memory[20542] <=  8'h00;      memory[20543] <=  8'h00;      memory[20544] <=  8'h00;      memory[20545] <=  8'h00;      memory[20546] <=  8'h00;      memory[20547] <=  8'h00;      memory[20548] <=  8'h00;      memory[20549] <=  8'h00;      memory[20550] <=  8'h00;      memory[20551] <=  8'h00;      memory[20552] <=  8'h00;      memory[20553] <=  8'h00;      memory[20554] <=  8'h00;      memory[20555] <=  8'h00;      memory[20556] <=  8'h00;      memory[20557] <=  8'h00;      memory[20558] <=  8'h00;      memory[20559] <=  8'h00;      memory[20560] <=  8'h00;      memory[20561] <=  8'h00;      memory[20562] <=  8'h00;      memory[20563] <=  8'h00;      memory[20564] <=  8'h00;      memory[20565] <=  8'h00;      memory[20566] <=  8'h00;      memory[20567] <=  8'h00;      memory[20568] <=  8'h00;      memory[20569] <=  8'h00;      memory[20570] <=  8'h00;      memory[20571] <=  8'h00;      memory[20572] <=  8'h00;      memory[20573] <=  8'h00;      memory[20574] <=  8'h00;      memory[20575] <=  8'h00;      memory[20576] <=  8'h00;      memory[20577] <=  8'h00;      memory[20578] <=  8'h00;      memory[20579] <=  8'h00;      memory[20580] <=  8'h00;      memory[20581] <=  8'h00;      memory[20582] <=  8'h00;      memory[20583] <=  8'h00;      memory[20584] <=  8'h00;      memory[20585] <=  8'h00;      memory[20586] <=  8'h00;      memory[20587] <=  8'h00;      memory[20588] <=  8'h00;      memory[20589] <=  8'h00;      memory[20590] <=  8'h00;      memory[20591] <=  8'h00;      memory[20592] <=  8'h00;      memory[20593] <=  8'h00;      memory[20594] <=  8'h00;      memory[20595] <=  8'h00;      memory[20596] <=  8'h00;      memory[20597] <=  8'h00;      memory[20598] <=  8'h00;      memory[20599] <=  8'h00;      memory[20600] <=  8'h00;      memory[20601] <=  8'h00;      memory[20602] <=  8'h00;      memory[20603] <=  8'h00;      memory[20604] <=  8'h00;      memory[20605] <=  8'h00;      memory[20606] <=  8'h00;      memory[20607] <=  8'h00;      memory[20608] <=  8'h00;      memory[20609] <=  8'h00;      memory[20610] <=  8'h00;      memory[20611] <=  8'h00;      memory[20612] <=  8'h00;      memory[20613] <=  8'h00;      memory[20614] <=  8'h00;      memory[20615] <=  8'h00;      memory[20616] <=  8'h00;      memory[20617] <=  8'h00;      memory[20618] <=  8'h00;      memory[20619] <=  8'h00;      memory[20620] <=  8'h00;      memory[20621] <=  8'h00;      memory[20622] <=  8'h00;      memory[20623] <=  8'h00;      memory[20624] <=  8'h00;      memory[20625] <=  8'h00;      memory[20626] <=  8'h00;      memory[20627] <=  8'h00;      memory[20628] <=  8'h00;      memory[20629] <=  8'h00;      memory[20630] <=  8'h00;      memory[20631] <=  8'h00;      memory[20632] <=  8'h00;      memory[20633] <=  8'h00;      memory[20634] <=  8'h00;      memory[20635] <=  8'h00;      memory[20636] <=  8'h00;      memory[20637] <=  8'h00;      memory[20638] <=  8'h00;      memory[20639] <=  8'h00;      memory[20640] <=  8'h00;      memory[20641] <=  8'h00;      memory[20642] <=  8'h00;      memory[20643] <=  8'h00;      memory[20644] <=  8'h00;      memory[20645] <=  8'h00;      memory[20646] <=  8'h00;      memory[20647] <=  8'h00;      memory[20648] <=  8'h00;      memory[20649] <=  8'h00;      memory[20650] <=  8'h00;      memory[20651] <=  8'h00;      memory[20652] <=  8'h00;      memory[20653] <=  8'h00;      memory[20654] <=  8'h00;      memory[20655] <=  8'h00;      memory[20656] <=  8'h00;      memory[20657] <=  8'h00;      memory[20658] <=  8'h00;      memory[20659] <=  8'h00;      memory[20660] <=  8'h00;      memory[20661] <=  8'h00;      memory[20662] <=  8'h00;      memory[20663] <=  8'h00;      memory[20664] <=  8'h00;      memory[20665] <=  8'h00;      memory[20666] <=  8'h00;      memory[20667] <=  8'h00;      memory[20668] <=  8'h00;      memory[20669] <=  8'h00;      memory[20670] <=  8'h00;      memory[20671] <=  8'h00;      memory[20672] <=  8'h00;      memory[20673] <=  8'h00;      memory[20674] <=  8'h00;      memory[20675] <=  8'h00;      memory[20676] <=  8'h00;      memory[20677] <=  8'h00;      memory[20678] <=  8'h00;      memory[20679] <=  8'h00;      memory[20680] <=  8'h00;      memory[20681] <=  8'h00;      memory[20682] <=  8'h00;      memory[20683] <=  8'h00;      memory[20684] <=  8'h00;      memory[20685] <=  8'h00;      memory[20686] <=  8'h00;      memory[20687] <=  8'h00;      memory[20688] <=  8'h00;      memory[20689] <=  8'h00;      memory[20690] <=  8'h00;      memory[20691] <=  8'h00;      memory[20692] <=  8'h00;      memory[20693] <=  8'h00;      memory[20694] <=  8'h00;      memory[20695] <=  8'h00;      memory[20696] <=  8'h00;      memory[20697] <=  8'h00;      memory[20698] <=  8'h00;      memory[20699] <=  8'h00;      memory[20700] <=  8'h00;      memory[20701] <=  8'h00;      memory[20702] <=  8'h00;      memory[20703] <=  8'h00;      memory[20704] <=  8'h00;      memory[20705] <=  8'h00;      memory[20706] <=  8'h00;      memory[20707] <=  8'h00;      memory[20708] <=  8'h00;      memory[20709] <=  8'h00;      memory[20710] <=  8'h00;      memory[20711] <=  8'h00;      memory[20712] <=  8'h00;      memory[20713] <=  8'h00;      memory[20714] <=  8'h00;      memory[20715] <=  8'h00;      memory[20716] <=  8'h00;      memory[20717] <=  8'h00;      memory[20718] <=  8'h00;      memory[20719] <=  8'h00;      memory[20720] <=  8'h00;      memory[20721] <=  8'h00;      memory[20722] <=  8'h00;      memory[20723] <=  8'h00;      memory[20724] <=  8'h00;      memory[20725] <=  8'h00;      memory[20726] <=  8'h00;      memory[20727] <=  8'h00;      memory[20728] <=  8'h00;      memory[20729] <=  8'h00;      memory[20730] <=  8'h00;      memory[20731] <=  8'h00;      memory[20732] <=  8'h00;      memory[20733] <=  8'h00;      memory[20734] <=  8'h00;      memory[20735] <=  8'h00;      memory[20736] <=  8'h00;      memory[20737] <=  8'h00;      memory[20738] <=  8'h00;      memory[20739] <=  8'h00;      memory[20740] <=  8'h00;      memory[20741] <=  8'h00;      memory[20742] <=  8'h00;      memory[20743] <=  8'h00;      memory[20744] <=  8'h00;      memory[20745] <=  8'h00;      memory[20746] <=  8'h00;      memory[20747] <=  8'h00;      memory[20748] <=  8'h00;      memory[20749] <=  8'h00;      memory[20750] <=  8'h00;      memory[20751] <=  8'h00;      memory[20752] <=  8'h00;      memory[20753] <=  8'h00;      memory[20754] <=  8'h00;      memory[20755] <=  8'h00;      memory[20756] <=  8'h00;      memory[20757] <=  8'h00;      memory[20758] <=  8'h00;      memory[20759] <=  8'h00;      memory[20760] <=  8'h00;      memory[20761] <=  8'h00;      memory[20762] <=  8'h00;      memory[20763] <=  8'h00;      memory[20764] <=  8'h00;      memory[20765] <=  8'h00;      memory[20766] <=  8'h00;      memory[20767] <=  8'h00;      memory[20768] <=  8'h00;      memory[20769] <=  8'h00;      memory[20770] <=  8'h00;      memory[20771] <=  8'h00;      memory[20772] <=  8'h00;      memory[20773] <=  8'h00;      memory[20774] <=  8'h00;      memory[20775] <=  8'h00;      memory[20776] <=  8'h00;      memory[20777] <=  8'h00;      memory[20778] <=  8'h00;      memory[20779] <=  8'h00;      memory[20780] <=  8'h00;      memory[20781] <=  8'h00;      memory[20782] <=  8'h00;      memory[20783] <=  8'h00;      memory[20784] <=  8'h00;      memory[20785] <=  8'h00;      memory[20786] <=  8'h00;      memory[20787] <=  8'h00;      memory[20788] <=  8'h00;      memory[20789] <=  8'h00;      memory[20790] <=  8'h00;      memory[20791] <=  8'h00;      memory[20792] <=  8'h00;      memory[20793] <=  8'h00;      memory[20794] <=  8'h00;      memory[20795] <=  8'h00;      memory[20796] <=  8'h00;      memory[20797] <=  8'h00;      memory[20798] <=  8'h00;      memory[20799] <=  8'h00;      memory[20800] <=  8'h00;      memory[20801] <=  8'h00;      memory[20802] <=  8'h00;      memory[20803] <=  8'h00;      memory[20804] <=  8'h00;      memory[20805] <=  8'h00;      memory[20806] <=  8'h00;      memory[20807] <=  8'h00;      memory[20808] <=  8'h00;      memory[20809] <=  8'h00;      memory[20810] <=  8'h00;      memory[20811] <=  8'h00;      memory[20812] <=  8'h00;      memory[20813] <=  8'h00;      memory[20814] <=  8'h00;      memory[20815] <=  8'h00;      memory[20816] <=  8'h00;      memory[20817] <=  8'h00;      memory[20818] <=  8'h00;      memory[20819] <=  8'h00;      memory[20820] <=  8'h00;      memory[20821] <=  8'h00;      memory[20822] <=  8'h00;      memory[20823] <=  8'h00;      memory[20824] <=  8'h00;      memory[20825] <=  8'h00;      memory[20826] <=  8'h00;      memory[20827] <=  8'h00;      memory[20828] <=  8'h00;      memory[20829] <=  8'h00;      memory[20830] <=  8'h00;      memory[20831] <=  8'h00;      memory[20832] <=  8'h00;      memory[20833] <=  8'h00;      memory[20834] <=  8'h00;      memory[20835] <=  8'h00;      memory[20836] <=  8'h00;      memory[20837] <=  8'h00;      memory[20838] <=  8'h00;      memory[20839] <=  8'h00;      memory[20840] <=  8'h00;      memory[20841] <=  8'h00;      memory[20842] <=  8'h00;      memory[20843] <=  8'h00;      memory[20844] <=  8'h00;      memory[20845] <=  8'h00;      memory[20846] <=  8'h00;      memory[20847] <=  8'h00;      memory[20848] <=  8'h00;      memory[20849] <=  8'h00;      memory[20850] <=  8'h00;      memory[20851] <=  8'h00;      memory[20852] <=  8'h00;      memory[20853] <=  8'h00;      memory[20854] <=  8'h00;      memory[20855] <=  8'h00;      memory[20856] <=  8'h00;      memory[20857] <=  8'h00;      memory[20858] <=  8'h00;      memory[20859] <=  8'h00;      memory[20860] <=  8'h00;      memory[20861] <=  8'h00;      memory[20862] <=  8'h00;      memory[20863] <=  8'h00;      memory[20864] <=  8'h00;      memory[20865] <=  8'h00;      memory[20866] <=  8'h00;      memory[20867] <=  8'h00;      memory[20868] <=  8'h00;      memory[20869] <=  8'h00;      memory[20870] <=  8'h00;      memory[20871] <=  8'h00;      memory[20872] <=  8'h00;      memory[20873] <=  8'h00;      memory[20874] <=  8'h00;      memory[20875] <=  8'h00;      memory[20876] <=  8'h00;      memory[20877] <=  8'h00;      memory[20878] <=  8'h00;      memory[20879] <=  8'h00;      memory[20880] <=  8'h00;      memory[20881] <=  8'h00;      memory[20882] <=  8'h00;      memory[20883] <=  8'h00;      memory[20884] <=  8'h00;      memory[20885] <=  8'h00;      memory[20886] <=  8'h00;      memory[20887] <=  8'h00;      memory[20888] <=  8'h00;      memory[20889] <=  8'h00;      memory[20890] <=  8'h00;      memory[20891] <=  8'h00;      memory[20892] <=  8'h00;      memory[20893] <=  8'h00;      memory[20894] <=  8'h00;      memory[20895] <=  8'h00;      memory[20896] <=  8'h00;      memory[20897] <=  8'h00;      memory[20898] <=  8'h00;      memory[20899] <=  8'h00;      memory[20900] <=  8'h00;      memory[20901] <=  8'h00;      memory[20902] <=  8'h00;      memory[20903] <=  8'h00;      memory[20904] <=  8'h00;      memory[20905] <=  8'h00;      memory[20906] <=  8'h00;      memory[20907] <=  8'h00;      memory[20908] <=  8'h00;      memory[20909] <=  8'h00;      memory[20910] <=  8'h00;      memory[20911] <=  8'h00;      memory[20912] <=  8'h00;      memory[20913] <=  8'h00;      memory[20914] <=  8'h00;      memory[20915] <=  8'h00;      memory[20916] <=  8'h00;      memory[20917] <=  8'h00;      memory[20918] <=  8'h00;      memory[20919] <=  8'h00;      memory[20920] <=  8'h00;      memory[20921] <=  8'h00;      memory[20922] <=  8'h00;      memory[20923] <=  8'h00;      memory[20924] <=  8'h00;      memory[20925] <=  8'h00;      memory[20926] <=  8'h00;      memory[20927] <=  8'h00;      memory[20928] <=  8'h00;      memory[20929] <=  8'h00;      memory[20930] <=  8'h00;      memory[20931] <=  8'h00;      memory[20932] <=  8'h00;      memory[20933] <=  8'h00;      memory[20934] <=  8'h00;      memory[20935] <=  8'h00;      memory[20936] <=  8'h00;      memory[20937] <=  8'h00;      memory[20938] <=  8'h00;      memory[20939] <=  8'h00;      memory[20940] <=  8'h00;      memory[20941] <=  8'h00;      memory[20942] <=  8'h00;      memory[20943] <=  8'h00;      memory[20944] <=  8'h00;      memory[20945] <=  8'h00;      memory[20946] <=  8'h00;      memory[20947] <=  8'h00;      memory[20948] <=  8'h00;      memory[20949] <=  8'h00;      memory[20950] <=  8'h00;      memory[20951] <=  8'h00;      memory[20952] <=  8'h00;      memory[20953] <=  8'h00;      memory[20954] <=  8'h00;      memory[20955] <=  8'h00;      memory[20956] <=  8'h00;      memory[20957] <=  8'h00;      memory[20958] <=  8'h00;      memory[20959] <=  8'h00;      memory[20960] <=  8'h00;      memory[20961] <=  8'h00;      memory[20962] <=  8'h00;      memory[20963] <=  8'h00;      memory[20964] <=  8'h00;      memory[20965] <=  8'h00;      memory[20966] <=  8'h00;      memory[20967] <=  8'h00;      memory[20968] <=  8'h00;      memory[20969] <=  8'h00;      memory[20970] <=  8'h00;      memory[20971] <=  8'h00;      memory[20972] <=  8'h00;      memory[20973] <=  8'h00;      memory[20974] <=  8'h00;      memory[20975] <=  8'h00;      memory[20976] <=  8'h00;      memory[20977] <=  8'h00;      memory[20978] <=  8'h00;      memory[20979] <=  8'h00;      memory[20980] <=  8'h00;      memory[20981] <=  8'h00;      memory[20982] <=  8'h00;      memory[20983] <=  8'h00;      memory[20984] <=  8'h00;      memory[20985] <=  8'h00;      memory[20986] <=  8'h00;      memory[20987] <=  8'h00;      memory[20988] <=  8'h00;      memory[20989] <=  8'h00;      memory[20990] <=  8'h00;      memory[20991] <=  8'h00;      memory[20992] <=  8'h00;      memory[20993] <=  8'h00;      memory[20994] <=  8'h00;      memory[20995] <=  8'h00;      memory[20996] <=  8'h00;      memory[20997] <=  8'h00;      memory[20998] <=  8'h00;      memory[20999] <=  8'h00;      memory[21000] <=  8'h00;      memory[21001] <=  8'h00;      memory[21002] <=  8'h00;      memory[21003] <=  8'h00;      memory[21004] <=  8'h00;      memory[21005] <=  8'h00;      memory[21006] <=  8'h00;      memory[21007] <=  8'h00;      memory[21008] <=  8'h00;      memory[21009] <=  8'h00;      memory[21010] <=  8'h00;      memory[21011] <=  8'h00;      memory[21012] <=  8'h00;      memory[21013] <=  8'h00;      memory[21014] <=  8'h00;      memory[21015] <=  8'h00;      memory[21016] <=  8'h00;      memory[21017] <=  8'h00;      memory[21018] <=  8'h00;      memory[21019] <=  8'h00;      memory[21020] <=  8'h00;      memory[21021] <=  8'h00;      memory[21022] <=  8'h00;      memory[21023] <=  8'h00;      memory[21024] <=  8'h00;      memory[21025] <=  8'h00;      memory[21026] <=  8'h00;      memory[21027] <=  8'h00;      memory[21028] <=  8'h00;      memory[21029] <=  8'h00;      memory[21030] <=  8'h00;      memory[21031] <=  8'h00;      memory[21032] <=  8'h00;      memory[21033] <=  8'h00;      memory[21034] <=  8'h00;      memory[21035] <=  8'h00;      memory[21036] <=  8'h00;      memory[21037] <=  8'h00;      memory[21038] <=  8'h00;      memory[21039] <=  8'h00;      memory[21040] <=  8'h00;      memory[21041] <=  8'h00;      memory[21042] <=  8'h00;      memory[21043] <=  8'h00;      memory[21044] <=  8'h00;      memory[21045] <=  8'h00;      memory[21046] <=  8'h00;      memory[21047] <=  8'h00;      memory[21048] <=  8'h00;      memory[21049] <=  8'h00;      memory[21050] <=  8'h00;      memory[21051] <=  8'h00;      memory[21052] <=  8'h00;      memory[21053] <=  8'h00;      memory[21054] <=  8'h00;      memory[21055] <=  8'h00;      memory[21056] <=  8'h00;      memory[21057] <=  8'h00;      memory[21058] <=  8'h00;      memory[21059] <=  8'h00;      memory[21060] <=  8'h00;      memory[21061] <=  8'h00;      memory[21062] <=  8'h00;      memory[21063] <=  8'h00;      memory[21064] <=  8'h00;      memory[21065] <=  8'h00;      memory[21066] <=  8'h00;      memory[21067] <=  8'h00;      memory[21068] <=  8'h00;      memory[21069] <=  8'h00;      memory[21070] <=  8'h00;      memory[21071] <=  8'h00;      memory[21072] <=  8'h00;      memory[21073] <=  8'h00;      memory[21074] <=  8'h00;      memory[21075] <=  8'h00;      memory[21076] <=  8'h00;      memory[21077] <=  8'h00;      memory[21078] <=  8'h00;      memory[21079] <=  8'h00;      memory[21080] <=  8'h00;      memory[21081] <=  8'h00;      memory[21082] <=  8'h00;      memory[21083] <=  8'h00;      memory[21084] <=  8'h00;      memory[21085] <=  8'h00;      memory[21086] <=  8'h00;      memory[21087] <=  8'h00;      memory[21088] <=  8'h00;      memory[21089] <=  8'h00;      memory[21090] <=  8'h00;      memory[21091] <=  8'h00;      memory[21092] <=  8'h00;      memory[21093] <=  8'h00;      memory[21094] <=  8'h00;      memory[21095] <=  8'h00;      memory[21096] <=  8'h00;      memory[21097] <=  8'h00;      memory[21098] <=  8'h00;      memory[21099] <=  8'h00;      memory[21100] <=  8'h00;      memory[21101] <=  8'h00;      memory[21102] <=  8'h00;      memory[21103] <=  8'h00;      memory[21104] <=  8'h00;      memory[21105] <=  8'h00;      memory[21106] <=  8'h00;      memory[21107] <=  8'h00;      memory[21108] <=  8'h00;      memory[21109] <=  8'h00;      memory[21110] <=  8'h00;      memory[21111] <=  8'h00;      memory[21112] <=  8'h00;      memory[21113] <=  8'h00;      memory[21114] <=  8'h00;      memory[21115] <=  8'h00;      memory[21116] <=  8'h00;      memory[21117] <=  8'h00;      memory[21118] <=  8'h00;      memory[21119] <=  8'h00;      memory[21120] <=  8'h00;      memory[21121] <=  8'h00;      memory[21122] <=  8'h00;      memory[21123] <=  8'h00;      memory[21124] <=  8'h00;      memory[21125] <=  8'h00;      memory[21126] <=  8'h00;      memory[21127] <=  8'h00;      memory[21128] <=  8'h00;      memory[21129] <=  8'h00;      memory[21130] <=  8'h00;      memory[21131] <=  8'h00;      memory[21132] <=  8'h00;      memory[21133] <=  8'h00;      memory[21134] <=  8'h00;      memory[21135] <=  8'h00;      memory[21136] <=  8'h00;      memory[21137] <=  8'h00;      memory[21138] <=  8'h00;      memory[21139] <=  8'h00;      memory[21140] <=  8'h00;      memory[21141] <=  8'h00;      memory[21142] <=  8'h00;      memory[21143] <=  8'h00;      memory[21144] <=  8'h00;      memory[21145] <=  8'h00;      memory[21146] <=  8'h00;      memory[21147] <=  8'h00;      memory[21148] <=  8'h00;      memory[21149] <=  8'h00;      memory[21150] <=  8'h00;      memory[21151] <=  8'h00;      memory[21152] <=  8'h00;      memory[21153] <=  8'h00;      memory[21154] <=  8'h00;      memory[21155] <=  8'h00;      memory[21156] <=  8'h00;      memory[21157] <=  8'h00;      memory[21158] <=  8'h00;      memory[21159] <=  8'h00;      memory[21160] <=  8'h00;      memory[21161] <=  8'h00;      memory[21162] <=  8'h00;      memory[21163] <=  8'h00;      memory[21164] <=  8'h00;      memory[21165] <=  8'h00;      memory[21166] <=  8'h00;      memory[21167] <=  8'h00;      memory[21168] <=  8'h00;      memory[21169] <=  8'h00;      memory[21170] <=  8'h00;      memory[21171] <=  8'h00;      memory[21172] <=  8'h00;      memory[21173] <=  8'h00;      memory[21174] <=  8'h00;      memory[21175] <=  8'h00;      memory[21176] <=  8'h00;      memory[21177] <=  8'h00;      memory[21178] <=  8'h00;      memory[21179] <=  8'h00;      memory[21180] <=  8'h00;      memory[21181] <=  8'h00;      memory[21182] <=  8'h00;      memory[21183] <=  8'h00;      memory[21184] <=  8'h00;      memory[21185] <=  8'h00;      memory[21186] <=  8'h00;      memory[21187] <=  8'h00;      memory[21188] <=  8'h00;      memory[21189] <=  8'h00;      memory[21190] <=  8'h00;      memory[21191] <=  8'h00;      memory[21192] <=  8'h00;      memory[21193] <=  8'h00;      memory[21194] <=  8'h00;      memory[21195] <=  8'h00;      memory[21196] <=  8'h00;      memory[21197] <=  8'h00;      memory[21198] <=  8'h00;      memory[21199] <=  8'h00;      memory[21200] <=  8'h00;      memory[21201] <=  8'h00;      memory[21202] <=  8'h00;      memory[21203] <=  8'h00;      memory[21204] <=  8'h00;      memory[21205] <=  8'h00;      memory[21206] <=  8'h00;      memory[21207] <=  8'h00;      memory[21208] <=  8'h00;      memory[21209] <=  8'h00;      memory[21210] <=  8'h00;      memory[21211] <=  8'h00;      memory[21212] <=  8'h00;      memory[21213] <=  8'h00;      memory[21214] <=  8'h00;      memory[21215] <=  8'h00;      memory[21216] <=  8'h00;      memory[21217] <=  8'h00;      memory[21218] <=  8'h00;      memory[21219] <=  8'h00;      memory[21220] <=  8'h00;      memory[21221] <=  8'h00;      memory[21222] <=  8'h00;      memory[21223] <=  8'h00;      memory[21224] <=  8'h00;      memory[21225] <=  8'h00;      memory[21226] <=  8'h00;      memory[21227] <=  8'h00;      memory[21228] <=  8'h00;      memory[21229] <=  8'h00;      memory[21230] <=  8'h00;      memory[21231] <=  8'h00;      memory[21232] <=  8'h00;      memory[21233] <=  8'h00;      memory[21234] <=  8'h00;      memory[21235] <=  8'h00;      memory[21236] <=  8'h00;      memory[21237] <=  8'h00;      memory[21238] <=  8'h00;      memory[21239] <=  8'h00;      memory[21240] <=  8'h00;      memory[21241] <=  8'h00;      memory[21242] <=  8'h00;      memory[21243] <=  8'h00;      memory[21244] <=  8'h00;      memory[21245] <=  8'h00;      memory[21246] <=  8'h00;      memory[21247] <=  8'h00;      memory[21248] <=  8'h00;      memory[21249] <=  8'h00;      memory[21250] <=  8'h00;      memory[21251] <=  8'h00;      memory[21252] <=  8'h00;      memory[21253] <=  8'h00;      memory[21254] <=  8'h00;      memory[21255] <=  8'h00;      memory[21256] <=  8'h00;      memory[21257] <=  8'h00;      memory[21258] <=  8'h00;      memory[21259] <=  8'h00;      memory[21260] <=  8'h00;      memory[21261] <=  8'h00;      memory[21262] <=  8'h00;      memory[21263] <=  8'h00;      memory[21264] <=  8'h00;      memory[21265] <=  8'h00;      memory[21266] <=  8'h00;      memory[21267] <=  8'h00;      memory[21268] <=  8'h00;      memory[21269] <=  8'h00;      memory[21270] <=  8'h00;      memory[21271] <=  8'h00;      memory[21272] <=  8'h00;      memory[21273] <=  8'h00;      memory[21274] <=  8'h00;      memory[21275] <=  8'h00;      memory[21276] <=  8'h00;      memory[21277] <=  8'h00;      memory[21278] <=  8'h00;      memory[21279] <=  8'h00;      memory[21280] <=  8'h00;      memory[21281] <=  8'h00;      memory[21282] <=  8'h00;      memory[21283] <=  8'h00;      memory[21284] <=  8'h00;      memory[21285] <=  8'h00;      memory[21286] <=  8'h00;      memory[21287] <=  8'h00;      memory[21288] <=  8'h00;      memory[21289] <=  8'h00;      memory[21290] <=  8'h00;      memory[21291] <=  8'h00;      memory[21292] <=  8'h00;      memory[21293] <=  8'h00;      memory[21294] <=  8'h00;      memory[21295] <=  8'h00;      memory[21296] <=  8'h00;      memory[21297] <=  8'h00;      memory[21298] <=  8'h00;      memory[21299] <=  8'h00;      memory[21300] <=  8'h00;      memory[21301] <=  8'h00;      memory[21302] <=  8'h00;      memory[21303] <=  8'h00;      memory[21304] <=  8'h00;      memory[21305] <=  8'h00;      memory[21306] <=  8'h00;      memory[21307] <=  8'h00;      memory[21308] <=  8'h00;      memory[21309] <=  8'h00;      memory[21310] <=  8'h00;      memory[21311] <=  8'h00;      memory[21312] <=  8'h00;      memory[21313] <=  8'h00;      memory[21314] <=  8'h00;      memory[21315] <=  8'h00;      memory[21316] <=  8'h00;      memory[21317] <=  8'h00;      memory[21318] <=  8'h00;      memory[21319] <=  8'h00;      memory[21320] <=  8'h00;      memory[21321] <=  8'h00;      memory[21322] <=  8'h00;      memory[21323] <=  8'h00;      memory[21324] <=  8'h00;      memory[21325] <=  8'h00;      memory[21326] <=  8'h00;      memory[21327] <=  8'h00;      memory[21328] <=  8'h00;      memory[21329] <=  8'h00;      memory[21330] <=  8'h00;      memory[21331] <=  8'h00;      memory[21332] <=  8'h00;      memory[21333] <=  8'h00;      memory[21334] <=  8'h00;      memory[21335] <=  8'h00;      memory[21336] <=  8'h00;      memory[21337] <=  8'h00;      memory[21338] <=  8'h00;      memory[21339] <=  8'h00;      memory[21340] <=  8'h00;      memory[21341] <=  8'h00;      memory[21342] <=  8'h00;      memory[21343] <=  8'h00;      memory[21344] <=  8'h00;      memory[21345] <=  8'h00;      memory[21346] <=  8'h00;      memory[21347] <=  8'h00;      memory[21348] <=  8'h00;      memory[21349] <=  8'h00;      memory[21350] <=  8'h00;      memory[21351] <=  8'h00;      memory[21352] <=  8'h00;      memory[21353] <=  8'h00;      memory[21354] <=  8'h00;      memory[21355] <=  8'h00;      memory[21356] <=  8'h00;      memory[21357] <=  8'h00;      memory[21358] <=  8'h00;      memory[21359] <=  8'h00;      memory[21360] <=  8'h00;      memory[21361] <=  8'h00;      memory[21362] <=  8'h00;      memory[21363] <=  8'h00;      memory[21364] <=  8'h00;      memory[21365] <=  8'h00;      memory[21366] <=  8'h00;      memory[21367] <=  8'h00;      memory[21368] <=  8'h00;      memory[21369] <=  8'h00;      memory[21370] <=  8'h00;      memory[21371] <=  8'h00;      memory[21372] <=  8'h00;      memory[21373] <=  8'h00;      memory[21374] <=  8'h00;      memory[21375] <=  8'h00;      memory[21376] <=  8'h00;      memory[21377] <=  8'h00;      memory[21378] <=  8'h00;      memory[21379] <=  8'h00;      memory[21380] <=  8'h00;      memory[21381] <=  8'h00;      memory[21382] <=  8'h00;      memory[21383] <=  8'h00;      memory[21384] <=  8'h00;      memory[21385] <=  8'h00;      memory[21386] <=  8'h00;      memory[21387] <=  8'h00;      memory[21388] <=  8'h00;      memory[21389] <=  8'h00;      memory[21390] <=  8'h00;      memory[21391] <=  8'h00;      memory[21392] <=  8'h00;      memory[21393] <=  8'h00;      memory[21394] <=  8'h00;      memory[21395] <=  8'h00;      memory[21396] <=  8'h00;      memory[21397] <=  8'h00;      memory[21398] <=  8'h00;      memory[21399] <=  8'h00;      memory[21400] <=  8'h00;      memory[21401] <=  8'h00;      memory[21402] <=  8'h00;      memory[21403] <=  8'h00;      memory[21404] <=  8'h00;      memory[21405] <=  8'h00;      memory[21406] <=  8'h00;      memory[21407] <=  8'h00;      memory[21408] <=  8'h00;      memory[21409] <=  8'h00;      memory[21410] <=  8'h00;      memory[21411] <=  8'h00;      memory[21412] <=  8'h00;      memory[21413] <=  8'h00;      memory[21414] <=  8'h00;      memory[21415] <=  8'h00;      memory[21416] <=  8'h00;      memory[21417] <=  8'h00;      memory[21418] <=  8'h00;      memory[21419] <=  8'h00;      memory[21420] <=  8'h00;      memory[21421] <=  8'h00;      memory[21422] <=  8'h00;      memory[21423] <=  8'h00;      memory[21424] <=  8'h00;      memory[21425] <=  8'h00;      memory[21426] <=  8'h00;      memory[21427] <=  8'h00;      memory[21428] <=  8'h00;      memory[21429] <=  8'h00;      memory[21430] <=  8'h00;      memory[21431] <=  8'h00;      memory[21432] <=  8'h00;      memory[21433] <=  8'h00;      memory[21434] <=  8'h00;      memory[21435] <=  8'h00;      memory[21436] <=  8'h00;      memory[21437] <=  8'h00;      memory[21438] <=  8'h00;      memory[21439] <=  8'h00;      memory[21440] <=  8'h00;      memory[21441] <=  8'h00;      memory[21442] <=  8'h00;      memory[21443] <=  8'h00;      memory[21444] <=  8'h00;      memory[21445] <=  8'h00;      memory[21446] <=  8'h00;      memory[21447] <=  8'h00;      memory[21448] <=  8'h00;      memory[21449] <=  8'h00;      memory[21450] <=  8'h00;      memory[21451] <=  8'h00;      memory[21452] <=  8'h00;      memory[21453] <=  8'h00;      memory[21454] <=  8'h00;      memory[21455] <=  8'h00;      memory[21456] <=  8'h00;      memory[21457] <=  8'h00;      memory[21458] <=  8'h00;      memory[21459] <=  8'h00;      memory[21460] <=  8'h00;      memory[21461] <=  8'h00;      memory[21462] <=  8'h00;      memory[21463] <=  8'h00;      memory[21464] <=  8'h00;      memory[21465] <=  8'h00;      memory[21466] <=  8'h00;      memory[21467] <=  8'h00;      memory[21468] <=  8'h00;      memory[21469] <=  8'h00;      memory[21470] <=  8'h00;      memory[21471] <=  8'h00;      memory[21472] <=  8'h00;      memory[21473] <=  8'h00;      memory[21474] <=  8'h00;      memory[21475] <=  8'h00;      memory[21476] <=  8'h00;      memory[21477] <=  8'h00;      memory[21478] <=  8'h00;      memory[21479] <=  8'h00;      memory[21480] <=  8'h00;      memory[21481] <=  8'h00;      memory[21482] <=  8'h00;      memory[21483] <=  8'h00;      memory[21484] <=  8'h00;      memory[21485] <=  8'h00;      memory[21486] <=  8'h00;      memory[21487] <=  8'h00;      memory[21488] <=  8'h00;      memory[21489] <=  8'h00;      memory[21490] <=  8'h00;      memory[21491] <=  8'h00;      memory[21492] <=  8'h00;      memory[21493] <=  8'h00;      memory[21494] <=  8'h00;      memory[21495] <=  8'h00;      memory[21496] <=  8'h00;      memory[21497] <=  8'h00;      memory[21498] <=  8'h00;      memory[21499] <=  8'h00;      memory[21500] <=  8'h00;      memory[21501] <=  8'h00;      memory[21502] <=  8'h00;      memory[21503] <=  8'h00;      memory[21504] <=  8'h00;      memory[21505] <=  8'h00;      memory[21506] <=  8'h00;      memory[21507] <=  8'h00;      memory[21508] <=  8'h00;      memory[21509] <=  8'h00;      memory[21510] <=  8'h00;      memory[21511] <=  8'h00;      memory[21512] <=  8'h00;      memory[21513] <=  8'h00;      memory[21514] <=  8'h00;      memory[21515] <=  8'h00;      memory[21516] <=  8'h00;      memory[21517] <=  8'h00;      memory[21518] <=  8'h00;      memory[21519] <=  8'h00;      memory[21520] <=  8'h00;      memory[21521] <=  8'h00;      memory[21522] <=  8'h00;      memory[21523] <=  8'h00;      memory[21524] <=  8'h00;      memory[21525] <=  8'h00;      memory[21526] <=  8'h00;      memory[21527] <=  8'h00;      memory[21528] <=  8'h00;      memory[21529] <=  8'h00;      memory[21530] <=  8'h00;      memory[21531] <=  8'h00;      memory[21532] <=  8'h00;      memory[21533] <=  8'h00;      memory[21534] <=  8'h00;      memory[21535] <=  8'h00;      memory[21536] <=  8'h00;      memory[21537] <=  8'h00;      memory[21538] <=  8'h00;      memory[21539] <=  8'h00;      memory[21540] <=  8'h00;      memory[21541] <=  8'h00;      memory[21542] <=  8'h00;      memory[21543] <=  8'h00;      memory[21544] <=  8'h00;      memory[21545] <=  8'h00;      memory[21546] <=  8'h00;      memory[21547] <=  8'h00;      memory[21548] <=  8'h00;      memory[21549] <=  8'h00;      memory[21550] <=  8'h00;      memory[21551] <=  8'h00;      memory[21552] <=  8'h00;      memory[21553] <=  8'h00;      memory[21554] <=  8'h00;      memory[21555] <=  8'h00;      memory[21556] <=  8'h00;      memory[21557] <=  8'h00;      memory[21558] <=  8'h00;      memory[21559] <=  8'h00;      memory[21560] <=  8'h00;      memory[21561] <=  8'h00;      memory[21562] <=  8'h00;      memory[21563] <=  8'h00;      memory[21564] <=  8'h00;      memory[21565] <=  8'h00;      memory[21566] <=  8'h00;      memory[21567] <=  8'h00;      memory[21568] <=  8'h00;      memory[21569] <=  8'h00;      memory[21570] <=  8'h00;      memory[21571] <=  8'h00;      memory[21572] <=  8'h00;      memory[21573] <=  8'h00;      memory[21574] <=  8'h00;      memory[21575] <=  8'h00;      memory[21576] <=  8'h00;      memory[21577] <=  8'h00;      memory[21578] <=  8'h00;      memory[21579] <=  8'h00;      memory[21580] <=  8'h00;      memory[21581] <=  8'h00;      memory[21582] <=  8'h00;      memory[21583] <=  8'h00;      memory[21584] <=  8'h00;      memory[21585] <=  8'h00;      memory[21586] <=  8'h00;      memory[21587] <=  8'h00;      memory[21588] <=  8'h00;      memory[21589] <=  8'h00;      memory[21590] <=  8'h00;      memory[21591] <=  8'h00;      memory[21592] <=  8'h00;      memory[21593] <=  8'h00;      memory[21594] <=  8'h00;      memory[21595] <=  8'h00;      memory[21596] <=  8'h00;      memory[21597] <=  8'h00;      memory[21598] <=  8'h00;      memory[21599] <=  8'h00;      memory[21600] <=  8'h00;      memory[21601] <=  8'h00;      memory[21602] <=  8'h00;      memory[21603] <=  8'h00;      memory[21604] <=  8'h00;      memory[21605] <=  8'h00;      memory[21606] <=  8'h00;      memory[21607] <=  8'h00;      memory[21608] <=  8'h00;      memory[21609] <=  8'h00;      memory[21610] <=  8'h00;      memory[21611] <=  8'h00;      memory[21612] <=  8'h00;      memory[21613] <=  8'h00;      memory[21614] <=  8'h00;      memory[21615] <=  8'h00;      memory[21616] <=  8'h00;      memory[21617] <=  8'h00;      memory[21618] <=  8'h00;      memory[21619] <=  8'h00;      memory[21620] <=  8'h00;      memory[21621] <=  8'h00;      memory[21622] <=  8'h00;      memory[21623] <=  8'h00;      memory[21624] <=  8'h00;      memory[21625] <=  8'h00;      memory[21626] <=  8'h00;      memory[21627] <=  8'h00;      memory[21628] <=  8'h00;      memory[21629] <=  8'h00;      memory[21630] <=  8'h00;      memory[21631] <=  8'h00;      memory[21632] <=  8'h00;      memory[21633] <=  8'h00;      memory[21634] <=  8'h00;      memory[21635] <=  8'h00;      memory[21636] <=  8'h00;      memory[21637] <=  8'h00;      memory[21638] <=  8'h00;      memory[21639] <=  8'h00;      memory[21640] <=  8'h00;      memory[21641] <=  8'h00;      memory[21642] <=  8'h00;      memory[21643] <=  8'h00;      memory[21644] <=  8'h00;      memory[21645] <=  8'h00;      memory[21646] <=  8'h00;      memory[21647] <=  8'h00;      memory[21648] <=  8'h00;      memory[21649] <=  8'h00;      memory[21650] <=  8'h00;      memory[21651] <=  8'h00;      memory[21652] <=  8'h00;      memory[21653] <=  8'h00;      memory[21654] <=  8'h00;      memory[21655] <=  8'h00;      memory[21656] <=  8'h00;      memory[21657] <=  8'h00;      memory[21658] <=  8'h00;      memory[21659] <=  8'h00;      memory[21660] <=  8'h00;      memory[21661] <=  8'h00;      memory[21662] <=  8'h00;      memory[21663] <=  8'h00;      memory[21664] <=  8'h00;      memory[21665] <=  8'h00;      memory[21666] <=  8'h00;      memory[21667] <=  8'h00;      memory[21668] <=  8'h00;      memory[21669] <=  8'h00;      memory[21670] <=  8'h00;      memory[21671] <=  8'h00;      memory[21672] <=  8'h00;      memory[21673] <=  8'h00;      memory[21674] <=  8'h00;      memory[21675] <=  8'h00;      memory[21676] <=  8'h00;      memory[21677] <=  8'h00;      memory[21678] <=  8'h00;      memory[21679] <=  8'h00;      memory[21680] <=  8'h00;      memory[21681] <=  8'h00;      memory[21682] <=  8'h00;      memory[21683] <=  8'h00;      memory[21684] <=  8'h00;      memory[21685] <=  8'h00;      memory[21686] <=  8'h00;      memory[21687] <=  8'h00;      memory[21688] <=  8'h00;      memory[21689] <=  8'h00;      memory[21690] <=  8'h00;      memory[21691] <=  8'h00;      memory[21692] <=  8'h00;      memory[21693] <=  8'h00;      memory[21694] <=  8'h00;      memory[21695] <=  8'h00;      memory[21696] <=  8'h00;      memory[21697] <=  8'h00;      memory[21698] <=  8'h00;      memory[21699] <=  8'h00;      memory[21700] <=  8'h00;      memory[21701] <=  8'h00;      memory[21702] <=  8'h00;      memory[21703] <=  8'h00;      memory[21704] <=  8'h00;      memory[21705] <=  8'h00;      memory[21706] <=  8'h00;      memory[21707] <=  8'h00;      memory[21708] <=  8'h00;      memory[21709] <=  8'h00;      memory[21710] <=  8'h00;      memory[21711] <=  8'h00;      memory[21712] <=  8'h00;      memory[21713] <=  8'h00;      memory[21714] <=  8'h00;      memory[21715] <=  8'h00;      memory[21716] <=  8'h00;      memory[21717] <=  8'h00;      memory[21718] <=  8'h00;      memory[21719] <=  8'h00;      memory[21720] <=  8'h00;      memory[21721] <=  8'h00;      memory[21722] <=  8'h00;      memory[21723] <=  8'h00;      memory[21724] <=  8'h00;      memory[21725] <=  8'h00;      memory[21726] <=  8'h00;      memory[21727] <=  8'h00;      memory[21728] <=  8'h00;      memory[21729] <=  8'h00;      memory[21730] <=  8'h00;      memory[21731] <=  8'h00;      memory[21732] <=  8'h00;      memory[21733] <=  8'h00;      memory[21734] <=  8'h00;      memory[21735] <=  8'h00;      memory[21736] <=  8'h00;      memory[21737] <=  8'h00;      memory[21738] <=  8'h00;      memory[21739] <=  8'h00;      memory[21740] <=  8'h00;      memory[21741] <=  8'h00;      memory[21742] <=  8'h00;      memory[21743] <=  8'h00;      memory[21744] <=  8'h00;      memory[21745] <=  8'h00;      memory[21746] <=  8'h00;      memory[21747] <=  8'h00;      memory[21748] <=  8'h00;      memory[21749] <=  8'h00;      memory[21750] <=  8'h00;      memory[21751] <=  8'h00;      memory[21752] <=  8'h00;      memory[21753] <=  8'h00;      memory[21754] <=  8'h00;      memory[21755] <=  8'h00;      memory[21756] <=  8'h00;      memory[21757] <=  8'h00;      memory[21758] <=  8'h00;      memory[21759] <=  8'h00;      memory[21760] <=  8'h00;      memory[21761] <=  8'h00;      memory[21762] <=  8'h00;      memory[21763] <=  8'h00;      memory[21764] <=  8'h00;      memory[21765] <=  8'h00;      memory[21766] <=  8'h00;      memory[21767] <=  8'h00;      memory[21768] <=  8'h00;      memory[21769] <=  8'h00;      memory[21770] <=  8'h00;      memory[21771] <=  8'h00;      memory[21772] <=  8'h00;      memory[21773] <=  8'h00;      memory[21774] <=  8'h00;      memory[21775] <=  8'h00;      memory[21776] <=  8'h00;      memory[21777] <=  8'h00;      memory[21778] <=  8'h00;      memory[21779] <=  8'h00;      memory[21780] <=  8'h00;      memory[21781] <=  8'h00;      memory[21782] <=  8'h00;      memory[21783] <=  8'h00;      memory[21784] <=  8'h00;      memory[21785] <=  8'h00;      memory[21786] <=  8'h00;      memory[21787] <=  8'h00;      memory[21788] <=  8'h00;      memory[21789] <=  8'h00;      memory[21790] <=  8'h00;      memory[21791] <=  8'h00;      memory[21792] <=  8'h00;      memory[21793] <=  8'h00;      memory[21794] <=  8'h00;      memory[21795] <=  8'h00;      memory[21796] <=  8'h00;      memory[21797] <=  8'h00;      memory[21798] <=  8'h00;      memory[21799] <=  8'h00;      memory[21800] <=  8'h00;      memory[21801] <=  8'h00;      memory[21802] <=  8'h00;      memory[21803] <=  8'h00;      memory[21804] <=  8'h00;      memory[21805] <=  8'h00;      memory[21806] <=  8'h00;      memory[21807] <=  8'h00;      memory[21808] <=  8'h00;      memory[21809] <=  8'h00;      memory[21810] <=  8'h00;      memory[21811] <=  8'h00;      memory[21812] <=  8'h00;      memory[21813] <=  8'h00;      memory[21814] <=  8'h00;      memory[21815] <=  8'h00;      memory[21816] <=  8'h00;      memory[21817] <=  8'h00;      memory[21818] <=  8'h00;      memory[21819] <=  8'h00;      memory[21820] <=  8'h00;      memory[21821] <=  8'h00;      memory[21822] <=  8'h00;      memory[21823] <=  8'h00;      memory[21824] <=  8'h00;      memory[21825] <=  8'h00;      memory[21826] <=  8'h00;      memory[21827] <=  8'h00;      memory[21828] <=  8'h00;      memory[21829] <=  8'h00;      memory[21830] <=  8'h00;      memory[21831] <=  8'h00;      memory[21832] <=  8'h00;      memory[21833] <=  8'h00;      memory[21834] <=  8'h00;      memory[21835] <=  8'h00;      memory[21836] <=  8'h00;      memory[21837] <=  8'h00;      memory[21838] <=  8'h00;      memory[21839] <=  8'h00;      memory[21840] <=  8'h00;      memory[21841] <=  8'h00;      memory[21842] <=  8'h00;      memory[21843] <=  8'h00;      memory[21844] <=  8'h00;      memory[21845] <=  8'h00;      memory[21846] <=  8'h00;      memory[21847] <=  8'h00;      memory[21848] <=  8'h00;      memory[21849] <=  8'h00;      memory[21850] <=  8'h00;      memory[21851] <=  8'h00;      memory[21852] <=  8'h00;      memory[21853] <=  8'h00;      memory[21854] <=  8'h00;      memory[21855] <=  8'h00;      memory[21856] <=  8'h00;      memory[21857] <=  8'h00;      memory[21858] <=  8'h00;      memory[21859] <=  8'h00;      memory[21860] <=  8'h00;      memory[21861] <=  8'h00;      memory[21862] <=  8'h00;      memory[21863] <=  8'h00;      memory[21864] <=  8'h00;      memory[21865] <=  8'h00;      memory[21866] <=  8'h00;      memory[21867] <=  8'h00;      memory[21868] <=  8'h00;      memory[21869] <=  8'h00;      memory[21870] <=  8'h00;      memory[21871] <=  8'h00;      memory[21872] <=  8'h00;      memory[21873] <=  8'h00;      memory[21874] <=  8'h00;      memory[21875] <=  8'h00;      memory[21876] <=  8'h00;      memory[21877] <=  8'h00;      memory[21878] <=  8'h00;      memory[21879] <=  8'h00;      memory[21880] <=  8'h00;      memory[21881] <=  8'h00;      memory[21882] <=  8'h00;      memory[21883] <=  8'h00;      memory[21884] <=  8'h00;      memory[21885] <=  8'h00;      memory[21886] <=  8'h00;      memory[21887] <=  8'h00;      memory[21888] <=  8'h00;      memory[21889] <=  8'h00;      memory[21890] <=  8'h00;      memory[21891] <=  8'h00;      memory[21892] <=  8'h00;      memory[21893] <=  8'h00;      memory[21894] <=  8'h00;      memory[21895] <=  8'h00;      memory[21896] <=  8'h00;      memory[21897] <=  8'h00;      memory[21898] <=  8'h00;      memory[21899] <=  8'h00;      memory[21900] <=  8'h00;      memory[21901] <=  8'h00;      memory[21902] <=  8'h00;      memory[21903] <=  8'h00;      memory[21904] <=  8'h00;      memory[21905] <=  8'h00;      memory[21906] <=  8'h00;      memory[21907] <=  8'h00;      memory[21908] <=  8'h00;      memory[21909] <=  8'h00;      memory[21910] <=  8'h00;      memory[21911] <=  8'h00;      memory[21912] <=  8'h00;      memory[21913] <=  8'h00;      memory[21914] <=  8'h00;      memory[21915] <=  8'h00;      memory[21916] <=  8'h00;      memory[21917] <=  8'h00;      memory[21918] <=  8'h00;      memory[21919] <=  8'h00;      memory[21920] <=  8'h00;      memory[21921] <=  8'h00;      memory[21922] <=  8'h00;      memory[21923] <=  8'h00;      memory[21924] <=  8'h00;      memory[21925] <=  8'h00;      memory[21926] <=  8'h00;      memory[21927] <=  8'h00;      memory[21928] <=  8'h00;      memory[21929] <=  8'h00;      memory[21930] <=  8'h00;      memory[21931] <=  8'h00;      memory[21932] <=  8'h00;      memory[21933] <=  8'h00;      memory[21934] <=  8'h00;      memory[21935] <=  8'h00;      memory[21936] <=  8'h00;      memory[21937] <=  8'h00;      memory[21938] <=  8'h00;      memory[21939] <=  8'h00;      memory[21940] <=  8'h00;      memory[21941] <=  8'h00;      memory[21942] <=  8'h00;      memory[21943] <=  8'h00;      memory[21944] <=  8'h00;      memory[21945] <=  8'h00;      memory[21946] <=  8'h00;      memory[21947] <=  8'h00;      memory[21948] <=  8'h00;      memory[21949] <=  8'h00;      memory[21950] <=  8'h00;      memory[21951] <=  8'h00;      memory[21952] <=  8'h00;      memory[21953] <=  8'h00;      memory[21954] <=  8'h00;      memory[21955] <=  8'h00;      memory[21956] <=  8'h00;      memory[21957] <=  8'h00;      memory[21958] <=  8'h00;      memory[21959] <=  8'h00;      memory[21960] <=  8'h00;      memory[21961] <=  8'h00;      memory[21962] <=  8'h00;      memory[21963] <=  8'h00;      memory[21964] <=  8'h00;      memory[21965] <=  8'h00;      memory[21966] <=  8'h00;      memory[21967] <=  8'h00;      memory[21968] <=  8'h00;      memory[21969] <=  8'h00;      memory[21970] <=  8'h00;      memory[21971] <=  8'h00;      memory[21972] <=  8'h00;      memory[21973] <=  8'h00;      memory[21974] <=  8'h00;      memory[21975] <=  8'h00;      memory[21976] <=  8'h00;      memory[21977] <=  8'h00;      memory[21978] <=  8'h00;      memory[21979] <=  8'h00;      memory[21980] <=  8'h00;      memory[21981] <=  8'h00;      memory[21982] <=  8'h00;      memory[21983] <=  8'h00;      memory[21984] <=  8'h00;      memory[21985] <=  8'h00;      memory[21986] <=  8'h00;      memory[21987] <=  8'h00;      memory[21988] <=  8'h00;      memory[21989] <=  8'h00;      memory[21990] <=  8'h00;      memory[21991] <=  8'h00;      memory[21992] <=  8'h00;      memory[21993] <=  8'h00;      memory[21994] <=  8'h00;      memory[21995] <=  8'h00;      memory[21996] <=  8'h00;      memory[21997] <=  8'h00;      memory[21998] <=  8'h00;      memory[21999] <=  8'h00;      memory[22000] <=  8'h00;      memory[22001] <=  8'h00;      memory[22002] <=  8'h00;      memory[22003] <=  8'h00;      memory[22004] <=  8'h00;      memory[22005] <=  8'h00;      memory[22006] <=  8'h00;      memory[22007] <=  8'h00;      memory[22008] <=  8'h00;      memory[22009] <=  8'h00;      memory[22010] <=  8'h00;      memory[22011] <=  8'h00;      memory[22012] <=  8'h00;      memory[22013] <=  8'h00;      memory[22014] <=  8'h00;      memory[22015] <=  8'h00;      memory[22016] <=  8'h00;      memory[22017] <=  8'h00;      memory[22018] <=  8'h00;      memory[22019] <=  8'h00;      memory[22020] <=  8'h00;      memory[22021] <=  8'h00;      memory[22022] <=  8'h00;      memory[22023] <=  8'h00;      memory[22024] <=  8'h00;      memory[22025] <=  8'h00;      memory[22026] <=  8'h00;      memory[22027] <=  8'h00;      memory[22028] <=  8'h00;      memory[22029] <=  8'h00;      memory[22030] <=  8'h00;      memory[22031] <=  8'h00;      memory[22032] <=  8'h00;      memory[22033] <=  8'h00;      memory[22034] <=  8'h00;      memory[22035] <=  8'h00;      memory[22036] <=  8'h00;      memory[22037] <=  8'h00;      memory[22038] <=  8'h00;      memory[22039] <=  8'h00;      memory[22040] <=  8'h00;      memory[22041] <=  8'h00;      memory[22042] <=  8'h00;      memory[22043] <=  8'h00;      memory[22044] <=  8'h00;      memory[22045] <=  8'h00;      memory[22046] <=  8'h00;      memory[22047] <=  8'h00;      memory[22048] <=  8'h00;      memory[22049] <=  8'h00;      memory[22050] <=  8'h00;      memory[22051] <=  8'h00;      memory[22052] <=  8'h00;      memory[22053] <=  8'h00;      memory[22054] <=  8'h00;      memory[22055] <=  8'h00;      memory[22056] <=  8'h00;      memory[22057] <=  8'h00;      memory[22058] <=  8'h00;      memory[22059] <=  8'h00;      memory[22060] <=  8'h00;      memory[22061] <=  8'h00;      memory[22062] <=  8'h00;      memory[22063] <=  8'h00;      memory[22064] <=  8'h00;      memory[22065] <=  8'h00;      memory[22066] <=  8'h00;      memory[22067] <=  8'h00;      memory[22068] <=  8'h00;      memory[22069] <=  8'h00;      memory[22070] <=  8'h00;      memory[22071] <=  8'h00;      memory[22072] <=  8'h00;      memory[22073] <=  8'h00;      memory[22074] <=  8'h00;      memory[22075] <=  8'h00;      memory[22076] <=  8'h00;      memory[22077] <=  8'h00;      memory[22078] <=  8'h00;      memory[22079] <=  8'h00;      memory[22080] <=  8'h00;      memory[22081] <=  8'h00;      memory[22082] <=  8'h00;      memory[22083] <=  8'h00;      memory[22084] <=  8'h00;      memory[22085] <=  8'h00;      memory[22086] <=  8'h00;      memory[22087] <=  8'h00;      memory[22088] <=  8'h00;      memory[22089] <=  8'h00;      memory[22090] <=  8'h00;      memory[22091] <=  8'h00;      memory[22092] <=  8'h00;      memory[22093] <=  8'h00;      memory[22094] <=  8'h00;      memory[22095] <=  8'h00;      memory[22096] <=  8'h00;      memory[22097] <=  8'h00;      memory[22098] <=  8'h00;      memory[22099] <=  8'h00;      memory[22100] <=  8'h00;      memory[22101] <=  8'h00;      memory[22102] <=  8'h00;      memory[22103] <=  8'h00;      memory[22104] <=  8'h00;      memory[22105] <=  8'h00;      memory[22106] <=  8'h00;      memory[22107] <=  8'h00;      memory[22108] <=  8'h00;      memory[22109] <=  8'h00;      memory[22110] <=  8'h00;      memory[22111] <=  8'h00;      memory[22112] <=  8'h00;      memory[22113] <=  8'h00;      memory[22114] <=  8'h00;      memory[22115] <=  8'h00;      memory[22116] <=  8'h00;      memory[22117] <=  8'h00;      memory[22118] <=  8'h00;      memory[22119] <=  8'h00;      memory[22120] <=  8'h00;      memory[22121] <=  8'h00;      memory[22122] <=  8'h00;      memory[22123] <=  8'h00;      memory[22124] <=  8'h00;      memory[22125] <=  8'h00;      memory[22126] <=  8'h00;      memory[22127] <=  8'h00;      memory[22128] <=  8'h00;      memory[22129] <=  8'h00;      memory[22130] <=  8'h00;      memory[22131] <=  8'h00;      memory[22132] <=  8'h00;      memory[22133] <=  8'h00;      memory[22134] <=  8'h00;      memory[22135] <=  8'h00;      memory[22136] <=  8'h00;      memory[22137] <=  8'h00;      memory[22138] <=  8'h00;      memory[22139] <=  8'h00;      memory[22140] <=  8'h00;      memory[22141] <=  8'h00;      memory[22142] <=  8'h00;      memory[22143] <=  8'h00;      memory[22144] <=  8'h00;      memory[22145] <=  8'h00;      memory[22146] <=  8'h00;      memory[22147] <=  8'h00;      memory[22148] <=  8'h00;      memory[22149] <=  8'h00;      memory[22150] <=  8'h00;      memory[22151] <=  8'h00;      memory[22152] <=  8'h00;      memory[22153] <=  8'h00;      memory[22154] <=  8'h00;      memory[22155] <=  8'h00;      memory[22156] <=  8'h00;      memory[22157] <=  8'h00;      memory[22158] <=  8'h00;      memory[22159] <=  8'h00;      memory[22160] <=  8'h00;      memory[22161] <=  8'h00;      memory[22162] <=  8'h00;      memory[22163] <=  8'h00;      memory[22164] <=  8'h00;      memory[22165] <=  8'h00;      memory[22166] <=  8'h00;      memory[22167] <=  8'h00;      memory[22168] <=  8'h00;      memory[22169] <=  8'h00;      memory[22170] <=  8'h00;      memory[22171] <=  8'h00;      memory[22172] <=  8'h00;      memory[22173] <=  8'h00;      memory[22174] <=  8'h00;      memory[22175] <=  8'h00;      memory[22176] <=  8'h00;      memory[22177] <=  8'h00;      memory[22178] <=  8'h00;      memory[22179] <=  8'h00;      memory[22180] <=  8'h00;      memory[22181] <=  8'h00;      memory[22182] <=  8'h00;      memory[22183] <=  8'h00;      memory[22184] <=  8'h00;      memory[22185] <=  8'h00;      memory[22186] <=  8'h00;      memory[22187] <=  8'h00;      memory[22188] <=  8'h00;      memory[22189] <=  8'h00;      memory[22190] <=  8'h00;      memory[22191] <=  8'h00;      memory[22192] <=  8'h00;      memory[22193] <=  8'h00;      memory[22194] <=  8'h00;      memory[22195] <=  8'h00;      memory[22196] <=  8'h00;      memory[22197] <=  8'h00;      memory[22198] <=  8'h00;      memory[22199] <=  8'h00;      memory[22200] <=  8'h00;      memory[22201] <=  8'h00;      memory[22202] <=  8'h00;      memory[22203] <=  8'h00;      memory[22204] <=  8'h00;      memory[22205] <=  8'h00;      memory[22206] <=  8'h00;      memory[22207] <=  8'h00;      memory[22208] <=  8'h00;      memory[22209] <=  8'h00;      memory[22210] <=  8'h00;      memory[22211] <=  8'h00;      memory[22212] <=  8'h00;      memory[22213] <=  8'h00;      memory[22214] <=  8'h00;      memory[22215] <=  8'h00;      memory[22216] <=  8'h00;      memory[22217] <=  8'h00;      memory[22218] <=  8'h00;      memory[22219] <=  8'h00;      memory[22220] <=  8'h00;      memory[22221] <=  8'h00;      memory[22222] <=  8'h00;      memory[22223] <=  8'h00;      memory[22224] <=  8'h00;      memory[22225] <=  8'h00;      memory[22226] <=  8'h00;      memory[22227] <=  8'h00;      memory[22228] <=  8'h00;      memory[22229] <=  8'h00;      memory[22230] <=  8'h00;      memory[22231] <=  8'h00;      memory[22232] <=  8'h00;      memory[22233] <=  8'h00;      memory[22234] <=  8'h00;      memory[22235] <=  8'h00;      memory[22236] <=  8'h00;      memory[22237] <=  8'h00;      memory[22238] <=  8'h00;      memory[22239] <=  8'h00;      memory[22240] <=  8'h00;      memory[22241] <=  8'h00;      memory[22242] <=  8'h00;      memory[22243] <=  8'h00;      memory[22244] <=  8'h00;      memory[22245] <=  8'h00;      memory[22246] <=  8'h00;      memory[22247] <=  8'h00;      memory[22248] <=  8'h00;      memory[22249] <=  8'h00;      memory[22250] <=  8'h00;      memory[22251] <=  8'h00;      memory[22252] <=  8'h00;      memory[22253] <=  8'h00;      memory[22254] <=  8'h00;      memory[22255] <=  8'h00;      memory[22256] <=  8'h00;      memory[22257] <=  8'h00;      memory[22258] <=  8'h00;      memory[22259] <=  8'h00;      memory[22260] <=  8'h00;      memory[22261] <=  8'h00;      memory[22262] <=  8'h00;      memory[22263] <=  8'h00;      memory[22264] <=  8'h00;      memory[22265] <=  8'h00;      memory[22266] <=  8'h00;      memory[22267] <=  8'h00;      memory[22268] <=  8'h00;      memory[22269] <=  8'h00;      memory[22270] <=  8'h00;      memory[22271] <=  8'h00;      memory[22272] <=  8'h00;      memory[22273] <=  8'h00;      memory[22274] <=  8'h00;      memory[22275] <=  8'h00;      memory[22276] <=  8'h00;      memory[22277] <=  8'h00;      memory[22278] <=  8'h00;      memory[22279] <=  8'h00;      memory[22280] <=  8'h00;      memory[22281] <=  8'h00;      memory[22282] <=  8'h00;      memory[22283] <=  8'h00;      memory[22284] <=  8'h00;      memory[22285] <=  8'h00;      memory[22286] <=  8'h00;      memory[22287] <=  8'h00;      memory[22288] <=  8'h00;      memory[22289] <=  8'h00;      memory[22290] <=  8'h00;      memory[22291] <=  8'h00;      memory[22292] <=  8'h00;      memory[22293] <=  8'h00;      memory[22294] <=  8'h00;      memory[22295] <=  8'h00;      memory[22296] <=  8'h00;      memory[22297] <=  8'h00;      memory[22298] <=  8'h00;      memory[22299] <=  8'h00;      memory[22300] <=  8'h00;      memory[22301] <=  8'h00;      memory[22302] <=  8'h00;      memory[22303] <=  8'h00;      memory[22304] <=  8'h00;      memory[22305] <=  8'h00;      memory[22306] <=  8'h00;      memory[22307] <=  8'h00;      memory[22308] <=  8'h00;      memory[22309] <=  8'h00;      memory[22310] <=  8'h00;      memory[22311] <=  8'h00;      memory[22312] <=  8'h00;      memory[22313] <=  8'h00;      memory[22314] <=  8'h00;      memory[22315] <=  8'h00;      memory[22316] <=  8'h00;      memory[22317] <=  8'h00;      memory[22318] <=  8'h00;      memory[22319] <=  8'h00;      memory[22320] <=  8'h00;      memory[22321] <=  8'h00;      memory[22322] <=  8'h00;      memory[22323] <=  8'h00;      memory[22324] <=  8'h00;      memory[22325] <=  8'h00;      memory[22326] <=  8'h00;      memory[22327] <=  8'h00;      memory[22328] <=  8'h00;      memory[22329] <=  8'h00;      memory[22330] <=  8'h00;      memory[22331] <=  8'h00;      memory[22332] <=  8'h00;      memory[22333] <=  8'h00;      memory[22334] <=  8'h00;      memory[22335] <=  8'h00;      memory[22336] <=  8'h00;      memory[22337] <=  8'h00;      memory[22338] <=  8'h00;      memory[22339] <=  8'h00;      memory[22340] <=  8'h00;      memory[22341] <=  8'h00;      memory[22342] <=  8'h00;      memory[22343] <=  8'h00;      memory[22344] <=  8'h00;      memory[22345] <=  8'h00;      memory[22346] <=  8'h00;      memory[22347] <=  8'h00;      memory[22348] <=  8'h00;      memory[22349] <=  8'h00;      memory[22350] <=  8'h00;      memory[22351] <=  8'h00;      memory[22352] <=  8'h00;      memory[22353] <=  8'h00;      memory[22354] <=  8'h00;      memory[22355] <=  8'h00;      memory[22356] <=  8'h00;      memory[22357] <=  8'h00;      memory[22358] <=  8'h00;      memory[22359] <=  8'h00;      memory[22360] <=  8'h00;      memory[22361] <=  8'h00;      memory[22362] <=  8'h00;      memory[22363] <=  8'h00;      memory[22364] <=  8'h00;      memory[22365] <=  8'h00;      memory[22366] <=  8'h00;      memory[22367] <=  8'h00;      memory[22368] <=  8'h00;      memory[22369] <=  8'h00;      memory[22370] <=  8'h00;      memory[22371] <=  8'h00;      memory[22372] <=  8'h00;      memory[22373] <=  8'h00;      memory[22374] <=  8'h00;      memory[22375] <=  8'h00;      memory[22376] <=  8'h00;      memory[22377] <=  8'h00;      memory[22378] <=  8'h00;      memory[22379] <=  8'h00;      memory[22380] <=  8'h00;      memory[22381] <=  8'h00;      memory[22382] <=  8'h00;      memory[22383] <=  8'h00;      memory[22384] <=  8'h00;      memory[22385] <=  8'h00;      memory[22386] <=  8'h00;      memory[22387] <=  8'h00;      memory[22388] <=  8'h00;      memory[22389] <=  8'h00;      memory[22390] <=  8'h00;      memory[22391] <=  8'h00;      memory[22392] <=  8'h00;      memory[22393] <=  8'h00;      memory[22394] <=  8'h00;      memory[22395] <=  8'h00;      memory[22396] <=  8'h00;      memory[22397] <=  8'h00;      memory[22398] <=  8'h00;      memory[22399] <=  8'h00;      memory[22400] <=  8'h00;      memory[22401] <=  8'h00;      memory[22402] <=  8'h00;      memory[22403] <=  8'h00;      memory[22404] <=  8'h00;      memory[22405] <=  8'h00;      memory[22406] <=  8'h00;      memory[22407] <=  8'h00;      memory[22408] <=  8'h00;      memory[22409] <=  8'h00;      memory[22410] <=  8'h00;      memory[22411] <=  8'h00;      memory[22412] <=  8'h00;      memory[22413] <=  8'h00;      memory[22414] <=  8'h00;      memory[22415] <=  8'h00;      memory[22416] <=  8'h00;      memory[22417] <=  8'h00;      memory[22418] <=  8'h00;      memory[22419] <=  8'h00;      memory[22420] <=  8'h00;      memory[22421] <=  8'h00;      memory[22422] <=  8'h00;      memory[22423] <=  8'h00;      memory[22424] <=  8'h00;      memory[22425] <=  8'h00;      memory[22426] <=  8'h00;      memory[22427] <=  8'h00;      memory[22428] <=  8'h00;      memory[22429] <=  8'h00;      memory[22430] <=  8'h00;      memory[22431] <=  8'h00;      memory[22432] <=  8'h00;      memory[22433] <=  8'h00;      memory[22434] <=  8'h00;      memory[22435] <=  8'h00;      memory[22436] <=  8'h00;      memory[22437] <=  8'h00;      memory[22438] <=  8'h00;      memory[22439] <=  8'h00;      memory[22440] <=  8'h00;      memory[22441] <=  8'h00;      memory[22442] <=  8'h00;      memory[22443] <=  8'h00;      memory[22444] <=  8'h00;      memory[22445] <=  8'h00;      memory[22446] <=  8'h00;      memory[22447] <=  8'h00;      memory[22448] <=  8'h00;      memory[22449] <=  8'h00;      memory[22450] <=  8'h00;      memory[22451] <=  8'h00;      memory[22452] <=  8'h00;      memory[22453] <=  8'h00;      memory[22454] <=  8'h00;      memory[22455] <=  8'h00;      memory[22456] <=  8'h00;      memory[22457] <=  8'h00;      memory[22458] <=  8'h00;      memory[22459] <=  8'h00;      memory[22460] <=  8'h00;      memory[22461] <=  8'h00;      memory[22462] <=  8'h00;      memory[22463] <=  8'h00;      memory[22464] <=  8'h00;      memory[22465] <=  8'h00;      memory[22466] <=  8'h00;      memory[22467] <=  8'h00;      memory[22468] <=  8'h00;      memory[22469] <=  8'h00;      memory[22470] <=  8'h00;      memory[22471] <=  8'h00;      memory[22472] <=  8'h00;      memory[22473] <=  8'h00;      memory[22474] <=  8'h00;      memory[22475] <=  8'h00;      memory[22476] <=  8'h00;      memory[22477] <=  8'h00;      memory[22478] <=  8'h00;      memory[22479] <=  8'h00;      memory[22480] <=  8'h00;      memory[22481] <=  8'h00;      memory[22482] <=  8'h00;      memory[22483] <=  8'h00;      memory[22484] <=  8'h00;      memory[22485] <=  8'h00;      memory[22486] <=  8'h00;      memory[22487] <=  8'h00;      memory[22488] <=  8'h00;      memory[22489] <=  8'h00;      memory[22490] <=  8'h00;      memory[22491] <=  8'h00;      memory[22492] <=  8'h00;      memory[22493] <=  8'h00;      memory[22494] <=  8'h00;      memory[22495] <=  8'h00;      memory[22496] <=  8'h00;      memory[22497] <=  8'h00;      memory[22498] <=  8'h00;      memory[22499] <=  8'h00;      memory[22500] <=  8'h00;      memory[22501] <=  8'h00;      memory[22502] <=  8'h00;      memory[22503] <=  8'h00;      memory[22504] <=  8'h00;      memory[22505] <=  8'h00;      memory[22506] <=  8'h00;      memory[22507] <=  8'h00;      memory[22508] <=  8'h00;      memory[22509] <=  8'h00;      memory[22510] <=  8'h00;      memory[22511] <=  8'h00;      memory[22512] <=  8'h00;      memory[22513] <=  8'h00;      memory[22514] <=  8'h00;      memory[22515] <=  8'h00;      memory[22516] <=  8'h00;      memory[22517] <=  8'h00;      memory[22518] <=  8'h00;      memory[22519] <=  8'h00;      memory[22520] <=  8'h00;      memory[22521] <=  8'h00;      memory[22522] <=  8'h00;      memory[22523] <=  8'h00;      memory[22524] <=  8'h00;      memory[22525] <=  8'h00;      memory[22526] <=  8'h00;      memory[22527] <=  8'h00;      memory[22528] <=  8'h00;      memory[22529] <=  8'h00;      memory[22530] <=  8'h00;      memory[22531] <=  8'h00;      memory[22532] <=  8'h00;      memory[22533] <=  8'h00;      memory[22534] <=  8'h00;      memory[22535] <=  8'h00;      memory[22536] <=  8'h00;      memory[22537] <=  8'h00;      memory[22538] <=  8'h00;      memory[22539] <=  8'h00;      memory[22540] <=  8'h00;      memory[22541] <=  8'h00;      memory[22542] <=  8'h00;      memory[22543] <=  8'h00;      memory[22544] <=  8'h00;      memory[22545] <=  8'h00;      memory[22546] <=  8'h00;      memory[22547] <=  8'h00;      memory[22548] <=  8'h00;      memory[22549] <=  8'h00;      memory[22550] <=  8'h00;      memory[22551] <=  8'h00;      memory[22552] <=  8'h00;      memory[22553] <=  8'h00;      memory[22554] <=  8'h00;      memory[22555] <=  8'h00;      memory[22556] <=  8'h00;      memory[22557] <=  8'h00;      memory[22558] <=  8'h00;      memory[22559] <=  8'h00;      memory[22560] <=  8'h00;      memory[22561] <=  8'h00;      memory[22562] <=  8'h00;      memory[22563] <=  8'h00;      memory[22564] <=  8'h00;      memory[22565] <=  8'h00;      memory[22566] <=  8'h00;      memory[22567] <=  8'h00;      memory[22568] <=  8'h00;      memory[22569] <=  8'h00;      memory[22570] <=  8'h00;      memory[22571] <=  8'h00;      memory[22572] <=  8'h00;      memory[22573] <=  8'h00;      memory[22574] <=  8'h00;      memory[22575] <=  8'h00;      memory[22576] <=  8'h00;      memory[22577] <=  8'h00;      memory[22578] <=  8'h00;      memory[22579] <=  8'h00;      memory[22580] <=  8'h00;      memory[22581] <=  8'h00;      memory[22582] <=  8'h00;      memory[22583] <=  8'h00;      memory[22584] <=  8'h00;      memory[22585] <=  8'h00;      memory[22586] <=  8'h00;      memory[22587] <=  8'h00;      memory[22588] <=  8'h00;      memory[22589] <=  8'h00;      memory[22590] <=  8'h00;      memory[22591] <=  8'h00;      memory[22592] <=  8'h00;      memory[22593] <=  8'h00;      memory[22594] <=  8'h00;      memory[22595] <=  8'h00;      memory[22596] <=  8'h00;      memory[22597] <=  8'h00;      memory[22598] <=  8'h00;      memory[22599] <=  8'h00;      memory[22600] <=  8'h00;      memory[22601] <=  8'h00;      memory[22602] <=  8'h00;      memory[22603] <=  8'h00;      memory[22604] <=  8'h00;      memory[22605] <=  8'h00;      memory[22606] <=  8'h00;      memory[22607] <=  8'h00;      memory[22608] <=  8'h00;      memory[22609] <=  8'h00;      memory[22610] <=  8'h00;      memory[22611] <=  8'h00;      memory[22612] <=  8'h00;      memory[22613] <=  8'h00;      memory[22614] <=  8'h00;      memory[22615] <=  8'h00;      memory[22616] <=  8'h00;      memory[22617] <=  8'h00;      memory[22618] <=  8'h00;      memory[22619] <=  8'h00;      memory[22620] <=  8'h00;      memory[22621] <=  8'h00;      memory[22622] <=  8'h00;      memory[22623] <=  8'h00;      memory[22624] <=  8'h00;      memory[22625] <=  8'h00;      memory[22626] <=  8'h00;      memory[22627] <=  8'h00;      memory[22628] <=  8'h00;      memory[22629] <=  8'h00;      memory[22630] <=  8'h00;      memory[22631] <=  8'h00;      memory[22632] <=  8'h00;      memory[22633] <=  8'h00;      memory[22634] <=  8'h00;      memory[22635] <=  8'h00;      memory[22636] <=  8'h00;      memory[22637] <=  8'h00;      memory[22638] <=  8'h00;      memory[22639] <=  8'h00;      memory[22640] <=  8'h00;      memory[22641] <=  8'h00;      memory[22642] <=  8'h00;      memory[22643] <=  8'h00;      memory[22644] <=  8'h00;      memory[22645] <=  8'h00;      memory[22646] <=  8'h00;      memory[22647] <=  8'h00;      memory[22648] <=  8'h00;      memory[22649] <=  8'h00;      memory[22650] <=  8'h00;      memory[22651] <=  8'h00;      memory[22652] <=  8'h00;      memory[22653] <=  8'h00;      memory[22654] <=  8'h00;      memory[22655] <=  8'h00;      memory[22656] <=  8'h00;      memory[22657] <=  8'h00;      memory[22658] <=  8'h00;      memory[22659] <=  8'h00;      memory[22660] <=  8'h00;      memory[22661] <=  8'h00;      memory[22662] <=  8'h00;      memory[22663] <=  8'h00;      memory[22664] <=  8'h00;      memory[22665] <=  8'h00;      memory[22666] <=  8'h00;      memory[22667] <=  8'h00;      memory[22668] <=  8'h00;      memory[22669] <=  8'h00;      memory[22670] <=  8'h00;      memory[22671] <=  8'h00;      memory[22672] <=  8'h00;      memory[22673] <=  8'h00;      memory[22674] <=  8'h00;      memory[22675] <=  8'h00;      memory[22676] <=  8'h00;      memory[22677] <=  8'h00;      memory[22678] <=  8'h00;      memory[22679] <=  8'h00;      memory[22680] <=  8'h00;      memory[22681] <=  8'h00;      memory[22682] <=  8'h00;      memory[22683] <=  8'h00;      memory[22684] <=  8'h00;      memory[22685] <=  8'h00;      memory[22686] <=  8'h00;      memory[22687] <=  8'h00;      memory[22688] <=  8'h00;      memory[22689] <=  8'h00;      memory[22690] <=  8'h00;      memory[22691] <=  8'h00;      memory[22692] <=  8'h00;      memory[22693] <=  8'h00;      memory[22694] <=  8'h00;      memory[22695] <=  8'h00;      memory[22696] <=  8'h00;      memory[22697] <=  8'h00;      memory[22698] <=  8'h00;      memory[22699] <=  8'h00;      memory[22700] <=  8'h00;      memory[22701] <=  8'h00;      memory[22702] <=  8'h00;      memory[22703] <=  8'h00;      memory[22704] <=  8'h00;      memory[22705] <=  8'h00;      memory[22706] <=  8'h00;      memory[22707] <=  8'h00;      memory[22708] <=  8'h00;      memory[22709] <=  8'h00;      memory[22710] <=  8'h00;      memory[22711] <=  8'h00;      memory[22712] <=  8'h00;      memory[22713] <=  8'h00;      memory[22714] <=  8'h00;      memory[22715] <=  8'h00;      memory[22716] <=  8'h00;      memory[22717] <=  8'h00;      memory[22718] <=  8'h00;      memory[22719] <=  8'h00;      memory[22720] <=  8'h00;      memory[22721] <=  8'h00;      memory[22722] <=  8'h00;      memory[22723] <=  8'h00;      memory[22724] <=  8'h00;      memory[22725] <=  8'h00;      memory[22726] <=  8'h00;      memory[22727] <=  8'h00;      memory[22728] <=  8'h00;      memory[22729] <=  8'h00;      memory[22730] <=  8'h00;      memory[22731] <=  8'h00;      memory[22732] <=  8'h00;      memory[22733] <=  8'h00;      memory[22734] <=  8'h00;      memory[22735] <=  8'h00;      memory[22736] <=  8'h00;      memory[22737] <=  8'h00;      memory[22738] <=  8'h00;      memory[22739] <=  8'h00;      memory[22740] <=  8'h00;      memory[22741] <=  8'h00;      memory[22742] <=  8'h00;      memory[22743] <=  8'h00;      memory[22744] <=  8'h00;      memory[22745] <=  8'h00;      memory[22746] <=  8'h00;      memory[22747] <=  8'h00;      memory[22748] <=  8'h00;      memory[22749] <=  8'h00;      memory[22750] <=  8'h00;      memory[22751] <=  8'h00;      memory[22752] <=  8'h00;      memory[22753] <=  8'h00;      memory[22754] <=  8'h00;      memory[22755] <=  8'h00;      memory[22756] <=  8'h00;      memory[22757] <=  8'h00;      memory[22758] <=  8'h00;      memory[22759] <=  8'h00;      memory[22760] <=  8'h00;      memory[22761] <=  8'h00;      memory[22762] <=  8'h00;      memory[22763] <=  8'h00;      memory[22764] <=  8'h00;      memory[22765] <=  8'h00;      memory[22766] <=  8'h00;      memory[22767] <=  8'h00;      memory[22768] <=  8'h00;      memory[22769] <=  8'h00;      memory[22770] <=  8'h00;      memory[22771] <=  8'h00;      memory[22772] <=  8'h00;      memory[22773] <=  8'h00;      memory[22774] <=  8'h00;      memory[22775] <=  8'h00;      memory[22776] <=  8'h00;      memory[22777] <=  8'h00;      memory[22778] <=  8'h00;      memory[22779] <=  8'h00;      memory[22780] <=  8'h00;      memory[22781] <=  8'h00;      memory[22782] <=  8'h00;      memory[22783] <=  8'h00;      memory[22784] <=  8'h00;      memory[22785] <=  8'h00;      memory[22786] <=  8'h00;      memory[22787] <=  8'h00;      memory[22788] <=  8'h00;      memory[22789] <=  8'h00;      memory[22790] <=  8'h00;      memory[22791] <=  8'h00;      memory[22792] <=  8'h00;      memory[22793] <=  8'h00;      memory[22794] <=  8'h00;      memory[22795] <=  8'h00;      memory[22796] <=  8'h00;      memory[22797] <=  8'h00;      memory[22798] <=  8'h00;      memory[22799] <=  8'h00;      memory[22800] <=  8'h00;      memory[22801] <=  8'h00;      memory[22802] <=  8'h00;      memory[22803] <=  8'h00;      memory[22804] <=  8'h00;      memory[22805] <=  8'h00;      memory[22806] <=  8'h00;      memory[22807] <=  8'h00;      memory[22808] <=  8'h00;      memory[22809] <=  8'h00;      memory[22810] <=  8'h00;      memory[22811] <=  8'h00;      memory[22812] <=  8'h00;      memory[22813] <=  8'h00;      memory[22814] <=  8'h00;      memory[22815] <=  8'h00;      memory[22816] <=  8'h00;      memory[22817] <=  8'h00;      memory[22818] <=  8'h00;      memory[22819] <=  8'h00;      memory[22820] <=  8'h00;      memory[22821] <=  8'h00;      memory[22822] <=  8'h00;      memory[22823] <=  8'h00;      memory[22824] <=  8'h00;      memory[22825] <=  8'h00;      memory[22826] <=  8'h00;      memory[22827] <=  8'h00;      memory[22828] <=  8'h00;      memory[22829] <=  8'h00;      memory[22830] <=  8'h00;      memory[22831] <=  8'h00;      memory[22832] <=  8'h00;      memory[22833] <=  8'h00;      memory[22834] <=  8'h00;      memory[22835] <=  8'h00;      memory[22836] <=  8'h00;      memory[22837] <=  8'h00;      memory[22838] <=  8'h00;      memory[22839] <=  8'h00;      memory[22840] <=  8'h00;      memory[22841] <=  8'h00;      memory[22842] <=  8'h00;      memory[22843] <=  8'h00;      memory[22844] <=  8'h00;      memory[22845] <=  8'h00;      memory[22846] <=  8'h00;      memory[22847] <=  8'h00;      memory[22848] <=  8'h00;      memory[22849] <=  8'h00;      memory[22850] <=  8'h00;      memory[22851] <=  8'h00;      memory[22852] <=  8'h00;      memory[22853] <=  8'h00;      memory[22854] <=  8'h00;      memory[22855] <=  8'h00;      memory[22856] <=  8'h00;      memory[22857] <=  8'h00;      memory[22858] <=  8'h00;      memory[22859] <=  8'h00;      memory[22860] <=  8'h00;      memory[22861] <=  8'h00;      memory[22862] <=  8'h00;      memory[22863] <=  8'h00;      memory[22864] <=  8'h00;      memory[22865] <=  8'h00;      memory[22866] <=  8'h00;      memory[22867] <=  8'h00;      memory[22868] <=  8'h00;      memory[22869] <=  8'h00;      memory[22870] <=  8'h00;      memory[22871] <=  8'h00;      memory[22872] <=  8'h00;      memory[22873] <=  8'h00;      memory[22874] <=  8'h00;      memory[22875] <=  8'h00;      memory[22876] <=  8'h00;      memory[22877] <=  8'h00;      memory[22878] <=  8'h00;      memory[22879] <=  8'h00;      memory[22880] <=  8'h00;      memory[22881] <=  8'h00;      memory[22882] <=  8'h00;      memory[22883] <=  8'h00;      memory[22884] <=  8'h00;      memory[22885] <=  8'h00;      memory[22886] <=  8'h00;      memory[22887] <=  8'h00;      memory[22888] <=  8'h00;      memory[22889] <=  8'h00;      memory[22890] <=  8'h00;      memory[22891] <=  8'h00;      memory[22892] <=  8'h00;      memory[22893] <=  8'h00;      memory[22894] <=  8'h00;      memory[22895] <=  8'h00;      memory[22896] <=  8'h00;      memory[22897] <=  8'h00;      memory[22898] <=  8'h00;      memory[22899] <=  8'h00;      memory[22900] <=  8'h00;      memory[22901] <=  8'h00;      memory[22902] <=  8'h00;      memory[22903] <=  8'h00;      memory[22904] <=  8'h00;      memory[22905] <=  8'h00;      memory[22906] <=  8'h00;      memory[22907] <=  8'h00;      memory[22908] <=  8'h00;      memory[22909] <=  8'h00;      memory[22910] <=  8'h00;      memory[22911] <=  8'h00;      memory[22912] <=  8'h00;      memory[22913] <=  8'h00;      memory[22914] <=  8'h00;      memory[22915] <=  8'h00;      memory[22916] <=  8'h00;      memory[22917] <=  8'h00;      memory[22918] <=  8'h00;      memory[22919] <=  8'h00;      memory[22920] <=  8'h00;      memory[22921] <=  8'h00;      memory[22922] <=  8'h00;      memory[22923] <=  8'h00;      memory[22924] <=  8'h00;      memory[22925] <=  8'h00;      memory[22926] <=  8'h00;      memory[22927] <=  8'h00;      memory[22928] <=  8'h00;      memory[22929] <=  8'h00;      memory[22930] <=  8'h00;      memory[22931] <=  8'h00;      memory[22932] <=  8'h00;      memory[22933] <=  8'h00;      memory[22934] <=  8'h00;      memory[22935] <=  8'h00;      memory[22936] <=  8'h00;      memory[22937] <=  8'h00;      memory[22938] <=  8'h00;      memory[22939] <=  8'h00;      memory[22940] <=  8'h00;      memory[22941] <=  8'h00;      memory[22942] <=  8'h00;      memory[22943] <=  8'h00;      memory[22944] <=  8'h00;      memory[22945] <=  8'h00;      memory[22946] <=  8'h00;      memory[22947] <=  8'h00;      memory[22948] <=  8'h00;      memory[22949] <=  8'h00;      memory[22950] <=  8'h00;      memory[22951] <=  8'h00;      memory[22952] <=  8'h00;      memory[22953] <=  8'h00;      memory[22954] <=  8'h00;      memory[22955] <=  8'h00;      memory[22956] <=  8'h00;      memory[22957] <=  8'h00;      memory[22958] <=  8'h00;      memory[22959] <=  8'h00;      memory[22960] <=  8'h00;      memory[22961] <=  8'h00;      memory[22962] <=  8'h00;      memory[22963] <=  8'h00;      memory[22964] <=  8'h00;      memory[22965] <=  8'h00;      memory[22966] <=  8'h00;      memory[22967] <=  8'h00;      memory[22968] <=  8'h00;      memory[22969] <=  8'h00;      memory[22970] <=  8'h00;      memory[22971] <=  8'h00;      memory[22972] <=  8'h00;      memory[22973] <=  8'h00;      memory[22974] <=  8'h00;      memory[22975] <=  8'h00;      memory[22976] <=  8'h00;      memory[22977] <=  8'h00;      memory[22978] <=  8'h00;      memory[22979] <=  8'h00;      memory[22980] <=  8'h00;      memory[22981] <=  8'h00;      memory[22982] <=  8'h00;      memory[22983] <=  8'h00;      memory[22984] <=  8'h00;      memory[22985] <=  8'h00;      memory[22986] <=  8'h00;      memory[22987] <=  8'h00;      memory[22988] <=  8'h00;      memory[22989] <=  8'h00;      memory[22990] <=  8'h00;      memory[22991] <=  8'h00;      memory[22992] <=  8'h00;      memory[22993] <=  8'h00;      memory[22994] <=  8'h00;      memory[22995] <=  8'h00;      memory[22996] <=  8'h00;      memory[22997] <=  8'h00;      memory[22998] <=  8'h00;      memory[22999] <=  8'h00;      memory[23000] <=  8'h00;      memory[23001] <=  8'h00;      memory[23002] <=  8'h00;      memory[23003] <=  8'h00;      memory[23004] <=  8'h00;      memory[23005] <=  8'h00;      memory[23006] <=  8'h00;      memory[23007] <=  8'h00;      memory[23008] <=  8'h00;      memory[23009] <=  8'h00;      memory[23010] <=  8'h00;      memory[23011] <=  8'h00;      memory[23012] <=  8'h00;      memory[23013] <=  8'h00;      memory[23014] <=  8'h00;      memory[23015] <=  8'h00;      memory[23016] <=  8'h00;      memory[23017] <=  8'h00;      memory[23018] <=  8'h00;      memory[23019] <=  8'h00;      memory[23020] <=  8'h00;      memory[23021] <=  8'h00;      memory[23022] <=  8'h00;      memory[23023] <=  8'h00;      memory[23024] <=  8'h00;      memory[23025] <=  8'h00;      memory[23026] <=  8'h00;      memory[23027] <=  8'h00;      memory[23028] <=  8'h00;      memory[23029] <=  8'h00;      memory[23030] <=  8'h00;      memory[23031] <=  8'h00;      memory[23032] <=  8'h00;      memory[23033] <=  8'h00;      memory[23034] <=  8'h00;      memory[23035] <=  8'h00;      memory[23036] <=  8'h00;      memory[23037] <=  8'h00;      memory[23038] <=  8'h00;      memory[23039] <=  8'h00;      memory[23040] <=  8'h00;      memory[23041] <=  8'h00;      memory[23042] <=  8'h00;      memory[23043] <=  8'h00;      memory[23044] <=  8'h00;      memory[23045] <=  8'h00;      memory[23046] <=  8'h00;      memory[23047] <=  8'h00;      memory[23048] <=  8'h00;      memory[23049] <=  8'h00;      memory[23050] <=  8'h00;      memory[23051] <=  8'h00;      memory[23052] <=  8'h00;      memory[23053] <=  8'h00;      memory[23054] <=  8'h00;      memory[23055] <=  8'h00;      memory[23056] <=  8'h00;      memory[23057] <=  8'h00;      memory[23058] <=  8'h00;      memory[23059] <=  8'h00;      memory[23060] <=  8'h00;      memory[23061] <=  8'h00;      memory[23062] <=  8'h00;      memory[23063] <=  8'h00;      memory[23064] <=  8'h00;      memory[23065] <=  8'h00;      memory[23066] <=  8'h00;      memory[23067] <=  8'h00;      memory[23068] <=  8'h00;      memory[23069] <=  8'h00;      memory[23070] <=  8'h00;      memory[23071] <=  8'h00;      memory[23072] <=  8'h00;      memory[23073] <=  8'h00;      memory[23074] <=  8'h00;      memory[23075] <=  8'h00;      memory[23076] <=  8'h00;      memory[23077] <=  8'h00;      memory[23078] <=  8'h00;      memory[23079] <=  8'h00;      memory[23080] <=  8'h00;      memory[23081] <=  8'h00;      memory[23082] <=  8'h00;      memory[23083] <=  8'h00;      memory[23084] <=  8'h00;      memory[23085] <=  8'h00;      memory[23086] <=  8'h00;      memory[23087] <=  8'h00;      memory[23088] <=  8'h00;      memory[23089] <=  8'h00;      memory[23090] <=  8'h00;      memory[23091] <=  8'h00;      memory[23092] <=  8'h00;      memory[23093] <=  8'h00;      memory[23094] <=  8'h00;      memory[23095] <=  8'h00;      memory[23096] <=  8'h00;      memory[23097] <=  8'h00;      memory[23098] <=  8'h00;      memory[23099] <=  8'h00;      memory[23100] <=  8'h00;      memory[23101] <=  8'h00;      memory[23102] <=  8'h00;      memory[23103] <=  8'h00;      memory[23104] <=  8'h00;      memory[23105] <=  8'h00;      memory[23106] <=  8'h00;      memory[23107] <=  8'h00;      memory[23108] <=  8'h00;      memory[23109] <=  8'h00;      memory[23110] <=  8'h00;      memory[23111] <=  8'h00;      memory[23112] <=  8'h00;      memory[23113] <=  8'h00;      memory[23114] <=  8'h00;      memory[23115] <=  8'h00;      memory[23116] <=  8'h00;      memory[23117] <=  8'h00;      memory[23118] <=  8'h00;      memory[23119] <=  8'h00;      memory[23120] <=  8'h00;      memory[23121] <=  8'h00;      memory[23122] <=  8'h00;      memory[23123] <=  8'h00;      memory[23124] <=  8'h00;      memory[23125] <=  8'h00;      memory[23126] <=  8'h00;      memory[23127] <=  8'h00;      memory[23128] <=  8'h00;      memory[23129] <=  8'h00;      memory[23130] <=  8'h00;      memory[23131] <=  8'h00;      memory[23132] <=  8'h00;      memory[23133] <=  8'h00;      memory[23134] <=  8'h00;      memory[23135] <=  8'h00;      memory[23136] <=  8'h00;      memory[23137] <=  8'h00;      memory[23138] <=  8'h00;      memory[23139] <=  8'h00;      memory[23140] <=  8'h00;      memory[23141] <=  8'h00;      memory[23142] <=  8'h00;      memory[23143] <=  8'h00;      memory[23144] <=  8'h00;      memory[23145] <=  8'h00;      memory[23146] <=  8'h00;      memory[23147] <=  8'h00;      memory[23148] <=  8'h00;      memory[23149] <=  8'h00;      memory[23150] <=  8'h00;      memory[23151] <=  8'h00;      memory[23152] <=  8'h00;      memory[23153] <=  8'h00;      memory[23154] <=  8'h00;      memory[23155] <=  8'h00;      memory[23156] <=  8'h00;      memory[23157] <=  8'h00;      memory[23158] <=  8'h00;      memory[23159] <=  8'h00;      memory[23160] <=  8'h00;      memory[23161] <=  8'h00;      memory[23162] <=  8'h00;      memory[23163] <=  8'h00;      memory[23164] <=  8'h00;      memory[23165] <=  8'h00;      memory[23166] <=  8'h00;      memory[23167] <=  8'h00;      memory[23168] <=  8'h00;      memory[23169] <=  8'h00;      memory[23170] <=  8'h00;      memory[23171] <=  8'h00;      memory[23172] <=  8'h00;      memory[23173] <=  8'h00;      memory[23174] <=  8'h00;      memory[23175] <=  8'h00;      memory[23176] <=  8'h00;      memory[23177] <=  8'h00;      memory[23178] <=  8'h00;      memory[23179] <=  8'h00;      memory[23180] <=  8'h00;      memory[23181] <=  8'h00;      memory[23182] <=  8'h00;      memory[23183] <=  8'h00;      memory[23184] <=  8'h00;      memory[23185] <=  8'h00;      memory[23186] <=  8'h00;      memory[23187] <=  8'h00;      memory[23188] <=  8'h00;      memory[23189] <=  8'h00;      memory[23190] <=  8'h00;      memory[23191] <=  8'h00;      memory[23192] <=  8'h00;      memory[23193] <=  8'h00;      memory[23194] <=  8'h00;      memory[23195] <=  8'h00;      memory[23196] <=  8'h00;      memory[23197] <=  8'h00;      memory[23198] <=  8'h00;      memory[23199] <=  8'h00;      memory[23200] <=  8'h00;      memory[23201] <=  8'h00;      memory[23202] <=  8'h00;      memory[23203] <=  8'h00;      memory[23204] <=  8'h00;      memory[23205] <=  8'h00;      memory[23206] <=  8'h00;      memory[23207] <=  8'h00;      memory[23208] <=  8'h00;      memory[23209] <=  8'h00;      memory[23210] <=  8'h00;      memory[23211] <=  8'h00;      memory[23212] <=  8'h00;      memory[23213] <=  8'h00;      memory[23214] <=  8'h00;      memory[23215] <=  8'h00;      memory[23216] <=  8'h00;      memory[23217] <=  8'h00;      memory[23218] <=  8'h00;      memory[23219] <=  8'h00;      memory[23220] <=  8'h00;      memory[23221] <=  8'h00;      memory[23222] <=  8'h00;      memory[23223] <=  8'h00;      memory[23224] <=  8'h00;      memory[23225] <=  8'h00;      memory[23226] <=  8'h00;      memory[23227] <=  8'h00;      memory[23228] <=  8'h00;      memory[23229] <=  8'h00;      memory[23230] <=  8'h00;      memory[23231] <=  8'h00;      memory[23232] <=  8'h00;      memory[23233] <=  8'h00;      memory[23234] <=  8'h00;      memory[23235] <=  8'h00;      memory[23236] <=  8'h00;      memory[23237] <=  8'h00;      memory[23238] <=  8'h00;      memory[23239] <=  8'h00;      memory[23240] <=  8'h00;      memory[23241] <=  8'h00;      memory[23242] <=  8'h00;      memory[23243] <=  8'h00;      memory[23244] <=  8'h00;      memory[23245] <=  8'h00;      memory[23246] <=  8'h00;      memory[23247] <=  8'h00;      memory[23248] <=  8'h00;      memory[23249] <=  8'h00;      memory[23250] <=  8'h00;      memory[23251] <=  8'h00;      memory[23252] <=  8'h00;      memory[23253] <=  8'h00;      memory[23254] <=  8'h00;      memory[23255] <=  8'h00;      memory[23256] <=  8'h00;      memory[23257] <=  8'h00;      memory[23258] <=  8'h00;      memory[23259] <=  8'h00;      memory[23260] <=  8'h00;      memory[23261] <=  8'h00;      memory[23262] <=  8'h00;      memory[23263] <=  8'h00;      memory[23264] <=  8'h00;      memory[23265] <=  8'h00;      memory[23266] <=  8'h00;      memory[23267] <=  8'h00;      memory[23268] <=  8'h00;      memory[23269] <=  8'h00;      memory[23270] <=  8'h00;      memory[23271] <=  8'h00;      memory[23272] <=  8'h00;      memory[23273] <=  8'h00;      memory[23274] <=  8'h00;      memory[23275] <=  8'h00;      memory[23276] <=  8'h00;      memory[23277] <=  8'h00;      memory[23278] <=  8'h00;      memory[23279] <=  8'h00;      memory[23280] <=  8'h00;      memory[23281] <=  8'h00;      memory[23282] <=  8'h00;      memory[23283] <=  8'h00;      memory[23284] <=  8'h00;      memory[23285] <=  8'h00;      memory[23286] <=  8'h00;      memory[23287] <=  8'h00;      memory[23288] <=  8'h00;      memory[23289] <=  8'h00;      memory[23290] <=  8'h00;      memory[23291] <=  8'h00;      memory[23292] <=  8'h00;      memory[23293] <=  8'h00;      memory[23294] <=  8'h00;      memory[23295] <=  8'h00;      memory[23296] <=  8'h00;      memory[23297] <=  8'h00;      memory[23298] <=  8'h00;      memory[23299] <=  8'h00;      memory[23300] <=  8'h00;      memory[23301] <=  8'h00;      memory[23302] <=  8'h00;      memory[23303] <=  8'h00;      memory[23304] <=  8'h00;      memory[23305] <=  8'h00;      memory[23306] <=  8'h00;      memory[23307] <=  8'h00;      memory[23308] <=  8'h00;      memory[23309] <=  8'h00;      memory[23310] <=  8'h00;      memory[23311] <=  8'h00;      memory[23312] <=  8'h00;      memory[23313] <=  8'h00;      memory[23314] <=  8'h00;      memory[23315] <=  8'h00;      memory[23316] <=  8'h00;      memory[23317] <=  8'h00;      memory[23318] <=  8'h00;      memory[23319] <=  8'h00;      memory[23320] <=  8'h00;      memory[23321] <=  8'h00;      memory[23322] <=  8'h00;      memory[23323] <=  8'h00;      memory[23324] <=  8'h00;      memory[23325] <=  8'h00;      memory[23326] <=  8'h00;      memory[23327] <=  8'h00;      memory[23328] <=  8'h00;      memory[23329] <=  8'h00;      memory[23330] <=  8'h00;      memory[23331] <=  8'h00;      memory[23332] <=  8'h00;      memory[23333] <=  8'h00;      memory[23334] <=  8'h00;      memory[23335] <=  8'h00;      memory[23336] <=  8'h00;      memory[23337] <=  8'h00;      memory[23338] <=  8'h00;      memory[23339] <=  8'h00;      memory[23340] <=  8'h00;      memory[23341] <=  8'h00;      memory[23342] <=  8'h00;      memory[23343] <=  8'h00;      memory[23344] <=  8'h00;      memory[23345] <=  8'h00;      memory[23346] <=  8'h00;      memory[23347] <=  8'h00;      memory[23348] <=  8'h00;      memory[23349] <=  8'h00;      memory[23350] <=  8'h00;      memory[23351] <=  8'h00;      memory[23352] <=  8'h00;      memory[23353] <=  8'h00;      memory[23354] <=  8'h00;      memory[23355] <=  8'h00;      memory[23356] <=  8'h00;      memory[23357] <=  8'h00;      memory[23358] <=  8'h00;      memory[23359] <=  8'h00;      memory[23360] <=  8'h00;      memory[23361] <=  8'h00;      memory[23362] <=  8'h00;      memory[23363] <=  8'h00;      memory[23364] <=  8'h00;      memory[23365] <=  8'h00;      memory[23366] <=  8'h00;      memory[23367] <=  8'h00;      memory[23368] <=  8'h00;      memory[23369] <=  8'h00;      memory[23370] <=  8'h00;      memory[23371] <=  8'h00;      memory[23372] <=  8'h00;      memory[23373] <=  8'h00;      memory[23374] <=  8'h00;      memory[23375] <=  8'h00;      memory[23376] <=  8'h00;      memory[23377] <=  8'h00;      memory[23378] <=  8'h00;      memory[23379] <=  8'h00;      memory[23380] <=  8'h00;      memory[23381] <=  8'h00;      memory[23382] <=  8'h00;      memory[23383] <=  8'h00;      memory[23384] <=  8'h00;      memory[23385] <=  8'h00;      memory[23386] <=  8'h00;      memory[23387] <=  8'h00;      memory[23388] <=  8'h00;      memory[23389] <=  8'h00;      memory[23390] <=  8'h00;      memory[23391] <=  8'h00;      memory[23392] <=  8'h00;      memory[23393] <=  8'h00;      memory[23394] <=  8'h00;      memory[23395] <=  8'h00;      memory[23396] <=  8'h00;      memory[23397] <=  8'h00;      memory[23398] <=  8'h00;      memory[23399] <=  8'h00;      memory[23400] <=  8'h00;      memory[23401] <=  8'h00;      memory[23402] <=  8'h00;      memory[23403] <=  8'h00;      memory[23404] <=  8'h00;      memory[23405] <=  8'h00;      memory[23406] <=  8'h00;      memory[23407] <=  8'h00;      memory[23408] <=  8'h00;      memory[23409] <=  8'h00;      memory[23410] <=  8'h00;      memory[23411] <=  8'h00;      memory[23412] <=  8'h00;      memory[23413] <=  8'h00;      memory[23414] <=  8'h00;      memory[23415] <=  8'h00;      memory[23416] <=  8'h00;      memory[23417] <=  8'h00;      memory[23418] <=  8'h00;      memory[23419] <=  8'h00;      memory[23420] <=  8'h00;      memory[23421] <=  8'h00;      memory[23422] <=  8'h00;      memory[23423] <=  8'h00;      memory[23424] <=  8'h00;      memory[23425] <=  8'h00;      memory[23426] <=  8'h00;      memory[23427] <=  8'h00;      memory[23428] <=  8'h00;      memory[23429] <=  8'h00;      memory[23430] <=  8'h00;      memory[23431] <=  8'h00;      memory[23432] <=  8'h00;      memory[23433] <=  8'h00;      memory[23434] <=  8'h00;      memory[23435] <=  8'h00;      memory[23436] <=  8'h00;      memory[23437] <=  8'h00;      memory[23438] <=  8'h00;      memory[23439] <=  8'h00;      memory[23440] <=  8'h00;      memory[23441] <=  8'h00;      memory[23442] <=  8'h00;      memory[23443] <=  8'h00;      memory[23444] <=  8'h00;      memory[23445] <=  8'h00;      memory[23446] <=  8'h00;      memory[23447] <=  8'h00;      memory[23448] <=  8'h00;      memory[23449] <=  8'h00;      memory[23450] <=  8'h00;      memory[23451] <=  8'h00;      memory[23452] <=  8'h00;      memory[23453] <=  8'h00;      memory[23454] <=  8'h00;      memory[23455] <=  8'h00;      memory[23456] <=  8'h00;      memory[23457] <=  8'h00;      memory[23458] <=  8'h00;      memory[23459] <=  8'h00;      memory[23460] <=  8'h00;      memory[23461] <=  8'h00;      memory[23462] <=  8'h00;      memory[23463] <=  8'h00;      memory[23464] <=  8'h00;      memory[23465] <=  8'h00;      memory[23466] <=  8'h00;      memory[23467] <=  8'h00;      memory[23468] <=  8'h00;      memory[23469] <=  8'h00;      memory[23470] <=  8'h00;      memory[23471] <=  8'h00;      memory[23472] <=  8'h00;      memory[23473] <=  8'h00;      memory[23474] <=  8'h00;      memory[23475] <=  8'h00;      memory[23476] <=  8'h00;      memory[23477] <=  8'h00;      memory[23478] <=  8'h00;      memory[23479] <=  8'h00;      memory[23480] <=  8'h00;      memory[23481] <=  8'h00;      memory[23482] <=  8'h00;      memory[23483] <=  8'h00;      memory[23484] <=  8'h00;      memory[23485] <=  8'h00;      memory[23486] <=  8'h00;      memory[23487] <=  8'h00;      memory[23488] <=  8'h00;      memory[23489] <=  8'h00;      memory[23490] <=  8'h00;      memory[23491] <=  8'h00;      memory[23492] <=  8'h00;      memory[23493] <=  8'h00;      memory[23494] <=  8'h00;      memory[23495] <=  8'h00;      memory[23496] <=  8'h00;      memory[23497] <=  8'h00;      memory[23498] <=  8'h00;      memory[23499] <=  8'h00;      memory[23500] <=  8'h00;      memory[23501] <=  8'h00;      memory[23502] <=  8'h00;      memory[23503] <=  8'h00;      memory[23504] <=  8'h00;      memory[23505] <=  8'h00;      memory[23506] <=  8'h00;      memory[23507] <=  8'h00;      memory[23508] <=  8'h00;      memory[23509] <=  8'h00;      memory[23510] <=  8'h00;      memory[23511] <=  8'h00;      memory[23512] <=  8'h00;      memory[23513] <=  8'h00;      memory[23514] <=  8'h00;      memory[23515] <=  8'h00;      memory[23516] <=  8'h00;      memory[23517] <=  8'h00;      memory[23518] <=  8'h00;      memory[23519] <=  8'h00;      memory[23520] <=  8'h00;      memory[23521] <=  8'h00;      memory[23522] <=  8'h00;      memory[23523] <=  8'h00;      memory[23524] <=  8'h00;      memory[23525] <=  8'h00;      memory[23526] <=  8'h00;      memory[23527] <=  8'h00;      memory[23528] <=  8'h00;      memory[23529] <=  8'h00;      memory[23530] <=  8'h00;      memory[23531] <=  8'h00;      memory[23532] <=  8'h00;      memory[23533] <=  8'h00;      memory[23534] <=  8'h00;      memory[23535] <=  8'h00;      memory[23536] <=  8'h00;      memory[23537] <=  8'h00;      memory[23538] <=  8'h00;      memory[23539] <=  8'h00;      memory[23540] <=  8'h00;      memory[23541] <=  8'h00;      memory[23542] <=  8'h00;      memory[23543] <=  8'h00;      memory[23544] <=  8'h00;      memory[23545] <=  8'h00;      memory[23546] <=  8'h00;      memory[23547] <=  8'h00;      memory[23548] <=  8'h00;      memory[23549] <=  8'h00;      memory[23550] <=  8'h00;      memory[23551] <=  8'h00;      memory[23552] <=  8'h00;      memory[23553] <=  8'h00;      memory[23554] <=  8'h00;      memory[23555] <=  8'h00;      memory[23556] <=  8'h00;      memory[23557] <=  8'h00;      memory[23558] <=  8'h00;      memory[23559] <=  8'h00;      memory[23560] <=  8'h00;      memory[23561] <=  8'h00;      memory[23562] <=  8'h00;      memory[23563] <=  8'h00;      memory[23564] <=  8'h00;      memory[23565] <=  8'h00;      memory[23566] <=  8'h00;      memory[23567] <=  8'h00;      memory[23568] <=  8'h00;      memory[23569] <=  8'h00;      memory[23570] <=  8'h00;      memory[23571] <=  8'h00;      memory[23572] <=  8'h00;      memory[23573] <=  8'h00;      memory[23574] <=  8'h00;      memory[23575] <=  8'h00;      memory[23576] <=  8'h00;      memory[23577] <=  8'h00;      memory[23578] <=  8'h00;      memory[23579] <=  8'h00;      memory[23580] <=  8'h00;      memory[23581] <=  8'h00;      memory[23582] <=  8'h00;      memory[23583] <=  8'h00;      memory[23584] <=  8'h00;      memory[23585] <=  8'h00;      memory[23586] <=  8'h00;      memory[23587] <=  8'h00;      memory[23588] <=  8'h00;      memory[23589] <=  8'h00;      memory[23590] <=  8'h00;      memory[23591] <=  8'h00;      memory[23592] <=  8'h00;      memory[23593] <=  8'h00;      memory[23594] <=  8'h00;      memory[23595] <=  8'h00;      memory[23596] <=  8'h00;      memory[23597] <=  8'h00;      memory[23598] <=  8'h00;      memory[23599] <=  8'h00;      memory[23600] <=  8'h00;      memory[23601] <=  8'h00;      memory[23602] <=  8'h00;      memory[23603] <=  8'h00;      memory[23604] <=  8'h00;      memory[23605] <=  8'h00;      memory[23606] <=  8'h00;      memory[23607] <=  8'h00;      memory[23608] <=  8'h00;      memory[23609] <=  8'h00;      memory[23610] <=  8'h00;      memory[23611] <=  8'h00;      memory[23612] <=  8'h00;      memory[23613] <=  8'h00;      memory[23614] <=  8'h00;      memory[23615] <=  8'h00;      memory[23616] <=  8'h00;      memory[23617] <=  8'h00;      memory[23618] <=  8'h00;      memory[23619] <=  8'h00;      memory[23620] <=  8'h00;      memory[23621] <=  8'h00;      memory[23622] <=  8'h00;      memory[23623] <=  8'h00;      memory[23624] <=  8'h00;      memory[23625] <=  8'h00;      memory[23626] <=  8'h00;      memory[23627] <=  8'h00;      memory[23628] <=  8'h00;      memory[23629] <=  8'h00;      memory[23630] <=  8'h00;      memory[23631] <=  8'h00;      memory[23632] <=  8'h00;      memory[23633] <=  8'h00;      memory[23634] <=  8'h00;      memory[23635] <=  8'h00;      memory[23636] <=  8'h00;      memory[23637] <=  8'h00;      memory[23638] <=  8'h00;      memory[23639] <=  8'h00;      memory[23640] <=  8'h00;      memory[23641] <=  8'h00;      memory[23642] <=  8'h00;      memory[23643] <=  8'h00;      memory[23644] <=  8'h00;      memory[23645] <=  8'h00;      memory[23646] <=  8'h00;      memory[23647] <=  8'h00;      memory[23648] <=  8'h00;      memory[23649] <=  8'h00;      memory[23650] <=  8'h00;      memory[23651] <=  8'h00;      memory[23652] <=  8'h00;      memory[23653] <=  8'h00;      memory[23654] <=  8'h00;      memory[23655] <=  8'h00;      memory[23656] <=  8'h00;      memory[23657] <=  8'h00;      memory[23658] <=  8'h00;      memory[23659] <=  8'h00;      memory[23660] <=  8'h00;      memory[23661] <=  8'h00;      memory[23662] <=  8'h00;      memory[23663] <=  8'h00;      memory[23664] <=  8'h00;      memory[23665] <=  8'h00;      memory[23666] <=  8'h00;      memory[23667] <=  8'h00;      memory[23668] <=  8'h00;      memory[23669] <=  8'h00;      memory[23670] <=  8'h00;      memory[23671] <=  8'h00;      memory[23672] <=  8'h00;      memory[23673] <=  8'h00;      memory[23674] <=  8'h00;      memory[23675] <=  8'h00;      memory[23676] <=  8'h00;      memory[23677] <=  8'h00;      memory[23678] <=  8'h00;      memory[23679] <=  8'h00;      memory[23680] <=  8'h00;      memory[23681] <=  8'h00;      memory[23682] <=  8'h00;      memory[23683] <=  8'h00;      memory[23684] <=  8'h00;      memory[23685] <=  8'h00;      memory[23686] <=  8'h00;      memory[23687] <=  8'h00;      memory[23688] <=  8'h00;      memory[23689] <=  8'h00;      memory[23690] <=  8'h00;      memory[23691] <=  8'h00;      memory[23692] <=  8'h00;      memory[23693] <=  8'h00;      memory[23694] <=  8'h00;      memory[23695] <=  8'h00;      memory[23696] <=  8'h00;      memory[23697] <=  8'h00;      memory[23698] <=  8'h00;      memory[23699] <=  8'h00;      memory[23700] <=  8'h00;      memory[23701] <=  8'h00;      memory[23702] <=  8'h00;      memory[23703] <=  8'h00;      memory[23704] <=  8'h00;      memory[23705] <=  8'h00;      memory[23706] <=  8'h00;      memory[23707] <=  8'h00;      memory[23708] <=  8'h00;      memory[23709] <=  8'h00;      memory[23710] <=  8'h00;      memory[23711] <=  8'h00;      memory[23712] <=  8'h00;      memory[23713] <=  8'h00;      memory[23714] <=  8'h00;      memory[23715] <=  8'h00;      memory[23716] <=  8'h00;      memory[23717] <=  8'h00;      memory[23718] <=  8'h00;      memory[23719] <=  8'h00;      memory[23720] <=  8'h00;      memory[23721] <=  8'h00;      memory[23722] <=  8'h00;      memory[23723] <=  8'h00;      memory[23724] <=  8'h00;      memory[23725] <=  8'h00;      memory[23726] <=  8'h00;      memory[23727] <=  8'h00;      memory[23728] <=  8'h00;      memory[23729] <=  8'h00;      memory[23730] <=  8'h00;      memory[23731] <=  8'h00;      memory[23732] <=  8'h00;      memory[23733] <=  8'h00;      memory[23734] <=  8'h00;      memory[23735] <=  8'h00;      memory[23736] <=  8'h00;      memory[23737] <=  8'h00;      memory[23738] <=  8'h00;      memory[23739] <=  8'h00;      memory[23740] <=  8'h00;      memory[23741] <=  8'h00;      memory[23742] <=  8'h00;      memory[23743] <=  8'h00;      memory[23744] <=  8'h00;      memory[23745] <=  8'h00;      memory[23746] <=  8'h00;      memory[23747] <=  8'h00;      memory[23748] <=  8'h00;      memory[23749] <=  8'h00;      memory[23750] <=  8'h00;      memory[23751] <=  8'h00;      memory[23752] <=  8'h00;      memory[23753] <=  8'h00;      memory[23754] <=  8'h00;      memory[23755] <=  8'h00;      memory[23756] <=  8'h00;      memory[23757] <=  8'h00;      memory[23758] <=  8'h00;      memory[23759] <=  8'h00;      memory[23760] <=  8'h00;      memory[23761] <=  8'h00;      memory[23762] <=  8'h00;      memory[23763] <=  8'h00;      memory[23764] <=  8'h00;      memory[23765] <=  8'h00;      memory[23766] <=  8'h00;      memory[23767] <=  8'h00;      memory[23768] <=  8'h00;      memory[23769] <=  8'h00;      memory[23770] <=  8'h00;      memory[23771] <=  8'h00;      memory[23772] <=  8'h00;      memory[23773] <=  8'h00;      memory[23774] <=  8'h00;      memory[23775] <=  8'h00;      memory[23776] <=  8'h00;      memory[23777] <=  8'h00;      memory[23778] <=  8'h00;      memory[23779] <=  8'h00;      memory[23780] <=  8'h00;      memory[23781] <=  8'h00;      memory[23782] <=  8'h00;      memory[23783] <=  8'h00;      memory[23784] <=  8'h00;      memory[23785] <=  8'h00;      memory[23786] <=  8'h00;      memory[23787] <=  8'h00;      memory[23788] <=  8'h00;      memory[23789] <=  8'h00;      memory[23790] <=  8'h00;      memory[23791] <=  8'h00;      memory[23792] <=  8'h00;      memory[23793] <=  8'h00;      memory[23794] <=  8'h00;      memory[23795] <=  8'h00;      memory[23796] <=  8'h00;      memory[23797] <=  8'h00;      memory[23798] <=  8'h00;      memory[23799] <=  8'h00;      memory[23800] <=  8'h00;      memory[23801] <=  8'h00;      memory[23802] <=  8'h00;      memory[23803] <=  8'h00;      memory[23804] <=  8'h00;      memory[23805] <=  8'h00;      memory[23806] <=  8'h00;      memory[23807] <=  8'h00;      memory[23808] <=  8'h00;      memory[23809] <=  8'h00;      memory[23810] <=  8'h00;      memory[23811] <=  8'h00;      memory[23812] <=  8'h00;      memory[23813] <=  8'h00;      memory[23814] <=  8'h00;      memory[23815] <=  8'h00;      memory[23816] <=  8'h00;      memory[23817] <=  8'h00;      memory[23818] <=  8'h00;      memory[23819] <=  8'h00;      memory[23820] <=  8'h00;      memory[23821] <=  8'h00;      memory[23822] <=  8'h00;      memory[23823] <=  8'h00;      memory[23824] <=  8'h00;      memory[23825] <=  8'h00;      memory[23826] <=  8'h00;      memory[23827] <=  8'h00;      memory[23828] <=  8'h00;      memory[23829] <=  8'h00;      memory[23830] <=  8'h00;      memory[23831] <=  8'h00;      memory[23832] <=  8'h00;      memory[23833] <=  8'h00;      memory[23834] <=  8'h00;      memory[23835] <=  8'h00;      memory[23836] <=  8'h00;      memory[23837] <=  8'h00;      memory[23838] <=  8'h00;      memory[23839] <=  8'h00;      memory[23840] <=  8'h00;      memory[23841] <=  8'h00;      memory[23842] <=  8'h00;      memory[23843] <=  8'h00;      memory[23844] <=  8'h00;      memory[23845] <=  8'h00;      memory[23846] <=  8'h00;      memory[23847] <=  8'h00;      memory[23848] <=  8'h00;      memory[23849] <=  8'h00;      memory[23850] <=  8'h00;      memory[23851] <=  8'h00;      memory[23852] <=  8'h00;      memory[23853] <=  8'h00;      memory[23854] <=  8'h00;      memory[23855] <=  8'h00;      memory[23856] <=  8'h00;      memory[23857] <=  8'h00;      memory[23858] <=  8'h00;      memory[23859] <=  8'h00;      memory[23860] <=  8'h00;      memory[23861] <=  8'h00;      memory[23862] <=  8'h00;      memory[23863] <=  8'h00;      memory[23864] <=  8'h00;      memory[23865] <=  8'h00;      memory[23866] <=  8'h00;      memory[23867] <=  8'h00;      memory[23868] <=  8'h00;      memory[23869] <=  8'h00;      memory[23870] <=  8'h00;      memory[23871] <=  8'h00;      memory[23872] <=  8'h00;      memory[23873] <=  8'h00;      memory[23874] <=  8'h00;      memory[23875] <=  8'h00;      memory[23876] <=  8'h00;      memory[23877] <=  8'h00;      memory[23878] <=  8'h00;      memory[23879] <=  8'h00;      memory[23880] <=  8'h00;      memory[23881] <=  8'h00;      memory[23882] <=  8'h00;      memory[23883] <=  8'h00;      memory[23884] <=  8'h00;      memory[23885] <=  8'h00;      memory[23886] <=  8'h00;      memory[23887] <=  8'h00;      memory[23888] <=  8'h00;      memory[23889] <=  8'h00;      memory[23890] <=  8'h00;      memory[23891] <=  8'h00;      memory[23892] <=  8'h00;      memory[23893] <=  8'h00;      memory[23894] <=  8'h00;      memory[23895] <=  8'h00;      memory[23896] <=  8'h00;      memory[23897] <=  8'h00;      memory[23898] <=  8'h00;      memory[23899] <=  8'h00;      memory[23900] <=  8'h00;      memory[23901] <=  8'h00;      memory[23902] <=  8'h00;      memory[23903] <=  8'h00;      memory[23904] <=  8'h00;      memory[23905] <=  8'h00;      memory[23906] <=  8'h00;      memory[23907] <=  8'h00;      memory[23908] <=  8'h00;      memory[23909] <=  8'h00;      memory[23910] <=  8'h00;      memory[23911] <=  8'h00;      memory[23912] <=  8'h00;      memory[23913] <=  8'h00;      memory[23914] <=  8'h00;      memory[23915] <=  8'h00;      memory[23916] <=  8'h00;      memory[23917] <=  8'h00;      memory[23918] <=  8'h00;      memory[23919] <=  8'h00;      memory[23920] <=  8'h00;      memory[23921] <=  8'h00;      memory[23922] <=  8'h00;      memory[23923] <=  8'h00;      memory[23924] <=  8'h00;      memory[23925] <=  8'h00;      memory[23926] <=  8'h00;      memory[23927] <=  8'h00;      memory[23928] <=  8'h00;      memory[23929] <=  8'h00;      memory[23930] <=  8'h00;      memory[23931] <=  8'h00;      memory[23932] <=  8'h00;      memory[23933] <=  8'h00;      memory[23934] <=  8'h00;      memory[23935] <=  8'h00;      memory[23936] <=  8'h00;      memory[23937] <=  8'h00;      memory[23938] <=  8'h00;      memory[23939] <=  8'h00;      memory[23940] <=  8'h00;      memory[23941] <=  8'h00;      memory[23942] <=  8'h00;      memory[23943] <=  8'h00;      memory[23944] <=  8'h00;      memory[23945] <=  8'h00;      memory[23946] <=  8'h00;      memory[23947] <=  8'h00;      memory[23948] <=  8'h00;      memory[23949] <=  8'h00;      memory[23950] <=  8'h00;      memory[23951] <=  8'h00;      memory[23952] <=  8'h00;      memory[23953] <=  8'h00;      memory[23954] <=  8'h00;      memory[23955] <=  8'h00;      memory[23956] <=  8'h00;      memory[23957] <=  8'h00;      memory[23958] <=  8'h00;      memory[23959] <=  8'h00;      memory[23960] <=  8'h00;      memory[23961] <=  8'h00;      memory[23962] <=  8'h00;      memory[23963] <=  8'h00;      memory[23964] <=  8'h00;      memory[23965] <=  8'h00;      memory[23966] <=  8'h00;      memory[23967] <=  8'h00;      memory[23968] <=  8'h00;      memory[23969] <=  8'h00;      memory[23970] <=  8'h00;      memory[23971] <=  8'h00;      memory[23972] <=  8'h00;      memory[23973] <=  8'h00;      memory[23974] <=  8'h00;      memory[23975] <=  8'h00;      memory[23976] <=  8'h00;      memory[23977] <=  8'h00;      memory[23978] <=  8'h00;      memory[23979] <=  8'h00;      memory[23980] <=  8'h00;      memory[23981] <=  8'h00;      memory[23982] <=  8'h00;      memory[23983] <=  8'h00;      memory[23984] <=  8'h00;      memory[23985] <=  8'h00;      memory[23986] <=  8'h00;      memory[23987] <=  8'h00;      memory[23988] <=  8'h00;      memory[23989] <=  8'h00;      memory[23990] <=  8'h00;      memory[23991] <=  8'h00;      memory[23992] <=  8'h00;      memory[23993] <=  8'h00;      memory[23994] <=  8'h00;      memory[23995] <=  8'h00;      memory[23996] <=  8'h00;      memory[23997] <=  8'h00;      memory[23998] <=  8'h00;      memory[23999] <=  8'h00;      memory[24000] <=  8'h00;      memory[24001] <=  8'h00;      memory[24002] <=  8'h00;      memory[24003] <=  8'h00;      memory[24004] <=  8'h00;      memory[24005] <=  8'h00;      memory[24006] <=  8'h00;      memory[24007] <=  8'h00;      memory[24008] <=  8'h00;      memory[24009] <=  8'h00;      memory[24010] <=  8'h00;      memory[24011] <=  8'h00;      memory[24012] <=  8'h00;      memory[24013] <=  8'h00;      memory[24014] <=  8'h00;      memory[24015] <=  8'h00;      memory[24016] <=  8'h00;      memory[24017] <=  8'h00;      memory[24018] <=  8'h00;      memory[24019] <=  8'h00;      memory[24020] <=  8'h00;      memory[24021] <=  8'h00;      memory[24022] <=  8'h00;      memory[24023] <=  8'h00;      memory[24024] <=  8'h00;      memory[24025] <=  8'h00;      memory[24026] <=  8'h00;      memory[24027] <=  8'h00;      memory[24028] <=  8'h00;      memory[24029] <=  8'h00;      memory[24030] <=  8'h00;      memory[24031] <=  8'h00;      memory[24032] <=  8'h00;      memory[24033] <=  8'h00;      memory[24034] <=  8'h00;      memory[24035] <=  8'h00;      memory[24036] <=  8'h00;      memory[24037] <=  8'h00;      memory[24038] <=  8'h00;      memory[24039] <=  8'h00;      memory[24040] <=  8'h00;      memory[24041] <=  8'h00;      memory[24042] <=  8'h00;      memory[24043] <=  8'h00;      memory[24044] <=  8'h00;      memory[24045] <=  8'h00;      memory[24046] <=  8'h00;      memory[24047] <=  8'h00;      memory[24048] <=  8'h00;      memory[24049] <=  8'h00;      memory[24050] <=  8'h00;      memory[24051] <=  8'h00;      memory[24052] <=  8'h00;      memory[24053] <=  8'h00;      memory[24054] <=  8'h00;      memory[24055] <=  8'h00;      memory[24056] <=  8'h00;      memory[24057] <=  8'h00;      memory[24058] <=  8'h00;      memory[24059] <=  8'h00;      memory[24060] <=  8'h00;      memory[24061] <=  8'h00;      memory[24062] <=  8'h00;      memory[24063] <=  8'h00;      memory[24064] <=  8'h00;      memory[24065] <=  8'h00;      memory[24066] <=  8'h00;      memory[24067] <=  8'h00;      memory[24068] <=  8'h00;      memory[24069] <=  8'h00;      memory[24070] <=  8'h00;      memory[24071] <=  8'h00;      memory[24072] <=  8'h00;      memory[24073] <=  8'h00;      memory[24074] <=  8'h00;      memory[24075] <=  8'h00;      memory[24076] <=  8'h00;      memory[24077] <=  8'h00;      memory[24078] <=  8'h00;      memory[24079] <=  8'h00;      memory[24080] <=  8'h00;      memory[24081] <=  8'h00;      memory[24082] <=  8'h00;      memory[24083] <=  8'h00;      memory[24084] <=  8'h00;      memory[24085] <=  8'h00;      memory[24086] <=  8'h00;      memory[24087] <=  8'h00;      memory[24088] <=  8'h00;      memory[24089] <=  8'h00;      memory[24090] <=  8'h00;      memory[24091] <=  8'h00;      memory[24092] <=  8'h00;      memory[24093] <=  8'h00;      memory[24094] <=  8'h00;      memory[24095] <=  8'h00;      memory[24096] <=  8'h00;      memory[24097] <=  8'h00;      memory[24098] <=  8'h00;      memory[24099] <=  8'h00;      memory[24100] <=  8'h00;      memory[24101] <=  8'h00;      memory[24102] <=  8'h00;      memory[24103] <=  8'h00;      memory[24104] <=  8'h00;      memory[24105] <=  8'h00;      memory[24106] <=  8'h00;      memory[24107] <=  8'h00;      memory[24108] <=  8'h00;      memory[24109] <=  8'h00;      memory[24110] <=  8'h00;      memory[24111] <=  8'h00;      memory[24112] <=  8'h00;      memory[24113] <=  8'h00;      memory[24114] <=  8'h00;      memory[24115] <=  8'h00;      memory[24116] <=  8'h00;      memory[24117] <=  8'h00;      memory[24118] <=  8'h00;      memory[24119] <=  8'h00;      memory[24120] <=  8'h00;      memory[24121] <=  8'h00;      memory[24122] <=  8'h00;      memory[24123] <=  8'h00;      memory[24124] <=  8'h00;      memory[24125] <=  8'h00;      memory[24126] <=  8'h00;      memory[24127] <=  8'h00;      memory[24128] <=  8'h00;      memory[24129] <=  8'h00;      memory[24130] <=  8'h00;      memory[24131] <=  8'h00;      memory[24132] <=  8'h00;      memory[24133] <=  8'h00;      memory[24134] <=  8'h00;      memory[24135] <=  8'h00;      memory[24136] <=  8'h00;      memory[24137] <=  8'h00;      memory[24138] <=  8'h00;      memory[24139] <=  8'h00;      memory[24140] <=  8'h00;      memory[24141] <=  8'h00;      memory[24142] <=  8'h00;      memory[24143] <=  8'h00;      memory[24144] <=  8'h00;      memory[24145] <=  8'h00;      memory[24146] <=  8'h00;      memory[24147] <=  8'h00;      memory[24148] <=  8'h00;      memory[24149] <=  8'h00;      memory[24150] <=  8'h00;      memory[24151] <=  8'h00;      memory[24152] <=  8'h00;      memory[24153] <=  8'h00;      memory[24154] <=  8'h00;      memory[24155] <=  8'h00;      memory[24156] <=  8'h00;      memory[24157] <=  8'h00;      memory[24158] <=  8'h00;      memory[24159] <=  8'h00;      memory[24160] <=  8'h00;      memory[24161] <=  8'h00;      memory[24162] <=  8'h00;      memory[24163] <=  8'h00;      memory[24164] <=  8'h00;      memory[24165] <=  8'h00;      memory[24166] <=  8'h00;      memory[24167] <=  8'h00;      memory[24168] <=  8'h00;      memory[24169] <=  8'h00;      memory[24170] <=  8'h00;      memory[24171] <=  8'h00;      memory[24172] <=  8'h00;      memory[24173] <=  8'h00;      memory[24174] <=  8'h00;      memory[24175] <=  8'h00;      memory[24176] <=  8'h00;      memory[24177] <=  8'h00;      memory[24178] <=  8'h00;      memory[24179] <=  8'h00;      memory[24180] <=  8'h00;      memory[24181] <=  8'h00;      memory[24182] <=  8'h00;      memory[24183] <=  8'h00;      memory[24184] <=  8'h00;      memory[24185] <=  8'h00;      memory[24186] <=  8'h00;      memory[24187] <=  8'h00;      memory[24188] <=  8'h00;      memory[24189] <=  8'h00;      memory[24190] <=  8'h00;      memory[24191] <=  8'h00;      memory[24192] <=  8'h00;      memory[24193] <=  8'h00;      memory[24194] <=  8'h00;      memory[24195] <=  8'h00;      memory[24196] <=  8'h00;      memory[24197] <=  8'h00;      memory[24198] <=  8'h00;      memory[24199] <=  8'h00;      memory[24200] <=  8'h00;      memory[24201] <=  8'h00;      memory[24202] <=  8'h00;      memory[24203] <=  8'h00;      memory[24204] <=  8'h00;      memory[24205] <=  8'h00;      memory[24206] <=  8'h00;      memory[24207] <=  8'h00;      memory[24208] <=  8'h00;      memory[24209] <=  8'h00;      memory[24210] <=  8'h00;      memory[24211] <=  8'h00;      memory[24212] <=  8'h00;      memory[24213] <=  8'h00;      memory[24214] <=  8'h00;      memory[24215] <=  8'h00;      memory[24216] <=  8'h00;      memory[24217] <=  8'h00;      memory[24218] <=  8'h00;      memory[24219] <=  8'h00;      memory[24220] <=  8'h00;      memory[24221] <=  8'h00;      memory[24222] <=  8'h00;      memory[24223] <=  8'h00;      memory[24224] <=  8'h00;      memory[24225] <=  8'h00;      memory[24226] <=  8'h00;      memory[24227] <=  8'h00;      memory[24228] <=  8'h00;      memory[24229] <=  8'h00;      memory[24230] <=  8'h00;      memory[24231] <=  8'h00;      memory[24232] <=  8'h00;      memory[24233] <=  8'h00;      memory[24234] <=  8'h00;      memory[24235] <=  8'h00;      memory[24236] <=  8'h00;      memory[24237] <=  8'h00;      memory[24238] <=  8'h00;      memory[24239] <=  8'h00;      memory[24240] <=  8'h00;      memory[24241] <=  8'h00;      memory[24242] <=  8'h00;      memory[24243] <=  8'h00;      memory[24244] <=  8'h00;      memory[24245] <=  8'h00;      memory[24246] <=  8'h00;      memory[24247] <=  8'h00;      memory[24248] <=  8'h00;      memory[24249] <=  8'h00;      memory[24250] <=  8'h00;      memory[24251] <=  8'h00;      memory[24252] <=  8'h00;      memory[24253] <=  8'h00;      memory[24254] <=  8'h00;      memory[24255] <=  8'h00;      memory[24256] <=  8'h00;      memory[24257] <=  8'h00;      memory[24258] <=  8'h00;      memory[24259] <=  8'h00;      memory[24260] <=  8'h00;      memory[24261] <=  8'h00;      memory[24262] <=  8'h00;      memory[24263] <=  8'h00;      memory[24264] <=  8'h00;      memory[24265] <=  8'h00;      memory[24266] <=  8'h00;      memory[24267] <=  8'h00;      memory[24268] <=  8'h00;      memory[24269] <=  8'h00;      memory[24270] <=  8'h00;      memory[24271] <=  8'h00;      memory[24272] <=  8'h00;      memory[24273] <=  8'h00;      memory[24274] <=  8'h00;      memory[24275] <=  8'h00;      memory[24276] <=  8'h00;      memory[24277] <=  8'h00;      memory[24278] <=  8'h00;      memory[24279] <=  8'h00;      memory[24280] <=  8'h00;      memory[24281] <=  8'h00;      memory[24282] <=  8'h00;      memory[24283] <=  8'h00;      memory[24284] <=  8'h00;      memory[24285] <=  8'h00;      memory[24286] <=  8'h00;      memory[24287] <=  8'h00;      memory[24288] <=  8'h00;      memory[24289] <=  8'h00;      memory[24290] <=  8'h00;      memory[24291] <=  8'h00;      memory[24292] <=  8'h00;      memory[24293] <=  8'h00;      memory[24294] <=  8'h00;      memory[24295] <=  8'h00;      memory[24296] <=  8'h00;      memory[24297] <=  8'h00;      memory[24298] <=  8'h00;      memory[24299] <=  8'h00;      memory[24300] <=  8'h00;      memory[24301] <=  8'h00;      memory[24302] <=  8'h00;      memory[24303] <=  8'h00;      memory[24304] <=  8'h00;      memory[24305] <=  8'h00;      memory[24306] <=  8'h00;      memory[24307] <=  8'h00;      memory[24308] <=  8'h00;      memory[24309] <=  8'h00;      memory[24310] <=  8'h00;      memory[24311] <=  8'h00;      memory[24312] <=  8'h00;      memory[24313] <=  8'h00;      memory[24314] <=  8'h00;      memory[24315] <=  8'h00;      memory[24316] <=  8'h00;      memory[24317] <=  8'h00;      memory[24318] <=  8'h00;      memory[24319] <=  8'h00;      memory[24320] <=  8'h00;      memory[24321] <=  8'h00;      memory[24322] <=  8'h00;      memory[24323] <=  8'h00;      memory[24324] <=  8'h00;      memory[24325] <=  8'h00;      memory[24326] <=  8'h00;      memory[24327] <=  8'h00;      memory[24328] <=  8'h00;      memory[24329] <=  8'h00;      memory[24330] <=  8'h00;      memory[24331] <=  8'h00;      memory[24332] <=  8'h00;      memory[24333] <=  8'h00;      memory[24334] <=  8'h00;      memory[24335] <=  8'h00;      memory[24336] <=  8'h00;      memory[24337] <=  8'h00;      memory[24338] <=  8'h00;      memory[24339] <=  8'h00;      memory[24340] <=  8'h00;      memory[24341] <=  8'h00;      memory[24342] <=  8'h00;      memory[24343] <=  8'h00;      memory[24344] <=  8'h00;      memory[24345] <=  8'h00;      memory[24346] <=  8'h00;      memory[24347] <=  8'h00;      memory[24348] <=  8'h00;      memory[24349] <=  8'h00;      memory[24350] <=  8'h00;      memory[24351] <=  8'h00;      memory[24352] <=  8'h00;      memory[24353] <=  8'h00;      memory[24354] <=  8'h00;      memory[24355] <=  8'h00;      memory[24356] <=  8'h00;      memory[24357] <=  8'h00;      memory[24358] <=  8'h00;      memory[24359] <=  8'h00;      memory[24360] <=  8'h00;      memory[24361] <=  8'h00;      memory[24362] <=  8'h00;      memory[24363] <=  8'h00;      memory[24364] <=  8'h00;      memory[24365] <=  8'h00;      memory[24366] <=  8'h00;      memory[24367] <=  8'h00;      memory[24368] <=  8'h00;      memory[24369] <=  8'h00;      memory[24370] <=  8'h00;      memory[24371] <=  8'h00;      memory[24372] <=  8'h00;      memory[24373] <=  8'h00;      memory[24374] <=  8'h00;      memory[24375] <=  8'h00;      memory[24376] <=  8'h00;      memory[24377] <=  8'h00;      memory[24378] <=  8'h00;      memory[24379] <=  8'h00;      memory[24380] <=  8'h00;      memory[24381] <=  8'h00;      memory[24382] <=  8'h00;      memory[24383] <=  8'h00;      memory[24384] <=  8'h00;      memory[24385] <=  8'h00;      memory[24386] <=  8'h00;      memory[24387] <=  8'h00;      memory[24388] <=  8'h00;      memory[24389] <=  8'h00;      memory[24390] <=  8'h00;      memory[24391] <=  8'h00;      memory[24392] <=  8'h00;      memory[24393] <=  8'h00;      memory[24394] <=  8'h00;      memory[24395] <=  8'h00;      memory[24396] <=  8'h00;      memory[24397] <=  8'h00;      memory[24398] <=  8'h00;      memory[24399] <=  8'h00;      memory[24400] <=  8'h00;      memory[24401] <=  8'h00;      memory[24402] <=  8'h00;      memory[24403] <=  8'h00;      memory[24404] <=  8'h00;      memory[24405] <=  8'h00;      memory[24406] <=  8'h00;      memory[24407] <=  8'h00;      memory[24408] <=  8'h00;      memory[24409] <=  8'h00;      memory[24410] <=  8'h00;      memory[24411] <=  8'h00;      memory[24412] <=  8'h00;      memory[24413] <=  8'h00;      memory[24414] <=  8'h00;      memory[24415] <=  8'h00;      memory[24416] <=  8'h00;      memory[24417] <=  8'h00;      memory[24418] <=  8'h00;      memory[24419] <=  8'h00;      memory[24420] <=  8'h00;      memory[24421] <=  8'h00;      memory[24422] <=  8'h00;      memory[24423] <=  8'h00;      memory[24424] <=  8'h00;      memory[24425] <=  8'h00;      memory[24426] <=  8'h00;      memory[24427] <=  8'h00;      memory[24428] <=  8'h00;      memory[24429] <=  8'h00;      memory[24430] <=  8'h00;      memory[24431] <=  8'h00;      memory[24432] <=  8'h00;      memory[24433] <=  8'h00;      memory[24434] <=  8'h00;      memory[24435] <=  8'h00;      memory[24436] <=  8'h00;      memory[24437] <=  8'h00;      memory[24438] <=  8'h00;      memory[24439] <=  8'h00;      memory[24440] <=  8'h00;      memory[24441] <=  8'h00;      memory[24442] <=  8'h00;      memory[24443] <=  8'h00;      memory[24444] <=  8'h00;      memory[24445] <=  8'h00;      memory[24446] <=  8'h00;      memory[24447] <=  8'h00;      memory[24448] <=  8'h00;      memory[24449] <=  8'h00;      memory[24450] <=  8'h00;      memory[24451] <=  8'h00;      memory[24452] <=  8'h00;      memory[24453] <=  8'h00;      memory[24454] <=  8'h00;      memory[24455] <=  8'h00;      memory[24456] <=  8'h00;      memory[24457] <=  8'h00;      memory[24458] <=  8'h00;      memory[24459] <=  8'h00;      memory[24460] <=  8'h00;      memory[24461] <=  8'h00;      memory[24462] <=  8'h00;      memory[24463] <=  8'h00;      memory[24464] <=  8'h00;      memory[24465] <=  8'h00;      memory[24466] <=  8'h00;      memory[24467] <=  8'h00;      memory[24468] <=  8'h00;      memory[24469] <=  8'h00;      memory[24470] <=  8'h00;      memory[24471] <=  8'h00;      memory[24472] <=  8'h00;      memory[24473] <=  8'h00;      memory[24474] <=  8'h00;      memory[24475] <=  8'h00;      memory[24476] <=  8'h00;      memory[24477] <=  8'h00;      memory[24478] <=  8'h00;      memory[24479] <=  8'h00;      memory[24480] <=  8'h00;      memory[24481] <=  8'h00;      memory[24482] <=  8'h00;      memory[24483] <=  8'h00;      memory[24484] <=  8'h00;      memory[24485] <=  8'h00;      memory[24486] <=  8'h00;      memory[24487] <=  8'h00;      memory[24488] <=  8'h00;      memory[24489] <=  8'h00;      memory[24490] <=  8'h00;      memory[24491] <=  8'h00;      memory[24492] <=  8'h00;      memory[24493] <=  8'h00;      memory[24494] <=  8'h00;      memory[24495] <=  8'h00;      memory[24496] <=  8'h00;      memory[24497] <=  8'h00;      memory[24498] <=  8'h00;      memory[24499] <=  8'h00;      memory[24500] <=  8'h00;      memory[24501] <=  8'h00;      memory[24502] <=  8'h00;      memory[24503] <=  8'h00;      memory[24504] <=  8'h00;      memory[24505] <=  8'h00;      memory[24506] <=  8'h00;      memory[24507] <=  8'h00;      memory[24508] <=  8'h00;      memory[24509] <=  8'h00;      memory[24510] <=  8'h00;      memory[24511] <=  8'h00;      memory[24512] <=  8'h00;      memory[24513] <=  8'h00;      memory[24514] <=  8'h00;      memory[24515] <=  8'h00;      memory[24516] <=  8'h00;      memory[24517] <=  8'h00;      memory[24518] <=  8'h00;      memory[24519] <=  8'h00;      memory[24520] <=  8'h00;      memory[24521] <=  8'h00;      memory[24522] <=  8'h00;      memory[24523] <=  8'h00;      memory[24524] <=  8'h00;      memory[24525] <=  8'h00;      memory[24526] <=  8'h00;      memory[24527] <=  8'h00;      memory[24528] <=  8'h00;      memory[24529] <=  8'h00;      memory[24530] <=  8'h00;      memory[24531] <=  8'h00;      memory[24532] <=  8'h00;      memory[24533] <=  8'h00;      memory[24534] <=  8'h00;      memory[24535] <=  8'h00;      memory[24536] <=  8'h00;      memory[24537] <=  8'h00;      memory[24538] <=  8'h00;      memory[24539] <=  8'h00;      memory[24540] <=  8'h00;      memory[24541] <=  8'h00;      memory[24542] <=  8'h00;      memory[24543] <=  8'h00;      memory[24544] <=  8'h00;      memory[24545] <=  8'h00;      memory[24546] <=  8'h00;      memory[24547] <=  8'h00;      memory[24548] <=  8'h00;      memory[24549] <=  8'h00;      memory[24550] <=  8'h00;      memory[24551] <=  8'h00;      memory[24552] <=  8'h00;      memory[24553] <=  8'h00;      memory[24554] <=  8'h00;      memory[24555] <=  8'h00;      memory[24556] <=  8'h00;      memory[24557] <=  8'h00;      memory[24558] <=  8'h00;      memory[24559] <=  8'h00;      memory[24560] <=  8'h00;      memory[24561] <=  8'h00;      memory[24562] <=  8'h00;      memory[24563] <=  8'h00;      memory[24564] <=  8'h00;      memory[24565] <=  8'h00;      memory[24566] <=  8'h00;      memory[24567] <=  8'h00;      memory[24568] <=  8'h00;      memory[24569] <=  8'h00;      memory[24570] <=  8'h00;      memory[24571] <=  8'h00;      memory[24572] <=  8'h00;      memory[24573] <=  8'h00;      memory[24574] <=  8'h00;      memory[24575] <=  8'h00;      memory[24576] <=  8'h00;      memory[24577] <=  8'h00;      memory[24578] <=  8'h00;      memory[24579] <=  8'h00;      memory[24580] <=  8'h00;      memory[24581] <=  8'h00;      memory[24582] <=  8'h00;      memory[24583] <=  8'h00;      memory[24584] <=  8'h00;      memory[24585] <=  8'h00;      memory[24586] <=  8'h00;      memory[24587] <=  8'h00;      memory[24588] <=  8'h00;      memory[24589] <=  8'h00;      memory[24590] <=  8'h00;      memory[24591] <=  8'h00;      memory[24592] <=  8'h00;      memory[24593] <=  8'h00;      memory[24594] <=  8'h00;      memory[24595] <=  8'h00;      memory[24596] <=  8'h00;      memory[24597] <=  8'h00;      memory[24598] <=  8'h00;      memory[24599] <=  8'h00;      memory[24600] <=  8'h00;      memory[24601] <=  8'h00;      memory[24602] <=  8'h00;      memory[24603] <=  8'h00;      memory[24604] <=  8'h00;      memory[24605] <=  8'h00;      memory[24606] <=  8'h00;      memory[24607] <=  8'h00;      memory[24608] <=  8'h00;      memory[24609] <=  8'h00;      memory[24610] <=  8'h00;      memory[24611] <=  8'h00;      memory[24612] <=  8'h00;      memory[24613] <=  8'h00;      memory[24614] <=  8'h00;      memory[24615] <=  8'h00;      memory[24616] <=  8'h00;      memory[24617] <=  8'h00;      memory[24618] <=  8'h00;      memory[24619] <=  8'h00;      memory[24620] <=  8'h00;      memory[24621] <=  8'h00;      memory[24622] <=  8'h00;      memory[24623] <=  8'h00;      memory[24624] <=  8'h00;      memory[24625] <=  8'h00;      memory[24626] <=  8'h00;      memory[24627] <=  8'h00;      memory[24628] <=  8'h00;      memory[24629] <=  8'h00;      memory[24630] <=  8'h00;      memory[24631] <=  8'h00;      memory[24632] <=  8'h00;      memory[24633] <=  8'h00;      memory[24634] <=  8'h00;      memory[24635] <=  8'h00;      memory[24636] <=  8'h00;      memory[24637] <=  8'h00;      memory[24638] <=  8'h00;      memory[24639] <=  8'h00;      memory[24640] <=  8'h00;      memory[24641] <=  8'h00;      memory[24642] <=  8'h00;      memory[24643] <=  8'h00;      memory[24644] <=  8'h00;      memory[24645] <=  8'h00;      memory[24646] <=  8'h00;      memory[24647] <=  8'h00;      memory[24648] <=  8'h00;      memory[24649] <=  8'h00;      memory[24650] <=  8'h00;      memory[24651] <=  8'h00;      memory[24652] <=  8'h00;      memory[24653] <=  8'h00;      memory[24654] <=  8'h00;      memory[24655] <=  8'h00;      memory[24656] <=  8'h00;      memory[24657] <=  8'h00;      memory[24658] <=  8'h00;      memory[24659] <=  8'h00;      memory[24660] <=  8'h00;      memory[24661] <=  8'h00;      memory[24662] <=  8'h00;      memory[24663] <=  8'h00;      memory[24664] <=  8'h00;      memory[24665] <=  8'h00;      memory[24666] <=  8'h00;      memory[24667] <=  8'h00;      memory[24668] <=  8'h00;      memory[24669] <=  8'h00;      memory[24670] <=  8'h00;      memory[24671] <=  8'h00;      memory[24672] <=  8'h00;      memory[24673] <=  8'h00;      memory[24674] <=  8'h00;      memory[24675] <=  8'h00;      memory[24676] <=  8'h00;      memory[24677] <=  8'h00;      memory[24678] <=  8'h00;      memory[24679] <=  8'h00;      memory[24680] <=  8'h00;      memory[24681] <=  8'h00;      memory[24682] <=  8'h00;      memory[24683] <=  8'h00;      memory[24684] <=  8'h00;      memory[24685] <=  8'h00;      memory[24686] <=  8'h00;      memory[24687] <=  8'h00;      memory[24688] <=  8'h00;      memory[24689] <=  8'h00;      memory[24690] <=  8'h00;      memory[24691] <=  8'h00;      memory[24692] <=  8'h00;      memory[24693] <=  8'h00;      memory[24694] <=  8'h00;      memory[24695] <=  8'h00;      memory[24696] <=  8'h00;      memory[24697] <=  8'h00;      memory[24698] <=  8'h00;      memory[24699] <=  8'h00;      memory[24700] <=  8'h00;      memory[24701] <=  8'h00;      memory[24702] <=  8'h00;      memory[24703] <=  8'h00;      memory[24704] <=  8'h00;      memory[24705] <=  8'h00;      memory[24706] <=  8'h00;      memory[24707] <=  8'h00;      memory[24708] <=  8'h00;      memory[24709] <=  8'h00;      memory[24710] <=  8'h00;      memory[24711] <=  8'h00;      memory[24712] <=  8'h00;      memory[24713] <=  8'h00;      memory[24714] <=  8'h00;      memory[24715] <=  8'h00;      memory[24716] <=  8'h00;      memory[24717] <=  8'h00;      memory[24718] <=  8'h00;      memory[24719] <=  8'h00;      memory[24720] <=  8'h00;      memory[24721] <=  8'h00;      memory[24722] <=  8'h00;      memory[24723] <=  8'h00;      memory[24724] <=  8'h00;      memory[24725] <=  8'h00;      memory[24726] <=  8'h00;      memory[24727] <=  8'h00;      memory[24728] <=  8'h00;      memory[24729] <=  8'h00;      memory[24730] <=  8'h00;      memory[24731] <=  8'h00;      memory[24732] <=  8'h00;      memory[24733] <=  8'h00;      memory[24734] <=  8'h00;      memory[24735] <=  8'h00;      memory[24736] <=  8'h00;      memory[24737] <=  8'h00;      memory[24738] <=  8'h00;      memory[24739] <=  8'h00;      memory[24740] <=  8'h00;      memory[24741] <=  8'h00;      memory[24742] <=  8'h00;      memory[24743] <=  8'h00;      memory[24744] <=  8'h00;      memory[24745] <=  8'h00;      memory[24746] <=  8'h00;      memory[24747] <=  8'h00;      memory[24748] <=  8'h00;      memory[24749] <=  8'h00;      memory[24750] <=  8'h00;      memory[24751] <=  8'h00;      memory[24752] <=  8'h00;      memory[24753] <=  8'h00;      memory[24754] <=  8'h00;      memory[24755] <=  8'h00;      memory[24756] <=  8'h00;      memory[24757] <=  8'h00;      memory[24758] <=  8'h00;      memory[24759] <=  8'h00;      memory[24760] <=  8'h00;      memory[24761] <=  8'h00;      memory[24762] <=  8'h00;      memory[24763] <=  8'h00;      memory[24764] <=  8'h00;      memory[24765] <=  8'h00;      memory[24766] <=  8'h00;      memory[24767] <=  8'h00;      memory[24768] <=  8'h00;      memory[24769] <=  8'h00;      memory[24770] <=  8'h00;      memory[24771] <=  8'h00;      memory[24772] <=  8'h00;      memory[24773] <=  8'h00;      memory[24774] <=  8'h00;      memory[24775] <=  8'h00;      memory[24776] <=  8'h00;      memory[24777] <=  8'h00;      memory[24778] <=  8'h00;      memory[24779] <=  8'h00;      memory[24780] <=  8'h00;      memory[24781] <=  8'h00;      memory[24782] <=  8'h00;      memory[24783] <=  8'h00;      memory[24784] <=  8'h00;      memory[24785] <=  8'h00;      memory[24786] <=  8'h00;      memory[24787] <=  8'h00;      memory[24788] <=  8'h00;      memory[24789] <=  8'h00;      memory[24790] <=  8'h00;      memory[24791] <=  8'h00;      memory[24792] <=  8'h00;      memory[24793] <=  8'h00;      memory[24794] <=  8'h00;      memory[24795] <=  8'h00;      memory[24796] <=  8'h00;      memory[24797] <=  8'h00;      memory[24798] <=  8'h00;      memory[24799] <=  8'h00;      memory[24800] <=  8'h00;      memory[24801] <=  8'h00;      memory[24802] <=  8'h00;      memory[24803] <=  8'h00;      memory[24804] <=  8'h00;      memory[24805] <=  8'h00;      memory[24806] <=  8'h00;      memory[24807] <=  8'h00;      memory[24808] <=  8'h00;      memory[24809] <=  8'h00;      memory[24810] <=  8'h00;      memory[24811] <=  8'h00;      memory[24812] <=  8'h00;      memory[24813] <=  8'h00;      memory[24814] <=  8'h00;      memory[24815] <=  8'h00;      memory[24816] <=  8'h00;      memory[24817] <=  8'h00;      memory[24818] <=  8'h00;      memory[24819] <=  8'h00;      memory[24820] <=  8'h00;      memory[24821] <=  8'h00;      memory[24822] <=  8'h00;      memory[24823] <=  8'h00;      memory[24824] <=  8'h00;      memory[24825] <=  8'h00;      memory[24826] <=  8'h00;      memory[24827] <=  8'h00;      memory[24828] <=  8'h00;      memory[24829] <=  8'h00;      memory[24830] <=  8'h00;      memory[24831] <=  8'h00;      memory[24832] <=  8'h00;      memory[24833] <=  8'h00;      memory[24834] <=  8'h00;      memory[24835] <=  8'h00;      memory[24836] <=  8'h00;      memory[24837] <=  8'h00;      memory[24838] <=  8'h00;      memory[24839] <=  8'h00;      memory[24840] <=  8'h00;      memory[24841] <=  8'h00;      memory[24842] <=  8'h00;      memory[24843] <=  8'h00;      memory[24844] <=  8'h00;      memory[24845] <=  8'h00;      memory[24846] <=  8'h00;      memory[24847] <=  8'h00;      memory[24848] <=  8'h00;      memory[24849] <=  8'h00;      memory[24850] <=  8'h00;      memory[24851] <=  8'h00;      memory[24852] <=  8'h00;      memory[24853] <=  8'h00;      memory[24854] <=  8'h00;      memory[24855] <=  8'h00;      memory[24856] <=  8'h00;      memory[24857] <=  8'h00;      memory[24858] <=  8'h00;      memory[24859] <=  8'h00;      memory[24860] <=  8'h00;      memory[24861] <=  8'h00;      memory[24862] <=  8'h00;      memory[24863] <=  8'h00;      memory[24864] <=  8'h00;      memory[24865] <=  8'h00;      memory[24866] <=  8'h00;      memory[24867] <=  8'h00;      memory[24868] <=  8'h00;      memory[24869] <=  8'h00;      memory[24870] <=  8'h00;      memory[24871] <=  8'h00;      memory[24872] <=  8'h00;      memory[24873] <=  8'h00;      memory[24874] <=  8'h00;      memory[24875] <=  8'h00;      memory[24876] <=  8'h00;      memory[24877] <=  8'h00;      memory[24878] <=  8'h00;      memory[24879] <=  8'h00;      memory[24880] <=  8'h00;      memory[24881] <=  8'h00;      memory[24882] <=  8'h00;      memory[24883] <=  8'h00;      memory[24884] <=  8'h00;      memory[24885] <=  8'h00;      memory[24886] <=  8'h00;      memory[24887] <=  8'h00;      memory[24888] <=  8'h00;      memory[24889] <=  8'h00;      memory[24890] <=  8'h00;      memory[24891] <=  8'h00;      memory[24892] <=  8'h00;      memory[24893] <=  8'h00;      memory[24894] <=  8'h00;      memory[24895] <=  8'h00;      memory[24896] <=  8'h00;      memory[24897] <=  8'h00;      memory[24898] <=  8'h00;      memory[24899] <=  8'h00;      memory[24900] <=  8'h00;      memory[24901] <=  8'h00;      memory[24902] <=  8'h00;      memory[24903] <=  8'h00;      memory[24904] <=  8'h00;      memory[24905] <=  8'h00;      memory[24906] <=  8'h00;      memory[24907] <=  8'h00;      memory[24908] <=  8'h00;      memory[24909] <=  8'h00;      memory[24910] <=  8'h00;      memory[24911] <=  8'h00;      memory[24912] <=  8'h00;      memory[24913] <=  8'h00;      memory[24914] <=  8'h00;      memory[24915] <=  8'h00;      memory[24916] <=  8'h00;      memory[24917] <=  8'h00;      memory[24918] <=  8'h00;      memory[24919] <=  8'h00;      memory[24920] <=  8'h00;      memory[24921] <=  8'h00;      memory[24922] <=  8'h00;      memory[24923] <=  8'h00;      memory[24924] <=  8'h00;      memory[24925] <=  8'h00;      memory[24926] <=  8'h00;      memory[24927] <=  8'h00;      memory[24928] <=  8'h00;      memory[24929] <=  8'h00;      memory[24930] <=  8'h00;      memory[24931] <=  8'h00;      memory[24932] <=  8'h00;      memory[24933] <=  8'h00;      memory[24934] <=  8'h00;      memory[24935] <=  8'h00;      memory[24936] <=  8'h00;      memory[24937] <=  8'h00;      memory[24938] <=  8'h00;      memory[24939] <=  8'h00;      memory[24940] <=  8'h00;      memory[24941] <=  8'h00;      memory[24942] <=  8'h00;      memory[24943] <=  8'h00;      memory[24944] <=  8'h00;      memory[24945] <=  8'h00;      memory[24946] <=  8'h00;      memory[24947] <=  8'h00;      memory[24948] <=  8'h00;      memory[24949] <=  8'h00;      memory[24950] <=  8'h00;      memory[24951] <=  8'h00;      memory[24952] <=  8'h00;      memory[24953] <=  8'h00;      memory[24954] <=  8'h00;      memory[24955] <=  8'h00;      memory[24956] <=  8'h00;      memory[24957] <=  8'h00;      memory[24958] <=  8'h00;      memory[24959] <=  8'h00;      memory[24960] <=  8'h00;      memory[24961] <=  8'h00;      memory[24962] <=  8'h00;      memory[24963] <=  8'h00;      memory[24964] <=  8'h00;      memory[24965] <=  8'h00;      memory[24966] <=  8'h00;      memory[24967] <=  8'h00;      memory[24968] <=  8'h00;      memory[24969] <=  8'h00;      memory[24970] <=  8'h00;      memory[24971] <=  8'h00;      memory[24972] <=  8'h00;      memory[24973] <=  8'h00;      memory[24974] <=  8'h00;      memory[24975] <=  8'h00;      memory[24976] <=  8'h00;      memory[24977] <=  8'h00;      memory[24978] <=  8'h00;      memory[24979] <=  8'h00;      memory[24980] <=  8'h00;      memory[24981] <=  8'h00;      memory[24982] <=  8'h00;      memory[24983] <=  8'h00;      memory[24984] <=  8'h00;      memory[24985] <=  8'h00;      memory[24986] <=  8'h00;      memory[24987] <=  8'h00;      memory[24988] <=  8'h00;      memory[24989] <=  8'h00;      memory[24990] <=  8'h00;      memory[24991] <=  8'h00;      memory[24992] <=  8'h00;      memory[24993] <=  8'h00;      memory[24994] <=  8'h00;      memory[24995] <=  8'h00;      memory[24996] <=  8'h00;      memory[24997] <=  8'h00;      memory[24998] <=  8'h00;      memory[24999] <=  8'h00;      memory[25000] <=  8'h00;      memory[25001] <=  8'h00;      memory[25002] <=  8'h00;      memory[25003] <=  8'h00;      memory[25004] <=  8'h00;      memory[25005] <=  8'h00;      memory[25006] <=  8'h00;      memory[25007] <=  8'h00;      memory[25008] <=  8'h00;      memory[25009] <=  8'h00;      memory[25010] <=  8'h00;      memory[25011] <=  8'h00;      memory[25012] <=  8'h00;      memory[25013] <=  8'h00;      memory[25014] <=  8'h00;      memory[25015] <=  8'h00;      memory[25016] <=  8'h00;      memory[25017] <=  8'h00;      memory[25018] <=  8'h00;      memory[25019] <=  8'h00;      memory[25020] <=  8'h00;      memory[25021] <=  8'h00;      memory[25022] <=  8'h00;      memory[25023] <=  8'h00;      memory[25024] <=  8'h00;      memory[25025] <=  8'h00;      memory[25026] <=  8'h00;      memory[25027] <=  8'h00;      memory[25028] <=  8'h00;      memory[25029] <=  8'h00;      memory[25030] <=  8'h00;      memory[25031] <=  8'h00;      memory[25032] <=  8'h00;      memory[25033] <=  8'h00;      memory[25034] <=  8'h00;      memory[25035] <=  8'h00;      memory[25036] <=  8'h00;      memory[25037] <=  8'h00;      memory[25038] <=  8'h00;      memory[25039] <=  8'h00;      memory[25040] <=  8'h00;      memory[25041] <=  8'h00;      memory[25042] <=  8'h00;      memory[25043] <=  8'h00;      memory[25044] <=  8'h00;      memory[25045] <=  8'h00;      memory[25046] <=  8'h00;      memory[25047] <=  8'h00;      memory[25048] <=  8'h00;      memory[25049] <=  8'h00;      memory[25050] <=  8'h00;      memory[25051] <=  8'h00;      memory[25052] <=  8'h00;      memory[25053] <=  8'h00;      memory[25054] <=  8'h00;      memory[25055] <=  8'h00;      memory[25056] <=  8'h00;      memory[25057] <=  8'h00;      memory[25058] <=  8'h00;      memory[25059] <=  8'h00;      memory[25060] <=  8'h00;      memory[25061] <=  8'h00;      memory[25062] <=  8'h00;      memory[25063] <=  8'h00;      memory[25064] <=  8'h00;      memory[25065] <=  8'h00;      memory[25066] <=  8'h00;      memory[25067] <=  8'h00;      memory[25068] <=  8'h00;      memory[25069] <=  8'h00;      memory[25070] <=  8'h00;      memory[25071] <=  8'h00;      memory[25072] <=  8'h00;      memory[25073] <=  8'h00;      memory[25074] <=  8'h00;      memory[25075] <=  8'h00;      memory[25076] <=  8'h00;      memory[25077] <=  8'h00;      memory[25078] <=  8'h00;      memory[25079] <=  8'h00;      memory[25080] <=  8'h00;      memory[25081] <=  8'h00;      memory[25082] <=  8'h00;      memory[25083] <=  8'h00;      memory[25084] <=  8'h00;      memory[25085] <=  8'h00;      memory[25086] <=  8'h00;      memory[25087] <=  8'h00;      memory[25088] <=  8'h00;      memory[25089] <=  8'h00;      memory[25090] <=  8'h00;      memory[25091] <=  8'h00;      memory[25092] <=  8'h00;      memory[25093] <=  8'h00;      memory[25094] <=  8'h00;      memory[25095] <=  8'h00;      memory[25096] <=  8'h00;      memory[25097] <=  8'h00;      memory[25098] <=  8'h00;      memory[25099] <=  8'h00;      memory[25100] <=  8'h00;      memory[25101] <=  8'h00;      memory[25102] <=  8'h00;      memory[25103] <=  8'h00;      memory[25104] <=  8'h00;      memory[25105] <=  8'h00;      memory[25106] <=  8'h00;      memory[25107] <=  8'h00;      memory[25108] <=  8'h00;      memory[25109] <=  8'h00;      memory[25110] <=  8'h00;      memory[25111] <=  8'h00;      memory[25112] <=  8'h00;      memory[25113] <=  8'h00;      memory[25114] <=  8'h00;      memory[25115] <=  8'h00;      memory[25116] <=  8'h00;      memory[25117] <=  8'h00;      memory[25118] <=  8'h00;      memory[25119] <=  8'h00;      memory[25120] <=  8'h00;      memory[25121] <=  8'h00;      memory[25122] <=  8'h00;      memory[25123] <=  8'h00;      memory[25124] <=  8'h00;      memory[25125] <=  8'h00;      memory[25126] <=  8'h00;      memory[25127] <=  8'h00;      memory[25128] <=  8'h00;      memory[25129] <=  8'h00;      memory[25130] <=  8'h00;      memory[25131] <=  8'h00;      memory[25132] <=  8'h00;      memory[25133] <=  8'h00;      memory[25134] <=  8'h00;      memory[25135] <=  8'h00;      memory[25136] <=  8'h00;      memory[25137] <=  8'h00;      memory[25138] <=  8'h00;      memory[25139] <=  8'h00;      memory[25140] <=  8'h00;      memory[25141] <=  8'h00;      memory[25142] <=  8'h00;      memory[25143] <=  8'h00;      memory[25144] <=  8'h00;      memory[25145] <=  8'h00;      memory[25146] <=  8'h00;      memory[25147] <=  8'h00;      memory[25148] <=  8'h00;      memory[25149] <=  8'h00;      memory[25150] <=  8'h00;      memory[25151] <=  8'h00;      memory[25152] <=  8'h00;      memory[25153] <=  8'h00;      memory[25154] <=  8'h00;      memory[25155] <=  8'h00;      memory[25156] <=  8'h00;      memory[25157] <=  8'h00;      memory[25158] <=  8'h00;      memory[25159] <=  8'h00;      memory[25160] <=  8'h00;      memory[25161] <=  8'h00;      memory[25162] <=  8'h00;      memory[25163] <=  8'h00;      memory[25164] <=  8'h00;      memory[25165] <=  8'h00;      memory[25166] <=  8'h00;      memory[25167] <=  8'h00;      memory[25168] <=  8'h00;      memory[25169] <=  8'h00;      memory[25170] <=  8'h00;      memory[25171] <=  8'h00;      memory[25172] <=  8'h00;      memory[25173] <=  8'h00;      memory[25174] <=  8'h00;      memory[25175] <=  8'h00;      memory[25176] <=  8'h00;      memory[25177] <=  8'h00;      memory[25178] <=  8'h00;      memory[25179] <=  8'h00;      memory[25180] <=  8'h00;      memory[25181] <=  8'h00;      memory[25182] <=  8'h00;      memory[25183] <=  8'h00;      memory[25184] <=  8'h00;      memory[25185] <=  8'h00;      memory[25186] <=  8'h00;      memory[25187] <=  8'h00;      memory[25188] <=  8'h00;      memory[25189] <=  8'h00;      memory[25190] <=  8'h00;      memory[25191] <=  8'h00;      memory[25192] <=  8'h00;      memory[25193] <=  8'h00;      memory[25194] <=  8'h00;      memory[25195] <=  8'h00;      memory[25196] <=  8'h00;      memory[25197] <=  8'h00;      memory[25198] <=  8'h00;      memory[25199] <=  8'h00;      memory[25200] <=  8'h00;      memory[25201] <=  8'h00;      memory[25202] <=  8'h00;      memory[25203] <=  8'h00;      memory[25204] <=  8'h00;      memory[25205] <=  8'h00;      memory[25206] <=  8'h00;      memory[25207] <=  8'h00;      memory[25208] <=  8'h00;      memory[25209] <=  8'h00;      memory[25210] <=  8'h00;      memory[25211] <=  8'h00;      memory[25212] <=  8'h00;      memory[25213] <=  8'h00;      memory[25214] <=  8'h00;      memory[25215] <=  8'h00;      memory[25216] <=  8'h00;      memory[25217] <=  8'h00;      memory[25218] <=  8'h00;      memory[25219] <=  8'h00;      memory[25220] <=  8'h00;      memory[25221] <=  8'h00;      memory[25222] <=  8'h00;      memory[25223] <=  8'h00;      memory[25224] <=  8'h00;      memory[25225] <=  8'h00;      memory[25226] <=  8'h00;      memory[25227] <=  8'h00;      memory[25228] <=  8'h00;      memory[25229] <=  8'h00;      memory[25230] <=  8'h00;      memory[25231] <=  8'h00;      memory[25232] <=  8'h00;      memory[25233] <=  8'h00;      memory[25234] <=  8'h00;      memory[25235] <=  8'h00;      memory[25236] <=  8'h00;      memory[25237] <=  8'h00;      memory[25238] <=  8'h00;      memory[25239] <=  8'h00;      memory[25240] <=  8'h00;      memory[25241] <=  8'h00;      memory[25242] <=  8'h00;      memory[25243] <=  8'h00;      memory[25244] <=  8'h00;      memory[25245] <=  8'h00;      memory[25246] <=  8'h00;      memory[25247] <=  8'h00;      memory[25248] <=  8'h00;      memory[25249] <=  8'h00;      memory[25250] <=  8'h00;      memory[25251] <=  8'h00;      memory[25252] <=  8'h00;      memory[25253] <=  8'h00;      memory[25254] <=  8'h00;      memory[25255] <=  8'h00;      memory[25256] <=  8'h00;      memory[25257] <=  8'h00;      memory[25258] <=  8'h00;      memory[25259] <=  8'h00;      memory[25260] <=  8'h00;      memory[25261] <=  8'h00;      memory[25262] <=  8'h00;      memory[25263] <=  8'h00;      memory[25264] <=  8'h00;      memory[25265] <=  8'h00;      memory[25266] <=  8'h00;      memory[25267] <=  8'h00;      memory[25268] <=  8'h00;      memory[25269] <=  8'h00;      memory[25270] <=  8'h00;      memory[25271] <=  8'h00;      memory[25272] <=  8'h00;      memory[25273] <=  8'h00;      memory[25274] <=  8'h00;      memory[25275] <=  8'h00;      memory[25276] <=  8'h00;      memory[25277] <=  8'h00;      memory[25278] <=  8'h00;      memory[25279] <=  8'h00;      memory[25280] <=  8'h00;      memory[25281] <=  8'h00;      memory[25282] <=  8'h00;      memory[25283] <=  8'h00;      memory[25284] <=  8'h00;      memory[25285] <=  8'h00;      memory[25286] <=  8'h00;      memory[25287] <=  8'h00;      memory[25288] <=  8'h00;      memory[25289] <=  8'h00;      memory[25290] <=  8'h00;      memory[25291] <=  8'h00;      memory[25292] <=  8'h00;      memory[25293] <=  8'h00;      memory[25294] <=  8'h00;      memory[25295] <=  8'h00;      memory[25296] <=  8'h00;      memory[25297] <=  8'h00;      memory[25298] <=  8'h00;      memory[25299] <=  8'h00;      memory[25300] <=  8'h00;      memory[25301] <=  8'h00;      memory[25302] <=  8'h00;      memory[25303] <=  8'h00;      memory[25304] <=  8'h00;      memory[25305] <=  8'h00;      memory[25306] <=  8'h00;      memory[25307] <=  8'h00;      memory[25308] <=  8'h00;      memory[25309] <=  8'h00;      memory[25310] <=  8'h00;      memory[25311] <=  8'h00;      memory[25312] <=  8'h00;      memory[25313] <=  8'h00;      memory[25314] <=  8'h00;      memory[25315] <=  8'h00;      memory[25316] <=  8'h00;      memory[25317] <=  8'h00;      memory[25318] <=  8'h00;      memory[25319] <=  8'h00;      memory[25320] <=  8'h00;      memory[25321] <=  8'h00;      memory[25322] <=  8'h00;      memory[25323] <=  8'h00;      memory[25324] <=  8'h00;      memory[25325] <=  8'h00;      memory[25326] <=  8'h00;      memory[25327] <=  8'h00;      memory[25328] <=  8'h00;      memory[25329] <=  8'h00;      memory[25330] <=  8'h00;      memory[25331] <=  8'h00;      memory[25332] <=  8'h00;      memory[25333] <=  8'h00;      memory[25334] <=  8'h00;      memory[25335] <=  8'h00;      memory[25336] <=  8'h00;      memory[25337] <=  8'h00;      memory[25338] <=  8'h00;      memory[25339] <=  8'h00;      memory[25340] <=  8'h00;      memory[25341] <=  8'h00;      memory[25342] <=  8'h00;      memory[25343] <=  8'h00;      memory[25344] <=  8'h00;      memory[25345] <=  8'h00;      memory[25346] <=  8'h00;      memory[25347] <=  8'h00;      memory[25348] <=  8'h00;      memory[25349] <=  8'h00;      memory[25350] <=  8'h00;      memory[25351] <=  8'h00;      memory[25352] <=  8'h00;      memory[25353] <=  8'h00;      memory[25354] <=  8'h00;      memory[25355] <=  8'h00;      memory[25356] <=  8'h00;      memory[25357] <=  8'h00;      memory[25358] <=  8'h00;      memory[25359] <=  8'h00;      memory[25360] <=  8'h00;      memory[25361] <=  8'h00;      memory[25362] <=  8'h00;      memory[25363] <=  8'h00;      memory[25364] <=  8'h00;      memory[25365] <=  8'h00;      memory[25366] <=  8'h00;      memory[25367] <=  8'h00;      memory[25368] <=  8'h00;      memory[25369] <=  8'h00;      memory[25370] <=  8'h00;      memory[25371] <=  8'h00;      memory[25372] <=  8'h00;      memory[25373] <=  8'h00;      memory[25374] <=  8'h00;      memory[25375] <=  8'h00;      memory[25376] <=  8'h00;      memory[25377] <=  8'h00;      memory[25378] <=  8'h00;      memory[25379] <=  8'h00;      memory[25380] <=  8'h00;      memory[25381] <=  8'h00;      memory[25382] <=  8'h00;      memory[25383] <=  8'h00;      memory[25384] <=  8'h00;      memory[25385] <=  8'h00;      memory[25386] <=  8'h00;      memory[25387] <=  8'h00;      memory[25388] <=  8'h00;      memory[25389] <=  8'h00;      memory[25390] <=  8'h00;      memory[25391] <=  8'h00;      memory[25392] <=  8'h00;      memory[25393] <=  8'h00;      memory[25394] <=  8'h00;      memory[25395] <=  8'h00;      memory[25396] <=  8'h00;      memory[25397] <=  8'h00;      memory[25398] <=  8'h00;      memory[25399] <=  8'h00;      memory[25400] <=  8'h00;      memory[25401] <=  8'h00;      memory[25402] <=  8'h00;      memory[25403] <=  8'h00;      memory[25404] <=  8'h00;      memory[25405] <=  8'h00;      memory[25406] <=  8'h00;      memory[25407] <=  8'h00;      memory[25408] <=  8'h00;      memory[25409] <=  8'h00;      memory[25410] <=  8'h00;      memory[25411] <=  8'h00;      memory[25412] <=  8'h00;      memory[25413] <=  8'h00;      memory[25414] <=  8'h00;      memory[25415] <=  8'h00;      memory[25416] <=  8'h00;      memory[25417] <=  8'h00;      memory[25418] <=  8'h00;      memory[25419] <=  8'h00;      memory[25420] <=  8'h00;      memory[25421] <=  8'h00;      memory[25422] <=  8'h00;      memory[25423] <=  8'h00;      memory[25424] <=  8'h00;      memory[25425] <=  8'h00;      memory[25426] <=  8'h00;      memory[25427] <=  8'h00;      memory[25428] <=  8'h00;      memory[25429] <=  8'h00;      memory[25430] <=  8'h00;      memory[25431] <=  8'h00;      memory[25432] <=  8'h00;      memory[25433] <=  8'h00;      memory[25434] <=  8'h00;      memory[25435] <=  8'h00;      memory[25436] <=  8'h00;      memory[25437] <=  8'h00;      memory[25438] <=  8'h00;      memory[25439] <=  8'h00;      memory[25440] <=  8'h00;      memory[25441] <=  8'h00;      memory[25442] <=  8'h00;      memory[25443] <=  8'h00;      memory[25444] <=  8'h00;      memory[25445] <=  8'h00;      memory[25446] <=  8'h00;      memory[25447] <=  8'h00;      memory[25448] <=  8'h00;      memory[25449] <=  8'h00;      memory[25450] <=  8'h00;      memory[25451] <=  8'h00;      memory[25452] <=  8'h00;      memory[25453] <=  8'h00;      memory[25454] <=  8'h00;      memory[25455] <=  8'h00;      memory[25456] <=  8'h00;      memory[25457] <=  8'h00;      memory[25458] <=  8'h00;      memory[25459] <=  8'h00;      memory[25460] <=  8'h00;      memory[25461] <=  8'h00;      memory[25462] <=  8'h00;      memory[25463] <=  8'h00;      memory[25464] <=  8'h00;      memory[25465] <=  8'h00;      memory[25466] <=  8'h00;      memory[25467] <=  8'h00;      memory[25468] <=  8'h00;      memory[25469] <=  8'h00;      memory[25470] <=  8'h00;      memory[25471] <=  8'h00;      memory[25472] <=  8'h00;      memory[25473] <=  8'h00;      memory[25474] <=  8'h00;      memory[25475] <=  8'h00;      memory[25476] <=  8'h00;      memory[25477] <=  8'h00;      memory[25478] <=  8'h00;      memory[25479] <=  8'h00;      memory[25480] <=  8'h00;      memory[25481] <=  8'h00;      memory[25482] <=  8'h00;      memory[25483] <=  8'h00;      memory[25484] <=  8'h00;      memory[25485] <=  8'h00;      memory[25486] <=  8'h00;      memory[25487] <=  8'h00;      memory[25488] <=  8'h00;      memory[25489] <=  8'h00;      memory[25490] <=  8'h00;      memory[25491] <=  8'h00;      memory[25492] <=  8'h00;      memory[25493] <=  8'h00;      memory[25494] <=  8'h00;      memory[25495] <=  8'h00;      memory[25496] <=  8'h00;      memory[25497] <=  8'h00;      memory[25498] <=  8'h00;      memory[25499] <=  8'h00;      memory[25500] <=  8'h00;      memory[25501] <=  8'h00;      memory[25502] <=  8'h00;      memory[25503] <=  8'h00;      memory[25504] <=  8'h00;      memory[25505] <=  8'h00;      memory[25506] <=  8'h00;      memory[25507] <=  8'h00;      memory[25508] <=  8'h00;      memory[25509] <=  8'h00;      memory[25510] <=  8'h00;      memory[25511] <=  8'h00;      memory[25512] <=  8'h00;      memory[25513] <=  8'h00;      memory[25514] <=  8'h00;      memory[25515] <=  8'h00;      memory[25516] <=  8'h00;      memory[25517] <=  8'h00;      memory[25518] <=  8'h00;      memory[25519] <=  8'h00;      memory[25520] <=  8'h00;      memory[25521] <=  8'h00;      memory[25522] <=  8'h00;      memory[25523] <=  8'h00;      memory[25524] <=  8'h00;      memory[25525] <=  8'h00;      memory[25526] <=  8'h00;      memory[25527] <=  8'h00;      memory[25528] <=  8'h00;      memory[25529] <=  8'h00;      memory[25530] <=  8'h00;      memory[25531] <=  8'h00;      memory[25532] <=  8'h00;      memory[25533] <=  8'h00;      memory[25534] <=  8'h00;      memory[25535] <=  8'h00;      memory[25536] <=  8'h00;      memory[25537] <=  8'h00;      memory[25538] <=  8'h00;      memory[25539] <=  8'h00;      memory[25540] <=  8'h00;      memory[25541] <=  8'h00;      memory[25542] <=  8'h00;      memory[25543] <=  8'h00;      memory[25544] <=  8'h00;      memory[25545] <=  8'h00;      memory[25546] <=  8'h00;      memory[25547] <=  8'h00;      memory[25548] <=  8'h00;      memory[25549] <=  8'h00;      memory[25550] <=  8'h00;      memory[25551] <=  8'h00;      memory[25552] <=  8'h00;      memory[25553] <=  8'h00;      memory[25554] <=  8'h00;      memory[25555] <=  8'h00;      memory[25556] <=  8'h00;      memory[25557] <=  8'h00;      memory[25558] <=  8'h00;      memory[25559] <=  8'h00;      memory[25560] <=  8'h00;      memory[25561] <=  8'h00;      memory[25562] <=  8'h00;      memory[25563] <=  8'h00;      memory[25564] <=  8'h00;      memory[25565] <=  8'h00;      memory[25566] <=  8'h00;      memory[25567] <=  8'h00;      memory[25568] <=  8'h00;      memory[25569] <=  8'h00;      memory[25570] <=  8'h00;      memory[25571] <=  8'h00;      memory[25572] <=  8'h00;      memory[25573] <=  8'h00;      memory[25574] <=  8'h00;      memory[25575] <=  8'h00;      memory[25576] <=  8'h00;      memory[25577] <=  8'h00;      memory[25578] <=  8'h00;      memory[25579] <=  8'h00;      memory[25580] <=  8'h00;      memory[25581] <=  8'h00;      memory[25582] <=  8'h00;      memory[25583] <=  8'h00;      memory[25584] <=  8'h00;      memory[25585] <=  8'h00;      memory[25586] <=  8'h00;      memory[25587] <=  8'h00;      memory[25588] <=  8'h00;      memory[25589] <=  8'h00;      memory[25590] <=  8'h00;      memory[25591] <=  8'h00;      memory[25592] <=  8'h00;      memory[25593] <=  8'h00;      memory[25594] <=  8'h00;      memory[25595] <=  8'h00;      memory[25596] <=  8'h00;      memory[25597] <=  8'h00;      memory[25598] <=  8'h00;      memory[25599] <=  8'h00;      memory[25600] <=  8'h00;      memory[25601] <=  8'h00;      memory[25602] <=  8'h00;      memory[25603] <=  8'h00;      memory[25604] <=  8'h00;      memory[25605] <=  8'h00;      memory[25606] <=  8'h00;      memory[25607] <=  8'h00;      memory[25608] <=  8'h00;      memory[25609] <=  8'h00;      memory[25610] <=  8'h00;      memory[25611] <=  8'h00;      memory[25612] <=  8'h00;      memory[25613] <=  8'h00;      memory[25614] <=  8'h00;      memory[25615] <=  8'h00;      memory[25616] <=  8'h00;      memory[25617] <=  8'h00;      memory[25618] <=  8'h00;      memory[25619] <=  8'h00;      memory[25620] <=  8'h00;      memory[25621] <=  8'h00;      memory[25622] <=  8'h00;      memory[25623] <=  8'h00;      memory[25624] <=  8'h00;      memory[25625] <=  8'h00;      memory[25626] <=  8'h00;      memory[25627] <=  8'h00;      memory[25628] <=  8'h00;      memory[25629] <=  8'h00;      memory[25630] <=  8'h00;      memory[25631] <=  8'h00;      memory[25632] <=  8'h00;      memory[25633] <=  8'h00;      memory[25634] <=  8'h00;      memory[25635] <=  8'h00;      memory[25636] <=  8'h00;      memory[25637] <=  8'h00;      memory[25638] <=  8'h00;      memory[25639] <=  8'h00;      memory[25640] <=  8'h00;      memory[25641] <=  8'h00;      memory[25642] <=  8'h00;      memory[25643] <=  8'h00;      memory[25644] <=  8'h00;      memory[25645] <=  8'h00;      memory[25646] <=  8'h00;      memory[25647] <=  8'h00;      memory[25648] <=  8'h00;      memory[25649] <=  8'h00;      memory[25650] <=  8'h00;      memory[25651] <=  8'h00;      memory[25652] <=  8'h00;      memory[25653] <=  8'h00;      memory[25654] <=  8'h00;      memory[25655] <=  8'h00;      memory[25656] <=  8'h00;      memory[25657] <=  8'h00;      memory[25658] <=  8'h00;      memory[25659] <=  8'h00;      memory[25660] <=  8'h00;      memory[25661] <=  8'h00;      memory[25662] <=  8'h00;      memory[25663] <=  8'h00;      memory[25664] <=  8'h00;      memory[25665] <=  8'h00;      memory[25666] <=  8'h00;      memory[25667] <=  8'h00;      memory[25668] <=  8'h00;      memory[25669] <=  8'h00;      memory[25670] <=  8'h00;      memory[25671] <=  8'h00;      memory[25672] <=  8'h00;      memory[25673] <=  8'h00;      memory[25674] <=  8'h00;      memory[25675] <=  8'h00;      memory[25676] <=  8'h00;      memory[25677] <=  8'h00;      memory[25678] <=  8'h00;      memory[25679] <=  8'h00;      memory[25680] <=  8'h00;      memory[25681] <=  8'h00;      memory[25682] <=  8'h00;      memory[25683] <=  8'h00;      memory[25684] <=  8'h00;      memory[25685] <=  8'h00;      memory[25686] <=  8'h00;      memory[25687] <=  8'h00;      memory[25688] <=  8'h00;      memory[25689] <=  8'h00;      memory[25690] <=  8'h00;      memory[25691] <=  8'h00;      memory[25692] <=  8'h00;      memory[25693] <=  8'h00;      memory[25694] <=  8'h00;      memory[25695] <=  8'h00;      memory[25696] <=  8'h00;      memory[25697] <=  8'h00;      memory[25698] <=  8'h00;      memory[25699] <=  8'h00;      memory[25700] <=  8'h00;      memory[25701] <=  8'h00;      memory[25702] <=  8'h00;      memory[25703] <=  8'h00;      memory[25704] <=  8'h00;      memory[25705] <=  8'h00;      memory[25706] <=  8'h00;      memory[25707] <=  8'h00;      memory[25708] <=  8'h00;      memory[25709] <=  8'h00;      memory[25710] <=  8'h00;      memory[25711] <=  8'h00;      memory[25712] <=  8'h00;      memory[25713] <=  8'h00;      memory[25714] <=  8'h00;      memory[25715] <=  8'h00;      memory[25716] <=  8'h00;      memory[25717] <=  8'h00;      memory[25718] <=  8'h00;      memory[25719] <=  8'h00;      memory[25720] <=  8'h00;      memory[25721] <=  8'h00;      memory[25722] <=  8'h00;      memory[25723] <=  8'h00;      memory[25724] <=  8'h00;      memory[25725] <=  8'h00;      memory[25726] <=  8'h00;      memory[25727] <=  8'h00;      memory[25728] <=  8'h00;      memory[25729] <=  8'h00;      memory[25730] <=  8'h00;      memory[25731] <=  8'h00;      memory[25732] <=  8'h00;      memory[25733] <=  8'h00;      memory[25734] <=  8'h00;      memory[25735] <=  8'h00;      memory[25736] <=  8'h00;      memory[25737] <=  8'h00;      memory[25738] <=  8'h00;      memory[25739] <=  8'h00;      memory[25740] <=  8'h00;      memory[25741] <=  8'h00;      memory[25742] <=  8'h00;      memory[25743] <=  8'h00;      memory[25744] <=  8'h00;      memory[25745] <=  8'h00;      memory[25746] <=  8'h00;      memory[25747] <=  8'h00;      memory[25748] <=  8'h00;      memory[25749] <=  8'h00;      memory[25750] <=  8'h00;      memory[25751] <=  8'h00;      memory[25752] <=  8'h00;      memory[25753] <=  8'h00;      memory[25754] <=  8'h00;      memory[25755] <=  8'h00;      memory[25756] <=  8'h00;      memory[25757] <=  8'h00;      memory[25758] <=  8'h00;      memory[25759] <=  8'h00;      memory[25760] <=  8'h00;      memory[25761] <=  8'h00;      memory[25762] <=  8'h00;      memory[25763] <=  8'h00;      memory[25764] <=  8'h00;      memory[25765] <=  8'h00;      memory[25766] <=  8'h00;      memory[25767] <=  8'h00;      memory[25768] <=  8'h00;      memory[25769] <=  8'h00;      memory[25770] <=  8'h00;      memory[25771] <=  8'h00;      memory[25772] <=  8'h00;      memory[25773] <=  8'h00;      memory[25774] <=  8'h00;      memory[25775] <=  8'h00;      memory[25776] <=  8'h00;      memory[25777] <=  8'h00;      memory[25778] <=  8'h00;      memory[25779] <=  8'h00;      memory[25780] <=  8'h00;      memory[25781] <=  8'h00;      memory[25782] <=  8'h00;      memory[25783] <=  8'h00;      memory[25784] <=  8'h00;      memory[25785] <=  8'h00;      memory[25786] <=  8'h00;      memory[25787] <=  8'h00;      memory[25788] <=  8'h00;      memory[25789] <=  8'h00;      memory[25790] <=  8'h00;      memory[25791] <=  8'h00;      memory[25792] <=  8'h00;      memory[25793] <=  8'h00;      memory[25794] <=  8'h00;      memory[25795] <=  8'h00;      memory[25796] <=  8'h00;      memory[25797] <=  8'h00;      memory[25798] <=  8'h00;      memory[25799] <=  8'h00;      memory[25800] <=  8'h00;      memory[25801] <=  8'h00;      memory[25802] <=  8'h00;      memory[25803] <=  8'h00;      memory[25804] <=  8'h00;      memory[25805] <=  8'h00;      memory[25806] <=  8'h00;      memory[25807] <=  8'h00;      memory[25808] <=  8'h00;      memory[25809] <=  8'h00;      memory[25810] <=  8'h00;      memory[25811] <=  8'h00;      memory[25812] <=  8'h00;      memory[25813] <=  8'h00;      memory[25814] <=  8'h00;      memory[25815] <=  8'h00;      memory[25816] <=  8'h00;      memory[25817] <=  8'h00;      memory[25818] <=  8'h00;      memory[25819] <=  8'h00;      memory[25820] <=  8'h00;      memory[25821] <=  8'h00;      memory[25822] <=  8'h00;      memory[25823] <=  8'h00;      memory[25824] <=  8'h00;      memory[25825] <=  8'h00;      memory[25826] <=  8'h00;      memory[25827] <=  8'h00;      memory[25828] <=  8'h00;      memory[25829] <=  8'h00;      memory[25830] <=  8'h00;      memory[25831] <=  8'h00;      memory[25832] <=  8'h00;      memory[25833] <=  8'h00;      memory[25834] <=  8'h00;      memory[25835] <=  8'h00;      memory[25836] <=  8'h00;      memory[25837] <=  8'h00;      memory[25838] <=  8'h00;      memory[25839] <=  8'h00;      memory[25840] <=  8'h00;      memory[25841] <=  8'h00;      memory[25842] <=  8'h00;      memory[25843] <=  8'h00;      memory[25844] <=  8'h00;      memory[25845] <=  8'h00;      memory[25846] <=  8'h00;      memory[25847] <=  8'h00;      memory[25848] <=  8'h00;      memory[25849] <=  8'h00;      memory[25850] <=  8'h00;      memory[25851] <=  8'h00;      memory[25852] <=  8'h00;      memory[25853] <=  8'h00;      memory[25854] <=  8'h00;      memory[25855] <=  8'h00;      memory[25856] <=  8'h00;      memory[25857] <=  8'h00;      memory[25858] <=  8'h00;      memory[25859] <=  8'h00;      memory[25860] <=  8'h00;      memory[25861] <=  8'h00;      memory[25862] <=  8'h00;      memory[25863] <=  8'h00;      memory[25864] <=  8'h00;      memory[25865] <=  8'h00;      memory[25866] <=  8'h00;      memory[25867] <=  8'h00;      memory[25868] <=  8'h00;      memory[25869] <=  8'h00;      memory[25870] <=  8'h00;      memory[25871] <=  8'h00;      memory[25872] <=  8'h00;      memory[25873] <=  8'h00;      memory[25874] <=  8'h00;      memory[25875] <=  8'h00;      memory[25876] <=  8'h00;      memory[25877] <=  8'h00;      memory[25878] <=  8'h00;      memory[25879] <=  8'h00;      memory[25880] <=  8'h00;      memory[25881] <=  8'h00;      memory[25882] <=  8'h00;      memory[25883] <=  8'h00;      memory[25884] <=  8'h00;      memory[25885] <=  8'h00;      memory[25886] <=  8'h00;      memory[25887] <=  8'h00;      memory[25888] <=  8'h00;      memory[25889] <=  8'h00;      memory[25890] <=  8'h00;      memory[25891] <=  8'h00;      memory[25892] <=  8'h00;      memory[25893] <=  8'h00;      memory[25894] <=  8'h00;      memory[25895] <=  8'h00;      memory[25896] <=  8'h00;      memory[25897] <=  8'h00;      memory[25898] <=  8'h00;      memory[25899] <=  8'h00;      memory[25900] <=  8'h00;      memory[25901] <=  8'h00;      memory[25902] <=  8'h00;      memory[25903] <=  8'h00;      memory[25904] <=  8'h00;      memory[25905] <=  8'h00;      memory[25906] <=  8'h00;      memory[25907] <=  8'h00;      memory[25908] <=  8'h00;      memory[25909] <=  8'h00;      memory[25910] <=  8'h00;      memory[25911] <=  8'h00;      memory[25912] <=  8'h00;      memory[25913] <=  8'h00;      memory[25914] <=  8'h00;      memory[25915] <=  8'h00;      memory[25916] <=  8'h00;      memory[25917] <=  8'h00;      memory[25918] <=  8'h00;      memory[25919] <=  8'h00;      memory[25920] <=  8'h00;      memory[25921] <=  8'h00;      memory[25922] <=  8'h00;      memory[25923] <=  8'h00;      memory[25924] <=  8'h00;      memory[25925] <=  8'h00;      memory[25926] <=  8'h00;      memory[25927] <=  8'h00;      memory[25928] <=  8'h00;      memory[25929] <=  8'h00;      memory[25930] <=  8'h00;      memory[25931] <=  8'h00;      memory[25932] <=  8'h00;      memory[25933] <=  8'h00;      memory[25934] <=  8'h00;      memory[25935] <=  8'h00;      memory[25936] <=  8'h00;      memory[25937] <=  8'h00;      memory[25938] <=  8'h00;      memory[25939] <=  8'h00;      memory[25940] <=  8'h00;      memory[25941] <=  8'h00;      memory[25942] <=  8'h00;      memory[25943] <=  8'h00;      memory[25944] <=  8'h00;      memory[25945] <=  8'h00;      memory[25946] <=  8'h00;      memory[25947] <=  8'h00;      memory[25948] <=  8'h00;      memory[25949] <=  8'h00;      memory[25950] <=  8'h00;      memory[25951] <=  8'h00;      memory[25952] <=  8'h00;      memory[25953] <=  8'h00;      memory[25954] <=  8'h00;      memory[25955] <=  8'h00;      memory[25956] <=  8'h00;      memory[25957] <=  8'h00;      memory[25958] <=  8'h00;      memory[25959] <=  8'h00;      memory[25960] <=  8'h00;      memory[25961] <=  8'h00;      memory[25962] <=  8'h00;      memory[25963] <=  8'h00;      memory[25964] <=  8'h00;      memory[25965] <=  8'h00;      memory[25966] <=  8'h00;      memory[25967] <=  8'h00;      memory[25968] <=  8'h00;      memory[25969] <=  8'h00;      memory[25970] <=  8'h00;      memory[25971] <=  8'h00;      memory[25972] <=  8'h00;      memory[25973] <=  8'h00;      memory[25974] <=  8'h00;      memory[25975] <=  8'h00;      memory[25976] <=  8'h00;      memory[25977] <=  8'h00;      memory[25978] <=  8'h00;      memory[25979] <=  8'h00;      memory[25980] <=  8'h00;      memory[25981] <=  8'h00;      memory[25982] <=  8'h00;      memory[25983] <=  8'h00;      memory[25984] <=  8'h00;      memory[25985] <=  8'h00;      memory[25986] <=  8'h00;      memory[25987] <=  8'h00;      memory[25988] <=  8'h00;      memory[25989] <=  8'h00;      memory[25990] <=  8'h00;      memory[25991] <=  8'h00;      memory[25992] <=  8'h00;      memory[25993] <=  8'h00;      memory[25994] <=  8'h00;      memory[25995] <=  8'h00;      memory[25996] <=  8'h00;      memory[25997] <=  8'h00;      memory[25998] <=  8'h00;      memory[25999] <=  8'h00;      memory[26000] <=  8'h00;      memory[26001] <=  8'h00;      memory[26002] <=  8'h00;      memory[26003] <=  8'h00;      memory[26004] <=  8'h00;      memory[26005] <=  8'h00;      memory[26006] <=  8'h00;      memory[26007] <=  8'h00;      memory[26008] <=  8'h00;      memory[26009] <=  8'h00;      memory[26010] <=  8'h00;      memory[26011] <=  8'h00;      memory[26012] <=  8'h00;      memory[26013] <=  8'h00;      memory[26014] <=  8'h00;      memory[26015] <=  8'h00;      memory[26016] <=  8'h00;      memory[26017] <=  8'h00;      memory[26018] <=  8'h00;      memory[26019] <=  8'h00;      memory[26020] <=  8'h00;      memory[26021] <=  8'h00;      memory[26022] <=  8'h00;      memory[26023] <=  8'h00;      memory[26024] <=  8'h00;      memory[26025] <=  8'h00;      memory[26026] <=  8'h00;      memory[26027] <=  8'h00;      memory[26028] <=  8'h00;      memory[26029] <=  8'h00;      memory[26030] <=  8'h00;      memory[26031] <=  8'h00;      memory[26032] <=  8'h00;      memory[26033] <=  8'h00;      memory[26034] <=  8'h00;      memory[26035] <=  8'h00;      memory[26036] <=  8'h00;      memory[26037] <=  8'h00;      memory[26038] <=  8'h00;      memory[26039] <=  8'h00;      memory[26040] <=  8'h00;      memory[26041] <=  8'h00;      memory[26042] <=  8'h00;      memory[26043] <=  8'h00;      memory[26044] <=  8'h00;      memory[26045] <=  8'h00;      memory[26046] <=  8'h00;      memory[26047] <=  8'h00;      memory[26048] <=  8'h00;      memory[26049] <=  8'h00;      memory[26050] <=  8'h00;      memory[26051] <=  8'h00;      memory[26052] <=  8'h00;      memory[26053] <=  8'h00;      memory[26054] <=  8'h00;      memory[26055] <=  8'h00;      memory[26056] <=  8'h00;      memory[26057] <=  8'h00;      memory[26058] <=  8'h00;      memory[26059] <=  8'h00;      memory[26060] <=  8'h00;      memory[26061] <=  8'h00;      memory[26062] <=  8'h00;      memory[26063] <=  8'h00;      memory[26064] <=  8'h00;      memory[26065] <=  8'h00;      memory[26066] <=  8'h00;      memory[26067] <=  8'h00;      memory[26068] <=  8'h00;      memory[26069] <=  8'h00;      memory[26070] <=  8'h00;      memory[26071] <=  8'h00;      memory[26072] <=  8'h00;      memory[26073] <=  8'h00;      memory[26074] <=  8'h00;      memory[26075] <=  8'h00;      memory[26076] <=  8'h00;      memory[26077] <=  8'h00;      memory[26078] <=  8'h00;      memory[26079] <=  8'h00;      memory[26080] <=  8'h00;      memory[26081] <=  8'h00;      memory[26082] <=  8'h00;      memory[26083] <=  8'h00;      memory[26084] <=  8'h00;      memory[26085] <=  8'h00;      memory[26086] <=  8'h00;      memory[26087] <=  8'h00;      memory[26088] <=  8'h00;      memory[26089] <=  8'h00;      memory[26090] <=  8'h00;      memory[26091] <=  8'h00;      memory[26092] <=  8'h00;      memory[26093] <=  8'h00;      memory[26094] <=  8'h00;      memory[26095] <=  8'h00;      memory[26096] <=  8'h00;      memory[26097] <=  8'h00;      memory[26098] <=  8'h00;      memory[26099] <=  8'h00;      memory[26100] <=  8'h00;      memory[26101] <=  8'h00;      memory[26102] <=  8'h00;      memory[26103] <=  8'h00;      memory[26104] <=  8'h00;      memory[26105] <=  8'h00;      memory[26106] <=  8'h00;      memory[26107] <=  8'h00;      memory[26108] <=  8'h00;      memory[26109] <=  8'h00;      memory[26110] <=  8'h00;      memory[26111] <=  8'h00;      memory[26112] <=  8'h00;      memory[26113] <=  8'h00;      memory[26114] <=  8'h00;      memory[26115] <=  8'h00;      memory[26116] <=  8'h00;      memory[26117] <=  8'h00;      memory[26118] <=  8'h00;      memory[26119] <=  8'h00;      memory[26120] <=  8'h00;      memory[26121] <=  8'h00;      memory[26122] <=  8'h00;      memory[26123] <=  8'h00;      memory[26124] <=  8'h00;      memory[26125] <=  8'h00;      memory[26126] <=  8'h00;      memory[26127] <=  8'h00;      memory[26128] <=  8'h00;      memory[26129] <=  8'h00;      memory[26130] <=  8'h00;      memory[26131] <=  8'h00;      memory[26132] <=  8'h00;      memory[26133] <=  8'h00;      memory[26134] <=  8'h00;      memory[26135] <=  8'h00;      memory[26136] <=  8'h00;      memory[26137] <=  8'h00;      memory[26138] <=  8'h00;      memory[26139] <=  8'h00;      memory[26140] <=  8'h00;      memory[26141] <=  8'h00;      memory[26142] <=  8'h00;      memory[26143] <=  8'h00;      memory[26144] <=  8'h00;      memory[26145] <=  8'h00;      memory[26146] <=  8'h00;      memory[26147] <=  8'h00;      memory[26148] <=  8'h00;      memory[26149] <=  8'h00;      memory[26150] <=  8'h00;      memory[26151] <=  8'h00;      memory[26152] <=  8'h00;      memory[26153] <=  8'h00;      memory[26154] <=  8'h00;      memory[26155] <=  8'h00;      memory[26156] <=  8'h00;      memory[26157] <=  8'h00;      memory[26158] <=  8'h00;      memory[26159] <=  8'h00;      memory[26160] <=  8'h00;      memory[26161] <=  8'h00;      memory[26162] <=  8'h00;      memory[26163] <=  8'h00;      memory[26164] <=  8'h00;      memory[26165] <=  8'h00;      memory[26166] <=  8'h00;      memory[26167] <=  8'h00;      memory[26168] <=  8'h00;      memory[26169] <=  8'h00;      memory[26170] <=  8'h00;      memory[26171] <=  8'h00;      memory[26172] <=  8'h00;      memory[26173] <=  8'h00;      memory[26174] <=  8'h00;      memory[26175] <=  8'h00;      memory[26176] <=  8'h00;      memory[26177] <=  8'h00;      memory[26178] <=  8'h00;      memory[26179] <=  8'h00;      memory[26180] <=  8'h00;      memory[26181] <=  8'h00;      memory[26182] <=  8'h00;      memory[26183] <=  8'h00;      memory[26184] <=  8'h00;      memory[26185] <=  8'h00;      memory[26186] <=  8'h00;      memory[26187] <=  8'h00;      memory[26188] <=  8'h00;      memory[26189] <=  8'h00;      memory[26190] <=  8'h00;      memory[26191] <=  8'h00;      memory[26192] <=  8'h00;      memory[26193] <=  8'h00;      memory[26194] <=  8'h00;      memory[26195] <=  8'h00;      memory[26196] <=  8'h00;      memory[26197] <=  8'h00;      memory[26198] <=  8'h00;      memory[26199] <=  8'h00;      memory[26200] <=  8'h00;      memory[26201] <=  8'h00;      memory[26202] <=  8'h00;      memory[26203] <=  8'h00;      memory[26204] <=  8'h00;      memory[26205] <=  8'h00;      memory[26206] <=  8'h00;      memory[26207] <=  8'h00;      memory[26208] <=  8'h00;      memory[26209] <=  8'h00;      memory[26210] <=  8'h00;      memory[26211] <=  8'h00;      memory[26212] <=  8'h00;      memory[26213] <=  8'h00;      memory[26214] <=  8'h00;      memory[26215] <=  8'h00;      memory[26216] <=  8'h00;      memory[26217] <=  8'h00;      memory[26218] <=  8'h00;      memory[26219] <=  8'h00;      memory[26220] <=  8'h00;      memory[26221] <=  8'h00;      memory[26222] <=  8'h00;      memory[26223] <=  8'h00;      memory[26224] <=  8'h00;      memory[26225] <=  8'h00;      memory[26226] <=  8'h00;      memory[26227] <=  8'h00;      memory[26228] <=  8'h00;      memory[26229] <=  8'h00;      memory[26230] <=  8'h00;      memory[26231] <=  8'h00;      memory[26232] <=  8'h00;      memory[26233] <=  8'h00;      memory[26234] <=  8'h00;      memory[26235] <=  8'h00;      memory[26236] <=  8'h00;      memory[26237] <=  8'h00;      memory[26238] <=  8'h00;      memory[26239] <=  8'h00;      memory[26240] <=  8'h00;      memory[26241] <=  8'h00;      memory[26242] <=  8'h00;      memory[26243] <=  8'h00;      memory[26244] <=  8'h00;      memory[26245] <=  8'h00;      memory[26246] <=  8'h00;      memory[26247] <=  8'h00;      memory[26248] <=  8'h00;      memory[26249] <=  8'h00;      memory[26250] <=  8'h00;      memory[26251] <=  8'h00;      memory[26252] <=  8'h00;      memory[26253] <=  8'h00;      memory[26254] <=  8'h00;      memory[26255] <=  8'h00;      memory[26256] <=  8'h00;      memory[26257] <=  8'h00;      memory[26258] <=  8'h00;      memory[26259] <=  8'h00;      memory[26260] <=  8'h00;      memory[26261] <=  8'h00;      memory[26262] <=  8'h00;      memory[26263] <=  8'h00;      memory[26264] <=  8'h00;      memory[26265] <=  8'h00;      memory[26266] <=  8'h00;      memory[26267] <=  8'h00;      memory[26268] <=  8'h00;      memory[26269] <=  8'h00;      memory[26270] <=  8'h00;      memory[26271] <=  8'h00;      memory[26272] <=  8'h00;      memory[26273] <=  8'h00;      memory[26274] <=  8'h00;      memory[26275] <=  8'h00;      memory[26276] <=  8'h00;      memory[26277] <=  8'h00;      memory[26278] <=  8'h00;      memory[26279] <=  8'h00;      memory[26280] <=  8'h00;      memory[26281] <=  8'h00;      memory[26282] <=  8'h00;      memory[26283] <=  8'h00;      memory[26284] <=  8'h00;      memory[26285] <=  8'h00;      memory[26286] <=  8'h00;      memory[26287] <=  8'h00;      memory[26288] <=  8'h00;      memory[26289] <=  8'h00;      memory[26290] <=  8'h00;      memory[26291] <=  8'h00;      memory[26292] <=  8'h00;      memory[26293] <=  8'h00;      memory[26294] <=  8'h00;      memory[26295] <=  8'h00;      memory[26296] <=  8'h00;      memory[26297] <=  8'h00;      memory[26298] <=  8'h00;      memory[26299] <=  8'h00;      memory[26300] <=  8'h00;      memory[26301] <=  8'h00;      memory[26302] <=  8'h00;      memory[26303] <=  8'h00;      memory[26304] <=  8'h00;      memory[26305] <=  8'h00;      memory[26306] <=  8'h00;      memory[26307] <=  8'h00;      memory[26308] <=  8'h00;      memory[26309] <=  8'h00;      memory[26310] <=  8'h00;      memory[26311] <=  8'h00;      memory[26312] <=  8'h00;      memory[26313] <=  8'h00;      memory[26314] <=  8'h00;      memory[26315] <=  8'h00;      memory[26316] <=  8'h00;      memory[26317] <=  8'h00;      memory[26318] <=  8'h00;      memory[26319] <=  8'h00;      memory[26320] <=  8'h00;      memory[26321] <=  8'h00;      memory[26322] <=  8'h00;      memory[26323] <=  8'h00;      memory[26324] <=  8'h00;      memory[26325] <=  8'h00;      memory[26326] <=  8'h00;      memory[26327] <=  8'h00;      memory[26328] <=  8'h00;      memory[26329] <=  8'h00;      memory[26330] <=  8'h00;      memory[26331] <=  8'h00;      memory[26332] <=  8'h00;      memory[26333] <=  8'h00;      memory[26334] <=  8'h00;      memory[26335] <=  8'h00;      memory[26336] <=  8'h00;      memory[26337] <=  8'h00;      memory[26338] <=  8'h00;      memory[26339] <=  8'h00;      memory[26340] <=  8'h00;      memory[26341] <=  8'h00;      memory[26342] <=  8'h00;      memory[26343] <=  8'h00;      memory[26344] <=  8'h00;      memory[26345] <=  8'h00;      memory[26346] <=  8'h00;      memory[26347] <=  8'h00;      memory[26348] <=  8'h00;      memory[26349] <=  8'h00;      memory[26350] <=  8'h00;      memory[26351] <=  8'h00;      memory[26352] <=  8'h00;      memory[26353] <=  8'h00;      memory[26354] <=  8'h00;      memory[26355] <=  8'h00;      memory[26356] <=  8'h00;      memory[26357] <=  8'h00;      memory[26358] <=  8'h00;      memory[26359] <=  8'h00;      memory[26360] <=  8'h00;      memory[26361] <=  8'h00;      memory[26362] <=  8'h00;      memory[26363] <=  8'h00;      memory[26364] <=  8'h00;      memory[26365] <=  8'h00;      memory[26366] <=  8'h00;      memory[26367] <=  8'h00;      memory[26368] <=  8'h00;      memory[26369] <=  8'h00;      memory[26370] <=  8'h00;      memory[26371] <=  8'h00;      memory[26372] <=  8'h00;      memory[26373] <=  8'h00;      memory[26374] <=  8'h00;      memory[26375] <=  8'h00;      memory[26376] <=  8'h00;      memory[26377] <=  8'h00;      memory[26378] <=  8'h00;      memory[26379] <=  8'h00;      memory[26380] <=  8'h00;      memory[26381] <=  8'h00;      memory[26382] <=  8'h00;      memory[26383] <=  8'h00;      memory[26384] <=  8'h00;      memory[26385] <=  8'h00;      memory[26386] <=  8'h00;      memory[26387] <=  8'h00;      memory[26388] <=  8'h00;      memory[26389] <=  8'h00;      memory[26390] <=  8'h00;      memory[26391] <=  8'h00;      memory[26392] <=  8'h00;      memory[26393] <=  8'h00;      memory[26394] <=  8'h00;      memory[26395] <=  8'h00;      memory[26396] <=  8'h00;      memory[26397] <=  8'h00;      memory[26398] <=  8'h00;      memory[26399] <=  8'h00;      memory[26400] <=  8'h00;      memory[26401] <=  8'h00;      memory[26402] <=  8'h00;      memory[26403] <=  8'h00;      memory[26404] <=  8'h00;      memory[26405] <=  8'h00;      memory[26406] <=  8'h00;      memory[26407] <=  8'h00;      memory[26408] <=  8'h00;      memory[26409] <=  8'h00;      memory[26410] <=  8'h00;      memory[26411] <=  8'h00;      memory[26412] <=  8'h00;      memory[26413] <=  8'h00;      memory[26414] <=  8'h00;      memory[26415] <=  8'h00;      memory[26416] <=  8'h00;      memory[26417] <=  8'h00;      memory[26418] <=  8'h00;      memory[26419] <=  8'h00;      memory[26420] <=  8'h00;      memory[26421] <=  8'h00;      memory[26422] <=  8'h00;      memory[26423] <=  8'h00;      memory[26424] <=  8'h00;      memory[26425] <=  8'h00;      memory[26426] <=  8'h00;      memory[26427] <=  8'h00;      memory[26428] <=  8'h00;      memory[26429] <=  8'h00;      memory[26430] <=  8'h00;      memory[26431] <=  8'h00;      memory[26432] <=  8'h00;      memory[26433] <=  8'h00;      memory[26434] <=  8'h00;      memory[26435] <=  8'h00;      memory[26436] <=  8'h00;      memory[26437] <=  8'h00;      memory[26438] <=  8'h00;      memory[26439] <=  8'h00;      memory[26440] <=  8'h00;      memory[26441] <=  8'h00;      memory[26442] <=  8'h00;      memory[26443] <=  8'h00;      memory[26444] <=  8'h00;      memory[26445] <=  8'h00;      memory[26446] <=  8'h00;      memory[26447] <=  8'h00;      memory[26448] <=  8'h00;      memory[26449] <=  8'h00;      memory[26450] <=  8'h00;      memory[26451] <=  8'h00;      memory[26452] <=  8'h00;      memory[26453] <=  8'h00;      memory[26454] <=  8'h00;      memory[26455] <=  8'h00;      memory[26456] <=  8'h00;      memory[26457] <=  8'h00;      memory[26458] <=  8'h00;      memory[26459] <=  8'h00;      memory[26460] <=  8'h00;      memory[26461] <=  8'h00;      memory[26462] <=  8'h00;      memory[26463] <=  8'h00;      memory[26464] <=  8'h00;      memory[26465] <=  8'h00;      memory[26466] <=  8'h00;      memory[26467] <=  8'h00;      memory[26468] <=  8'h00;      memory[26469] <=  8'h00;      memory[26470] <=  8'h00;      memory[26471] <=  8'h00;      memory[26472] <=  8'h00;      memory[26473] <=  8'h00;      memory[26474] <=  8'h00;      memory[26475] <=  8'h00;      memory[26476] <=  8'h00;      memory[26477] <=  8'h00;      memory[26478] <=  8'h00;      memory[26479] <=  8'h00;      memory[26480] <=  8'h00;      memory[26481] <=  8'h00;      memory[26482] <=  8'h00;      memory[26483] <=  8'h00;      memory[26484] <=  8'h00;      memory[26485] <=  8'h00;      memory[26486] <=  8'h00;      memory[26487] <=  8'h00;      memory[26488] <=  8'h00;      memory[26489] <=  8'h00;      memory[26490] <=  8'h00;      memory[26491] <=  8'h00;      memory[26492] <=  8'h00;      memory[26493] <=  8'h00;      memory[26494] <=  8'h00;      memory[26495] <=  8'h00;      memory[26496] <=  8'h00;      memory[26497] <=  8'h00;      memory[26498] <=  8'h00;      memory[26499] <=  8'h00;      memory[26500] <=  8'h00;      memory[26501] <=  8'h00;      memory[26502] <=  8'h00;      memory[26503] <=  8'h00;      memory[26504] <=  8'h00;      memory[26505] <=  8'h00;      memory[26506] <=  8'h00;      memory[26507] <=  8'h00;      memory[26508] <=  8'h00;      memory[26509] <=  8'h00;      memory[26510] <=  8'h00;      memory[26511] <=  8'h00;      memory[26512] <=  8'h00;      memory[26513] <=  8'h00;      memory[26514] <=  8'h00;      memory[26515] <=  8'h00;      memory[26516] <=  8'h00;      memory[26517] <=  8'h00;      memory[26518] <=  8'h00;      memory[26519] <=  8'h00;      memory[26520] <=  8'h00;      memory[26521] <=  8'h00;      memory[26522] <=  8'h00;      memory[26523] <=  8'h00;      memory[26524] <=  8'h00;      memory[26525] <=  8'h00;      memory[26526] <=  8'h00;      memory[26527] <=  8'h00;      memory[26528] <=  8'h00;      memory[26529] <=  8'h00;      memory[26530] <=  8'h00;      memory[26531] <=  8'h00;      memory[26532] <=  8'h00;      memory[26533] <=  8'h00;      memory[26534] <=  8'h00;      memory[26535] <=  8'h00;      memory[26536] <=  8'h00;      memory[26537] <=  8'h00;      memory[26538] <=  8'h00;      memory[26539] <=  8'h00;      memory[26540] <=  8'h00;      memory[26541] <=  8'h00;      memory[26542] <=  8'h00;      memory[26543] <=  8'h00;      memory[26544] <=  8'h00;      memory[26545] <=  8'h00;      memory[26546] <=  8'h00;      memory[26547] <=  8'h00;      memory[26548] <=  8'h00;      memory[26549] <=  8'h00;      memory[26550] <=  8'h00;      memory[26551] <=  8'h00;      memory[26552] <=  8'h00;      memory[26553] <=  8'h00;      memory[26554] <=  8'h00;      memory[26555] <=  8'h00;      memory[26556] <=  8'h00;      memory[26557] <=  8'h00;      memory[26558] <=  8'h00;      memory[26559] <=  8'h00;      memory[26560] <=  8'h00;      memory[26561] <=  8'h00;      memory[26562] <=  8'h00;      memory[26563] <=  8'h00;      memory[26564] <=  8'h00;      memory[26565] <=  8'h00;      memory[26566] <=  8'h00;      memory[26567] <=  8'h00;      memory[26568] <=  8'h00;      memory[26569] <=  8'h00;      memory[26570] <=  8'h00;      memory[26571] <=  8'h00;      memory[26572] <=  8'h00;      memory[26573] <=  8'h00;      memory[26574] <=  8'h00;      memory[26575] <=  8'h00;      memory[26576] <=  8'h00;      memory[26577] <=  8'h00;      memory[26578] <=  8'h00;      memory[26579] <=  8'h00;      memory[26580] <=  8'h00;      memory[26581] <=  8'h00;      memory[26582] <=  8'h00;      memory[26583] <=  8'h00;      memory[26584] <=  8'h00;      memory[26585] <=  8'h00;      memory[26586] <=  8'h00;      memory[26587] <=  8'h00;      memory[26588] <=  8'h00;      memory[26589] <=  8'h00;      memory[26590] <=  8'h00;      memory[26591] <=  8'h00;      memory[26592] <=  8'h00;      memory[26593] <=  8'h00;      memory[26594] <=  8'h00;      memory[26595] <=  8'h00;      memory[26596] <=  8'h00;      memory[26597] <=  8'h00;      memory[26598] <=  8'h00;      memory[26599] <=  8'h00;      memory[26600] <=  8'h00;      memory[26601] <=  8'h00;      memory[26602] <=  8'h00;      memory[26603] <=  8'h00;      memory[26604] <=  8'h00;      memory[26605] <=  8'h00;      memory[26606] <=  8'h00;      memory[26607] <=  8'h00;      memory[26608] <=  8'h00;      memory[26609] <=  8'h00;      memory[26610] <=  8'h00;      memory[26611] <=  8'h00;      memory[26612] <=  8'h00;      memory[26613] <=  8'h00;      memory[26614] <=  8'h00;      memory[26615] <=  8'h00;      memory[26616] <=  8'h00;      memory[26617] <=  8'h00;      memory[26618] <=  8'h00;      memory[26619] <=  8'h00;      memory[26620] <=  8'h00;      memory[26621] <=  8'h00;      memory[26622] <=  8'h00;      memory[26623] <=  8'h00;      memory[26624] <=  8'h00;      memory[26625] <=  8'h00;      memory[26626] <=  8'h00;      memory[26627] <=  8'h00;      memory[26628] <=  8'h00;      memory[26629] <=  8'h00;      memory[26630] <=  8'h00;      memory[26631] <=  8'h00;      memory[26632] <=  8'h00;      memory[26633] <=  8'h00;      memory[26634] <=  8'h00;      memory[26635] <=  8'h00;      memory[26636] <=  8'h00;      memory[26637] <=  8'h00;      memory[26638] <=  8'h00;      memory[26639] <=  8'h00;      memory[26640] <=  8'h00;      memory[26641] <=  8'h00;      memory[26642] <=  8'h00;      memory[26643] <=  8'h00;      memory[26644] <=  8'h00;      memory[26645] <=  8'h00;      memory[26646] <=  8'h00;      memory[26647] <=  8'h00;      memory[26648] <=  8'h00;      memory[26649] <=  8'h00;      memory[26650] <=  8'h00;      memory[26651] <=  8'h00;      memory[26652] <=  8'h00;      memory[26653] <=  8'h00;      memory[26654] <=  8'h00;      memory[26655] <=  8'h00;      memory[26656] <=  8'h00;      memory[26657] <=  8'h00;      memory[26658] <=  8'h00;      memory[26659] <=  8'h00;      memory[26660] <=  8'h00;      memory[26661] <=  8'h00;      memory[26662] <=  8'h00;      memory[26663] <=  8'h00;      memory[26664] <=  8'h00;      memory[26665] <=  8'h00;      memory[26666] <=  8'h00;      memory[26667] <=  8'h00;      memory[26668] <=  8'h00;      memory[26669] <=  8'h00;      memory[26670] <=  8'h00;      memory[26671] <=  8'h00;      memory[26672] <=  8'h00;      memory[26673] <=  8'h00;      memory[26674] <=  8'h00;      memory[26675] <=  8'h00;      memory[26676] <=  8'h00;      memory[26677] <=  8'h00;      memory[26678] <=  8'h00;      memory[26679] <=  8'h00;      memory[26680] <=  8'h00;      memory[26681] <=  8'h00;      memory[26682] <=  8'h00;      memory[26683] <=  8'h00;      memory[26684] <=  8'h00;      memory[26685] <=  8'h00;      memory[26686] <=  8'h00;      memory[26687] <=  8'h00;      memory[26688] <=  8'h00;      memory[26689] <=  8'h00;      memory[26690] <=  8'h00;      memory[26691] <=  8'h00;      memory[26692] <=  8'h00;      memory[26693] <=  8'h00;      memory[26694] <=  8'h00;      memory[26695] <=  8'h00;      memory[26696] <=  8'h00;      memory[26697] <=  8'h00;      memory[26698] <=  8'h00;      memory[26699] <=  8'h00;      memory[26700] <=  8'h00;      memory[26701] <=  8'h00;      memory[26702] <=  8'h00;      memory[26703] <=  8'h00;      memory[26704] <=  8'h00;      memory[26705] <=  8'h00;      memory[26706] <=  8'h00;      memory[26707] <=  8'h00;      memory[26708] <=  8'h00;      memory[26709] <=  8'h00;      memory[26710] <=  8'h00;      memory[26711] <=  8'h00;      memory[26712] <=  8'h00;      memory[26713] <=  8'h00;      memory[26714] <=  8'h00;      memory[26715] <=  8'h00;      memory[26716] <=  8'h00;      memory[26717] <=  8'h00;      memory[26718] <=  8'h00;      memory[26719] <=  8'h00;      memory[26720] <=  8'h00;      memory[26721] <=  8'h00;      memory[26722] <=  8'h00;      memory[26723] <=  8'h00;      memory[26724] <=  8'h00;      memory[26725] <=  8'h00;      memory[26726] <=  8'h00;      memory[26727] <=  8'h00;      memory[26728] <=  8'h00;      memory[26729] <=  8'h00;      memory[26730] <=  8'h00;      memory[26731] <=  8'h00;      memory[26732] <=  8'h00;      memory[26733] <=  8'h00;      memory[26734] <=  8'h00;      memory[26735] <=  8'h00;      memory[26736] <=  8'h00;      memory[26737] <=  8'h00;      memory[26738] <=  8'h00;      memory[26739] <=  8'h00;      memory[26740] <=  8'h00;      memory[26741] <=  8'h00;      memory[26742] <=  8'h00;      memory[26743] <=  8'h00;      memory[26744] <=  8'h00;      memory[26745] <=  8'h00;      memory[26746] <=  8'h00;      memory[26747] <=  8'h00;      memory[26748] <=  8'h00;      memory[26749] <=  8'h00;      memory[26750] <=  8'h00;      memory[26751] <=  8'h00;      memory[26752] <=  8'h00;      memory[26753] <=  8'h00;      memory[26754] <=  8'h00;      memory[26755] <=  8'h00;      memory[26756] <=  8'h00;      memory[26757] <=  8'h00;      memory[26758] <=  8'h00;      memory[26759] <=  8'h00;      memory[26760] <=  8'h00;      memory[26761] <=  8'h00;      memory[26762] <=  8'h00;      memory[26763] <=  8'h00;      memory[26764] <=  8'h00;      memory[26765] <=  8'h00;      memory[26766] <=  8'h00;      memory[26767] <=  8'h00;      memory[26768] <=  8'h00;      memory[26769] <=  8'h00;      memory[26770] <=  8'h00;      memory[26771] <=  8'h00;      memory[26772] <=  8'h00;      memory[26773] <=  8'h00;      memory[26774] <=  8'h00;      memory[26775] <=  8'h00;      memory[26776] <=  8'h00;      memory[26777] <=  8'h00;      memory[26778] <=  8'h00;      memory[26779] <=  8'h00;      memory[26780] <=  8'h00;      memory[26781] <=  8'h00;      memory[26782] <=  8'h00;      memory[26783] <=  8'h00;      memory[26784] <=  8'h00;      memory[26785] <=  8'h00;      memory[26786] <=  8'h00;      memory[26787] <=  8'h00;      memory[26788] <=  8'h00;      memory[26789] <=  8'h00;      memory[26790] <=  8'h00;      memory[26791] <=  8'h00;      memory[26792] <=  8'h00;      memory[26793] <=  8'h00;      memory[26794] <=  8'h00;      memory[26795] <=  8'h00;      memory[26796] <=  8'h00;      memory[26797] <=  8'h00;      memory[26798] <=  8'h00;      memory[26799] <=  8'h00;      memory[26800] <=  8'h00;      memory[26801] <=  8'h00;      memory[26802] <=  8'h00;      memory[26803] <=  8'h00;      memory[26804] <=  8'h00;      memory[26805] <=  8'h00;      memory[26806] <=  8'h00;      memory[26807] <=  8'h00;      memory[26808] <=  8'h00;      memory[26809] <=  8'h00;      memory[26810] <=  8'h00;      memory[26811] <=  8'h00;      memory[26812] <=  8'h00;      memory[26813] <=  8'h00;      memory[26814] <=  8'h00;      memory[26815] <=  8'h00;      memory[26816] <=  8'h00;      memory[26817] <=  8'h00;      memory[26818] <=  8'h00;      memory[26819] <=  8'h00;      memory[26820] <=  8'h00;      memory[26821] <=  8'h00;      memory[26822] <=  8'h00;      memory[26823] <=  8'h00;      memory[26824] <=  8'h00;      memory[26825] <=  8'h00;      memory[26826] <=  8'h00;      memory[26827] <=  8'h00;      memory[26828] <=  8'h00;      memory[26829] <=  8'h00;      memory[26830] <=  8'h00;      memory[26831] <=  8'h00;      memory[26832] <=  8'h00;      memory[26833] <=  8'h00;      memory[26834] <=  8'h00;      memory[26835] <=  8'h00;      memory[26836] <=  8'h00;      memory[26837] <=  8'h00;      memory[26838] <=  8'h00;      memory[26839] <=  8'h00;      memory[26840] <=  8'h00;      memory[26841] <=  8'h00;      memory[26842] <=  8'h00;      memory[26843] <=  8'h00;      memory[26844] <=  8'h00;      memory[26845] <=  8'h00;      memory[26846] <=  8'h00;      memory[26847] <=  8'h00;      memory[26848] <=  8'h00;      memory[26849] <=  8'h00;      memory[26850] <=  8'h00;      memory[26851] <=  8'h00;      memory[26852] <=  8'h00;      memory[26853] <=  8'h00;      memory[26854] <=  8'h00;      memory[26855] <=  8'h00;      memory[26856] <=  8'h00;      memory[26857] <=  8'h00;      memory[26858] <=  8'h00;      memory[26859] <=  8'h00;      memory[26860] <=  8'h00;      memory[26861] <=  8'h00;      memory[26862] <=  8'h00;      memory[26863] <=  8'h00;      memory[26864] <=  8'h00;      memory[26865] <=  8'h00;      memory[26866] <=  8'h00;      memory[26867] <=  8'h00;      memory[26868] <=  8'h00;      memory[26869] <=  8'h00;      memory[26870] <=  8'h00;      memory[26871] <=  8'h00;      memory[26872] <=  8'h00;      memory[26873] <=  8'h00;      memory[26874] <=  8'h00;      memory[26875] <=  8'h00;      memory[26876] <=  8'h00;      memory[26877] <=  8'h00;      memory[26878] <=  8'h00;      memory[26879] <=  8'h00;      memory[26880] <=  8'h00;      memory[26881] <=  8'h00;      memory[26882] <=  8'h00;      memory[26883] <=  8'h00;      memory[26884] <=  8'h00;      memory[26885] <=  8'h00;      memory[26886] <=  8'h00;      memory[26887] <=  8'h00;      memory[26888] <=  8'h00;      memory[26889] <=  8'h00;      memory[26890] <=  8'h00;      memory[26891] <=  8'h00;      memory[26892] <=  8'h00;      memory[26893] <=  8'h00;      memory[26894] <=  8'h00;      memory[26895] <=  8'h00;      memory[26896] <=  8'h00;      memory[26897] <=  8'h00;      memory[26898] <=  8'h00;      memory[26899] <=  8'h00;      memory[26900] <=  8'h00;      memory[26901] <=  8'h00;      memory[26902] <=  8'h00;      memory[26903] <=  8'h00;      memory[26904] <=  8'h00;      memory[26905] <=  8'h00;      memory[26906] <=  8'h00;      memory[26907] <=  8'h00;      memory[26908] <=  8'h00;      memory[26909] <=  8'h00;      memory[26910] <=  8'h00;      memory[26911] <=  8'h00;      memory[26912] <=  8'h00;      memory[26913] <=  8'h00;      memory[26914] <=  8'h00;      memory[26915] <=  8'h00;      memory[26916] <=  8'h00;      memory[26917] <=  8'h00;      memory[26918] <=  8'h00;      memory[26919] <=  8'h00;      memory[26920] <=  8'h00;      memory[26921] <=  8'h00;      memory[26922] <=  8'h00;      memory[26923] <=  8'h00;      memory[26924] <=  8'h00;      memory[26925] <=  8'h00;      memory[26926] <=  8'h00;      memory[26927] <=  8'h00;      memory[26928] <=  8'h00;      memory[26929] <=  8'h00;      memory[26930] <=  8'h00;      memory[26931] <=  8'h00;      memory[26932] <=  8'h00;      memory[26933] <=  8'h00;      memory[26934] <=  8'h00;      memory[26935] <=  8'h00;      memory[26936] <=  8'h00;      memory[26937] <=  8'h00;      memory[26938] <=  8'h00;      memory[26939] <=  8'h00;      memory[26940] <=  8'h00;      memory[26941] <=  8'h00;      memory[26942] <=  8'h00;      memory[26943] <=  8'h00;      memory[26944] <=  8'h00;      memory[26945] <=  8'h00;      memory[26946] <=  8'h00;      memory[26947] <=  8'h00;      memory[26948] <=  8'h00;      memory[26949] <=  8'h00;      memory[26950] <=  8'h00;      memory[26951] <=  8'h00;      memory[26952] <=  8'h00;      memory[26953] <=  8'h00;      memory[26954] <=  8'h00;      memory[26955] <=  8'h00;      memory[26956] <=  8'h00;      memory[26957] <=  8'h00;      memory[26958] <=  8'h00;      memory[26959] <=  8'h00;      memory[26960] <=  8'h00;      memory[26961] <=  8'h00;      memory[26962] <=  8'h00;      memory[26963] <=  8'h00;      memory[26964] <=  8'h00;      memory[26965] <=  8'h00;      memory[26966] <=  8'h00;      memory[26967] <=  8'h00;      memory[26968] <=  8'h00;      memory[26969] <=  8'h00;      memory[26970] <=  8'h00;      memory[26971] <=  8'h00;      memory[26972] <=  8'h00;      memory[26973] <=  8'h00;      memory[26974] <=  8'h00;      memory[26975] <=  8'h00;      memory[26976] <=  8'h00;      memory[26977] <=  8'h00;      memory[26978] <=  8'h00;      memory[26979] <=  8'h00;      memory[26980] <=  8'h00;      memory[26981] <=  8'h00;      memory[26982] <=  8'h00;      memory[26983] <=  8'h00;      memory[26984] <=  8'h00;      memory[26985] <=  8'h00;      memory[26986] <=  8'h00;      memory[26987] <=  8'h00;      memory[26988] <=  8'h00;      memory[26989] <=  8'h00;      memory[26990] <=  8'h00;      memory[26991] <=  8'h00;      memory[26992] <=  8'h00;      memory[26993] <=  8'h00;      memory[26994] <=  8'h00;      memory[26995] <=  8'h00;      memory[26996] <=  8'h00;      memory[26997] <=  8'h00;      memory[26998] <=  8'h00;      memory[26999] <=  8'h00;      memory[27000] <=  8'h00;      memory[27001] <=  8'h00;      memory[27002] <=  8'h00;      memory[27003] <=  8'h00;      memory[27004] <=  8'h00;      memory[27005] <=  8'h00;      memory[27006] <=  8'h00;      memory[27007] <=  8'h00;      memory[27008] <=  8'h00;      memory[27009] <=  8'h00;      memory[27010] <=  8'h00;      memory[27011] <=  8'h00;      memory[27012] <=  8'h00;      memory[27013] <=  8'h00;      memory[27014] <=  8'h00;      memory[27015] <=  8'h00;      memory[27016] <=  8'h00;      memory[27017] <=  8'h00;      memory[27018] <=  8'h00;      memory[27019] <=  8'h00;      memory[27020] <=  8'h00;      memory[27021] <=  8'h00;      memory[27022] <=  8'h00;      memory[27023] <=  8'h00;      memory[27024] <=  8'h00;      memory[27025] <=  8'h00;      memory[27026] <=  8'h00;      memory[27027] <=  8'h00;      memory[27028] <=  8'h00;      memory[27029] <=  8'h00;      memory[27030] <=  8'h00;      memory[27031] <=  8'h00;      memory[27032] <=  8'h00;      memory[27033] <=  8'h00;      memory[27034] <=  8'h00;      memory[27035] <=  8'h00;      memory[27036] <=  8'h00;      memory[27037] <=  8'h00;      memory[27038] <=  8'h00;      memory[27039] <=  8'h00;      memory[27040] <=  8'h00;      memory[27041] <=  8'h00;      memory[27042] <=  8'h00;      memory[27043] <=  8'h00;      memory[27044] <=  8'h00;      memory[27045] <=  8'h00;      memory[27046] <=  8'h00;      memory[27047] <=  8'h00;      memory[27048] <=  8'h00;      memory[27049] <=  8'h00;      memory[27050] <=  8'h00;      memory[27051] <=  8'h00;      memory[27052] <=  8'h00;      memory[27053] <=  8'h00;      memory[27054] <=  8'h00;      memory[27055] <=  8'h00;      memory[27056] <=  8'h00;      memory[27057] <=  8'h00;      memory[27058] <=  8'h00;      memory[27059] <=  8'h00;      memory[27060] <=  8'h00;      memory[27061] <=  8'h00;      memory[27062] <=  8'h00;      memory[27063] <=  8'h00;      memory[27064] <=  8'h00;      memory[27065] <=  8'h00;      memory[27066] <=  8'h00;      memory[27067] <=  8'h00;      memory[27068] <=  8'h00;      memory[27069] <=  8'h00;      memory[27070] <=  8'h00;      memory[27071] <=  8'h00;      memory[27072] <=  8'h00;      memory[27073] <=  8'h00;      memory[27074] <=  8'h00;      memory[27075] <=  8'h00;      memory[27076] <=  8'h00;      memory[27077] <=  8'h00;      memory[27078] <=  8'h00;      memory[27079] <=  8'h00;      memory[27080] <=  8'h00;      memory[27081] <=  8'h00;      memory[27082] <=  8'h00;      memory[27083] <=  8'h00;      memory[27084] <=  8'h00;      memory[27085] <=  8'h00;      memory[27086] <=  8'h00;      memory[27087] <=  8'h00;      memory[27088] <=  8'h00;      memory[27089] <=  8'h00;      memory[27090] <=  8'h00;      memory[27091] <=  8'h00;      memory[27092] <=  8'h00;      memory[27093] <=  8'h00;      memory[27094] <=  8'h00;      memory[27095] <=  8'h00;      memory[27096] <=  8'h00;      memory[27097] <=  8'h00;      memory[27098] <=  8'h00;      memory[27099] <=  8'h00;      memory[27100] <=  8'h00;      memory[27101] <=  8'h00;      memory[27102] <=  8'h00;      memory[27103] <=  8'h00;      memory[27104] <=  8'h00;      memory[27105] <=  8'h00;      memory[27106] <=  8'h00;      memory[27107] <=  8'h00;      memory[27108] <=  8'h00;      memory[27109] <=  8'h00;      memory[27110] <=  8'h00;      memory[27111] <=  8'h00;      memory[27112] <=  8'h00;      memory[27113] <=  8'h00;      memory[27114] <=  8'h00;      memory[27115] <=  8'h00;      memory[27116] <=  8'h00;      memory[27117] <=  8'h00;      memory[27118] <=  8'h00;      memory[27119] <=  8'h00;      memory[27120] <=  8'h00;      memory[27121] <=  8'h00;      memory[27122] <=  8'h00;      memory[27123] <=  8'h00;      memory[27124] <=  8'h00;      memory[27125] <=  8'h00;      memory[27126] <=  8'h00;      memory[27127] <=  8'h00;      memory[27128] <=  8'h00;      memory[27129] <=  8'h00;      memory[27130] <=  8'h00;      memory[27131] <=  8'h00;      memory[27132] <=  8'h00;      memory[27133] <=  8'h00;      memory[27134] <=  8'h00;      memory[27135] <=  8'h00;      memory[27136] <=  8'h00;      memory[27137] <=  8'h00;      memory[27138] <=  8'h00;      memory[27139] <=  8'h00;      memory[27140] <=  8'h00;      memory[27141] <=  8'h00;      memory[27142] <=  8'h00;      memory[27143] <=  8'h00;      memory[27144] <=  8'h00;      memory[27145] <=  8'h00;      memory[27146] <=  8'h00;      memory[27147] <=  8'h00;      memory[27148] <=  8'h00;      memory[27149] <=  8'h00;      memory[27150] <=  8'h00;      memory[27151] <=  8'h00;      memory[27152] <=  8'h00;      memory[27153] <=  8'h00;      memory[27154] <=  8'h00;      memory[27155] <=  8'h00;      memory[27156] <=  8'h00;      memory[27157] <=  8'h00;      memory[27158] <=  8'h00;      memory[27159] <=  8'h00;      memory[27160] <=  8'h00;      memory[27161] <=  8'h00;      memory[27162] <=  8'h00;      memory[27163] <=  8'h00;      memory[27164] <=  8'h00;      memory[27165] <=  8'h00;      memory[27166] <=  8'h00;      memory[27167] <=  8'h00;      memory[27168] <=  8'h00;      memory[27169] <=  8'h00;      memory[27170] <=  8'h00;      memory[27171] <=  8'h00;      memory[27172] <=  8'h00;      memory[27173] <=  8'h00;      memory[27174] <=  8'h00;      memory[27175] <=  8'h00;      memory[27176] <=  8'h00;      memory[27177] <=  8'h00;      memory[27178] <=  8'h00;      memory[27179] <=  8'h00;      memory[27180] <=  8'h00;      memory[27181] <=  8'h00;      memory[27182] <=  8'h00;      memory[27183] <=  8'h00;      memory[27184] <=  8'h00;      memory[27185] <=  8'h00;      memory[27186] <=  8'h00;      memory[27187] <=  8'h00;      memory[27188] <=  8'h00;      memory[27189] <=  8'h00;      memory[27190] <=  8'h00;      memory[27191] <=  8'h00;      memory[27192] <=  8'h00;      memory[27193] <=  8'h00;      memory[27194] <=  8'h00;      memory[27195] <=  8'h00;      memory[27196] <=  8'h00;      memory[27197] <=  8'h00;      memory[27198] <=  8'h00;      memory[27199] <=  8'h00;      memory[27200] <=  8'h00;      memory[27201] <=  8'h00;      memory[27202] <=  8'h00;      memory[27203] <=  8'h00;      memory[27204] <=  8'h00;      memory[27205] <=  8'h00;      memory[27206] <=  8'h00;      memory[27207] <=  8'h00;      memory[27208] <=  8'h00;      memory[27209] <=  8'h00;      memory[27210] <=  8'h00;      memory[27211] <=  8'h00;      memory[27212] <=  8'h00;      memory[27213] <=  8'h00;      memory[27214] <=  8'h00;      memory[27215] <=  8'h00;      memory[27216] <=  8'h00;      memory[27217] <=  8'h00;      memory[27218] <=  8'h00;      memory[27219] <=  8'h00;      memory[27220] <=  8'h00;      memory[27221] <=  8'h00;      memory[27222] <=  8'h00;      memory[27223] <=  8'h00;      memory[27224] <=  8'h00;      memory[27225] <=  8'h00;      memory[27226] <=  8'h00;      memory[27227] <=  8'h00;      memory[27228] <=  8'h00;      memory[27229] <=  8'h00;      memory[27230] <=  8'h00;      memory[27231] <=  8'h00;      memory[27232] <=  8'h00;      memory[27233] <=  8'h00;      memory[27234] <=  8'h00;      memory[27235] <=  8'h00;      memory[27236] <=  8'h00;      memory[27237] <=  8'h00;      memory[27238] <=  8'h00;      memory[27239] <=  8'h00;      memory[27240] <=  8'h00;      memory[27241] <=  8'h00;      memory[27242] <=  8'h00;      memory[27243] <=  8'h00;      memory[27244] <=  8'h00;      memory[27245] <=  8'h00;      memory[27246] <=  8'h00;      memory[27247] <=  8'h00;      memory[27248] <=  8'h00;      memory[27249] <=  8'h00;      memory[27250] <=  8'h00;      memory[27251] <=  8'h00;      memory[27252] <=  8'h00;      memory[27253] <=  8'h00;      memory[27254] <=  8'h00;      memory[27255] <=  8'h00;      memory[27256] <=  8'h00;      memory[27257] <=  8'h00;      memory[27258] <=  8'h00;      memory[27259] <=  8'h00;      memory[27260] <=  8'h00;      memory[27261] <=  8'h00;      memory[27262] <=  8'h00;      memory[27263] <=  8'h00;      memory[27264] <=  8'h00;      memory[27265] <=  8'h00;      memory[27266] <=  8'h00;      memory[27267] <=  8'h00;      memory[27268] <=  8'h00;      memory[27269] <=  8'h00;      memory[27270] <=  8'h00;      memory[27271] <=  8'h00;      memory[27272] <=  8'h00;      memory[27273] <=  8'h00;      memory[27274] <=  8'h00;      memory[27275] <=  8'h00;      memory[27276] <=  8'h00;      memory[27277] <=  8'h00;      memory[27278] <=  8'h00;      memory[27279] <=  8'h00;      memory[27280] <=  8'h00;      memory[27281] <=  8'h00;      memory[27282] <=  8'h00;      memory[27283] <=  8'h00;      memory[27284] <=  8'h00;      memory[27285] <=  8'h00;      memory[27286] <=  8'h00;      memory[27287] <=  8'h00;      memory[27288] <=  8'h00;      memory[27289] <=  8'h00;      memory[27290] <=  8'h00;      memory[27291] <=  8'h00;      memory[27292] <=  8'h00;      memory[27293] <=  8'h00;      memory[27294] <=  8'h00;      memory[27295] <=  8'h00;      memory[27296] <=  8'h00;      memory[27297] <=  8'h00;      memory[27298] <=  8'h00;      memory[27299] <=  8'h00;      memory[27300] <=  8'h00;      memory[27301] <=  8'h00;      memory[27302] <=  8'h00;      memory[27303] <=  8'h00;      memory[27304] <=  8'h00;      memory[27305] <=  8'h00;      memory[27306] <=  8'h00;      memory[27307] <=  8'h00;      memory[27308] <=  8'h00;      memory[27309] <=  8'h00;      memory[27310] <=  8'h00;      memory[27311] <=  8'h00;      memory[27312] <=  8'h00;      memory[27313] <=  8'h00;      memory[27314] <=  8'h00;      memory[27315] <=  8'h00;      memory[27316] <=  8'h00;      memory[27317] <=  8'h00;      memory[27318] <=  8'h00;      memory[27319] <=  8'h00;      memory[27320] <=  8'h00;      memory[27321] <=  8'h00;      memory[27322] <=  8'h00;      memory[27323] <=  8'h00;      memory[27324] <=  8'h00;      memory[27325] <=  8'h00;      memory[27326] <=  8'h00;      memory[27327] <=  8'h00;      memory[27328] <=  8'h00;      memory[27329] <=  8'h00;      memory[27330] <=  8'h00;      memory[27331] <=  8'h00;      memory[27332] <=  8'h00;      memory[27333] <=  8'h00;      memory[27334] <=  8'h00;      memory[27335] <=  8'h00;      memory[27336] <=  8'h00;      memory[27337] <=  8'h00;      memory[27338] <=  8'h00;      memory[27339] <=  8'h00;      memory[27340] <=  8'h00;      memory[27341] <=  8'h00;      memory[27342] <=  8'h00;      memory[27343] <=  8'h00;      memory[27344] <=  8'h00;      memory[27345] <=  8'h00;      memory[27346] <=  8'h00;      memory[27347] <=  8'h00;      memory[27348] <=  8'h00;      memory[27349] <=  8'h00;      memory[27350] <=  8'h00;      memory[27351] <=  8'h00;      memory[27352] <=  8'h00;      memory[27353] <=  8'h00;      memory[27354] <=  8'h00;      memory[27355] <=  8'h00;      memory[27356] <=  8'h00;      memory[27357] <=  8'h00;      memory[27358] <=  8'h00;      memory[27359] <=  8'h00;      memory[27360] <=  8'h00;      memory[27361] <=  8'h00;      memory[27362] <=  8'h00;      memory[27363] <=  8'h00;      memory[27364] <=  8'h00;      memory[27365] <=  8'h00;      memory[27366] <=  8'h00;      memory[27367] <=  8'h00;      memory[27368] <=  8'h00;      memory[27369] <=  8'h00;      memory[27370] <=  8'h00;      memory[27371] <=  8'h00;      memory[27372] <=  8'h00;      memory[27373] <=  8'h00;      memory[27374] <=  8'h00;      memory[27375] <=  8'h00;      memory[27376] <=  8'h00;      memory[27377] <=  8'h00;      memory[27378] <=  8'h00;      memory[27379] <=  8'h00;      memory[27380] <=  8'h00;      memory[27381] <=  8'h00;      memory[27382] <=  8'h00;      memory[27383] <=  8'h00;      memory[27384] <=  8'h00;      memory[27385] <=  8'h00;      memory[27386] <=  8'h00;      memory[27387] <=  8'h00;      memory[27388] <=  8'h00;      memory[27389] <=  8'h00;      memory[27390] <=  8'h00;      memory[27391] <=  8'h00;      memory[27392] <=  8'h00;      memory[27393] <=  8'h00;      memory[27394] <=  8'h00;      memory[27395] <=  8'h00;      memory[27396] <=  8'h00;      memory[27397] <=  8'h00;      memory[27398] <=  8'h00;      memory[27399] <=  8'h00;      memory[27400] <=  8'h00;      memory[27401] <=  8'h00;      memory[27402] <=  8'h00;      memory[27403] <=  8'h00;      memory[27404] <=  8'h00;      memory[27405] <=  8'h00;      memory[27406] <=  8'h00;      memory[27407] <=  8'h00;      memory[27408] <=  8'h00;      memory[27409] <=  8'h00;      memory[27410] <=  8'h00;      memory[27411] <=  8'h00;      memory[27412] <=  8'h00;      memory[27413] <=  8'h00;      memory[27414] <=  8'h00;      memory[27415] <=  8'h00;      memory[27416] <=  8'h00;      memory[27417] <=  8'h00;      memory[27418] <=  8'h00;      memory[27419] <=  8'h00;      memory[27420] <=  8'h00;      memory[27421] <=  8'h00;      memory[27422] <=  8'h00;      memory[27423] <=  8'h00;      memory[27424] <=  8'h00;      memory[27425] <=  8'h00;      memory[27426] <=  8'h00;      memory[27427] <=  8'h00;      memory[27428] <=  8'h00;      memory[27429] <=  8'h00;      memory[27430] <=  8'h00;      memory[27431] <=  8'h00;      memory[27432] <=  8'h00;      memory[27433] <=  8'h00;      memory[27434] <=  8'h00;      memory[27435] <=  8'h00;      memory[27436] <=  8'h00;      memory[27437] <=  8'h00;      memory[27438] <=  8'h00;      memory[27439] <=  8'h00;      memory[27440] <=  8'h00;      memory[27441] <=  8'h00;      memory[27442] <=  8'h00;      memory[27443] <=  8'h00;      memory[27444] <=  8'h00;      memory[27445] <=  8'h00;      memory[27446] <=  8'h00;      memory[27447] <=  8'h00;      memory[27448] <=  8'h00;      memory[27449] <=  8'h00;      memory[27450] <=  8'h00;      memory[27451] <=  8'h00;      memory[27452] <=  8'h00;      memory[27453] <=  8'h00;      memory[27454] <=  8'h00;      memory[27455] <=  8'h00;      memory[27456] <=  8'h00;      memory[27457] <=  8'h00;      memory[27458] <=  8'h00;      memory[27459] <=  8'h00;      memory[27460] <=  8'h00;      memory[27461] <=  8'h00;      memory[27462] <=  8'h00;      memory[27463] <=  8'h00;      memory[27464] <=  8'h00;      memory[27465] <=  8'h00;      memory[27466] <=  8'h00;      memory[27467] <=  8'h00;      memory[27468] <=  8'h00;      memory[27469] <=  8'h00;      memory[27470] <=  8'h00;      memory[27471] <=  8'h00;      memory[27472] <=  8'h00;      memory[27473] <=  8'h00;      memory[27474] <=  8'h00;      memory[27475] <=  8'h00;      memory[27476] <=  8'h00;      memory[27477] <=  8'h00;      memory[27478] <=  8'h00;      memory[27479] <=  8'h00;      memory[27480] <=  8'h00;      memory[27481] <=  8'h00;      memory[27482] <=  8'h00;      memory[27483] <=  8'h00;      memory[27484] <=  8'h00;      memory[27485] <=  8'h00;      memory[27486] <=  8'h00;      memory[27487] <=  8'h00;      memory[27488] <=  8'h00;      memory[27489] <=  8'h00;      memory[27490] <=  8'h00;      memory[27491] <=  8'h00;      memory[27492] <=  8'h00;      memory[27493] <=  8'h00;      memory[27494] <=  8'h00;      memory[27495] <=  8'h00;      memory[27496] <=  8'h00;      memory[27497] <=  8'h00;      memory[27498] <=  8'h00;      memory[27499] <=  8'h00;      memory[27500] <=  8'h00;      memory[27501] <=  8'h00;      memory[27502] <=  8'h00;      memory[27503] <=  8'h00;      memory[27504] <=  8'h00;      memory[27505] <=  8'h00;      memory[27506] <=  8'h00;      memory[27507] <=  8'h00;      memory[27508] <=  8'h00;      memory[27509] <=  8'h00;      memory[27510] <=  8'h00;      memory[27511] <=  8'h00;      memory[27512] <=  8'h00;      memory[27513] <=  8'h00;      memory[27514] <=  8'h00;      memory[27515] <=  8'h00;      memory[27516] <=  8'h00;      memory[27517] <=  8'h00;      memory[27518] <=  8'h00;      memory[27519] <=  8'h00;      memory[27520] <=  8'h00;      memory[27521] <=  8'h00;      memory[27522] <=  8'h00;      memory[27523] <=  8'h00;      memory[27524] <=  8'h00;      memory[27525] <=  8'h00;      memory[27526] <=  8'h00;      memory[27527] <=  8'h00;      memory[27528] <=  8'h00;      memory[27529] <=  8'h00;      memory[27530] <=  8'h00;      memory[27531] <=  8'h00;      memory[27532] <=  8'h00;      memory[27533] <=  8'h00;      memory[27534] <=  8'h00;      memory[27535] <=  8'h00;      memory[27536] <=  8'h00;      memory[27537] <=  8'h00;      memory[27538] <=  8'h00;      memory[27539] <=  8'h00;      memory[27540] <=  8'h00;      memory[27541] <=  8'h00;      memory[27542] <=  8'h00;      memory[27543] <=  8'h00;      memory[27544] <=  8'h00;      memory[27545] <=  8'h00;      memory[27546] <=  8'h00;      memory[27547] <=  8'h00;      memory[27548] <=  8'h00;      memory[27549] <=  8'h00;      memory[27550] <=  8'h00;      memory[27551] <=  8'h00;      memory[27552] <=  8'h00;      memory[27553] <=  8'h00;      memory[27554] <=  8'h00;      memory[27555] <=  8'h00;      memory[27556] <=  8'h00;      memory[27557] <=  8'h00;      memory[27558] <=  8'h00;      memory[27559] <=  8'h00;      memory[27560] <=  8'h00;      memory[27561] <=  8'h00;      memory[27562] <=  8'h00;      memory[27563] <=  8'h00;      memory[27564] <=  8'h00;      memory[27565] <=  8'h00;      memory[27566] <=  8'h00;      memory[27567] <=  8'h00;      memory[27568] <=  8'h00;      memory[27569] <=  8'h00;      memory[27570] <=  8'h00;      memory[27571] <=  8'h00;      memory[27572] <=  8'h00;      memory[27573] <=  8'h00;      memory[27574] <=  8'h00;      memory[27575] <=  8'h00;      memory[27576] <=  8'h00;      memory[27577] <=  8'h00;      memory[27578] <=  8'h00;      memory[27579] <=  8'h00;      memory[27580] <=  8'h00;      memory[27581] <=  8'h00;      memory[27582] <=  8'h00;      memory[27583] <=  8'h00;      memory[27584] <=  8'h00;      memory[27585] <=  8'h00;      memory[27586] <=  8'h00;      memory[27587] <=  8'h00;      memory[27588] <=  8'h00;      memory[27589] <=  8'h00;      memory[27590] <=  8'h00;      memory[27591] <=  8'h00;      memory[27592] <=  8'h00;      memory[27593] <=  8'h00;      memory[27594] <=  8'h00;      memory[27595] <=  8'h00;      memory[27596] <=  8'h00;      memory[27597] <=  8'h00;      memory[27598] <=  8'h00;      memory[27599] <=  8'h00;      memory[27600] <=  8'h00;      memory[27601] <=  8'h00;      memory[27602] <=  8'h00;      memory[27603] <=  8'h00;      memory[27604] <=  8'h00;      memory[27605] <=  8'h00;      memory[27606] <=  8'h00;      memory[27607] <=  8'h00;      memory[27608] <=  8'h00;      memory[27609] <=  8'h00;      memory[27610] <=  8'h00;      memory[27611] <=  8'h00;      memory[27612] <=  8'h00;      memory[27613] <=  8'h00;      memory[27614] <=  8'h00;      memory[27615] <=  8'h00;      memory[27616] <=  8'h00;      memory[27617] <=  8'h00;      memory[27618] <=  8'h00;      memory[27619] <=  8'h00;      memory[27620] <=  8'h00;      memory[27621] <=  8'h00;      memory[27622] <=  8'h00;      memory[27623] <=  8'h00;      memory[27624] <=  8'h00;      memory[27625] <=  8'h00;      memory[27626] <=  8'h00;      memory[27627] <=  8'h00;      memory[27628] <=  8'h00;      memory[27629] <=  8'h00;      memory[27630] <=  8'h00;      memory[27631] <=  8'h00;      memory[27632] <=  8'h00;      memory[27633] <=  8'h00;      memory[27634] <=  8'h00;      memory[27635] <=  8'h00;      memory[27636] <=  8'h00;      memory[27637] <=  8'h00;      memory[27638] <=  8'h00;      memory[27639] <=  8'h00;      memory[27640] <=  8'h00;      memory[27641] <=  8'h00;      memory[27642] <=  8'h00;      memory[27643] <=  8'h00;      memory[27644] <=  8'h00;      memory[27645] <=  8'h00;      memory[27646] <=  8'h00;      memory[27647] <=  8'h00;      memory[27648] <=  8'h00;      memory[27649] <=  8'h00;      memory[27650] <=  8'h00;      memory[27651] <=  8'h00;      memory[27652] <=  8'h00;      memory[27653] <=  8'h00;      memory[27654] <=  8'h00;      memory[27655] <=  8'h00;      memory[27656] <=  8'h00;      memory[27657] <=  8'h00;      memory[27658] <=  8'h00;      memory[27659] <=  8'h00;      memory[27660] <=  8'h00;      memory[27661] <=  8'h00;      memory[27662] <=  8'h00;      memory[27663] <=  8'h00;      memory[27664] <=  8'h00;      memory[27665] <=  8'h00;      memory[27666] <=  8'h00;      memory[27667] <=  8'h00;      memory[27668] <=  8'h00;      memory[27669] <=  8'h00;      memory[27670] <=  8'h00;      memory[27671] <=  8'h00;      memory[27672] <=  8'h00;      memory[27673] <=  8'h00;      memory[27674] <=  8'h00;      memory[27675] <=  8'h00;      memory[27676] <=  8'h00;      memory[27677] <=  8'h00;      memory[27678] <=  8'h00;      memory[27679] <=  8'h00;      memory[27680] <=  8'h00;      memory[27681] <=  8'h00;      memory[27682] <=  8'h00;      memory[27683] <=  8'h00;      memory[27684] <=  8'h00;      memory[27685] <=  8'h00;      memory[27686] <=  8'h00;      memory[27687] <=  8'h00;      memory[27688] <=  8'h00;      memory[27689] <=  8'h00;      memory[27690] <=  8'h00;      memory[27691] <=  8'h00;      memory[27692] <=  8'h00;      memory[27693] <=  8'h00;      memory[27694] <=  8'h00;      memory[27695] <=  8'h00;      memory[27696] <=  8'h00;      memory[27697] <=  8'h00;      memory[27698] <=  8'h00;      memory[27699] <=  8'h00;      memory[27700] <=  8'h00;      memory[27701] <=  8'h00;      memory[27702] <=  8'h00;      memory[27703] <=  8'h00;      memory[27704] <=  8'h00;      memory[27705] <=  8'h00;      memory[27706] <=  8'h00;      memory[27707] <=  8'h00;      memory[27708] <=  8'h00;      memory[27709] <=  8'h00;      memory[27710] <=  8'h00;      memory[27711] <=  8'h00;      memory[27712] <=  8'h00;      memory[27713] <=  8'h00;      memory[27714] <=  8'h00;      memory[27715] <=  8'h00;      memory[27716] <=  8'h00;      memory[27717] <=  8'h00;      memory[27718] <=  8'h00;      memory[27719] <=  8'h00;      memory[27720] <=  8'h00;      memory[27721] <=  8'h00;      memory[27722] <=  8'h00;      memory[27723] <=  8'h00;      memory[27724] <=  8'h00;      memory[27725] <=  8'h00;      memory[27726] <=  8'h00;      memory[27727] <=  8'h00;      memory[27728] <=  8'h00;      memory[27729] <=  8'h00;      memory[27730] <=  8'h00;      memory[27731] <=  8'h00;      memory[27732] <=  8'h00;      memory[27733] <=  8'h00;      memory[27734] <=  8'h00;      memory[27735] <=  8'h00;      memory[27736] <=  8'h00;      memory[27737] <=  8'h00;      memory[27738] <=  8'h00;      memory[27739] <=  8'h00;      memory[27740] <=  8'h00;      memory[27741] <=  8'h00;      memory[27742] <=  8'h00;      memory[27743] <=  8'h00;      memory[27744] <=  8'h00;      memory[27745] <=  8'h00;      memory[27746] <=  8'h00;      memory[27747] <=  8'h00;      memory[27748] <=  8'h00;      memory[27749] <=  8'h00;      memory[27750] <=  8'h00;      memory[27751] <=  8'h00;      memory[27752] <=  8'h00;      memory[27753] <=  8'h00;      memory[27754] <=  8'h00;      memory[27755] <=  8'h00;      memory[27756] <=  8'h00;      memory[27757] <=  8'h00;      memory[27758] <=  8'h00;      memory[27759] <=  8'h00;      memory[27760] <=  8'h00;      memory[27761] <=  8'h00;      memory[27762] <=  8'h00;      memory[27763] <=  8'h00;      memory[27764] <=  8'h00;      memory[27765] <=  8'h00;      memory[27766] <=  8'h00;      memory[27767] <=  8'h00;      memory[27768] <=  8'h00;      memory[27769] <=  8'h00;      memory[27770] <=  8'h00;      memory[27771] <=  8'h00;      memory[27772] <=  8'h00;      memory[27773] <=  8'h00;      memory[27774] <=  8'h00;      memory[27775] <=  8'h00;      memory[27776] <=  8'h00;      memory[27777] <=  8'h00;      memory[27778] <=  8'h00;      memory[27779] <=  8'h00;      memory[27780] <=  8'h00;      memory[27781] <=  8'h00;      memory[27782] <=  8'h00;      memory[27783] <=  8'h00;      memory[27784] <=  8'h00;      memory[27785] <=  8'h00;      memory[27786] <=  8'h00;      memory[27787] <=  8'h00;      memory[27788] <=  8'h00;      memory[27789] <=  8'h00;      memory[27790] <=  8'h00;      memory[27791] <=  8'h00;      memory[27792] <=  8'h00;      memory[27793] <=  8'h00;      memory[27794] <=  8'h00;      memory[27795] <=  8'h00;      memory[27796] <=  8'h00;      memory[27797] <=  8'h00;      memory[27798] <=  8'h00;      memory[27799] <=  8'h00;      memory[27800] <=  8'h00;      memory[27801] <=  8'h00;      memory[27802] <=  8'h00;      memory[27803] <=  8'h00;      memory[27804] <=  8'h00;      memory[27805] <=  8'h00;      memory[27806] <=  8'h00;      memory[27807] <=  8'h00;      memory[27808] <=  8'h00;      memory[27809] <=  8'h00;      memory[27810] <=  8'h00;      memory[27811] <=  8'h00;      memory[27812] <=  8'h00;      memory[27813] <=  8'h00;      memory[27814] <=  8'h00;      memory[27815] <=  8'h00;      memory[27816] <=  8'h00;      memory[27817] <=  8'h00;      memory[27818] <=  8'h00;      memory[27819] <=  8'h00;      memory[27820] <=  8'h00;      memory[27821] <=  8'h00;      memory[27822] <=  8'h00;      memory[27823] <=  8'h00;      memory[27824] <=  8'h00;      memory[27825] <=  8'h00;      memory[27826] <=  8'h00;      memory[27827] <=  8'h00;      memory[27828] <=  8'h00;      memory[27829] <=  8'h00;      memory[27830] <=  8'h00;      memory[27831] <=  8'h00;      memory[27832] <=  8'h00;      memory[27833] <=  8'h00;      memory[27834] <=  8'h00;      memory[27835] <=  8'h00;      memory[27836] <=  8'h00;      memory[27837] <=  8'h00;      memory[27838] <=  8'h00;      memory[27839] <=  8'h00;      memory[27840] <=  8'h00;      memory[27841] <=  8'h00;      memory[27842] <=  8'h00;      memory[27843] <=  8'h00;      memory[27844] <=  8'h00;      memory[27845] <=  8'h00;      memory[27846] <=  8'h00;      memory[27847] <=  8'h00;      memory[27848] <=  8'h00;      memory[27849] <=  8'h00;      memory[27850] <=  8'h00;      memory[27851] <=  8'h00;      memory[27852] <=  8'h00;      memory[27853] <=  8'h00;      memory[27854] <=  8'h00;      memory[27855] <=  8'h00;      memory[27856] <=  8'h00;      memory[27857] <=  8'h00;      memory[27858] <=  8'h00;      memory[27859] <=  8'h00;      memory[27860] <=  8'h00;      memory[27861] <=  8'h00;      memory[27862] <=  8'h00;      memory[27863] <=  8'h00;      memory[27864] <=  8'h00;      memory[27865] <=  8'h00;      memory[27866] <=  8'h00;      memory[27867] <=  8'h00;      memory[27868] <=  8'h00;      memory[27869] <=  8'h00;      memory[27870] <=  8'h00;      memory[27871] <=  8'h00;      memory[27872] <=  8'h00;      memory[27873] <=  8'h00;      memory[27874] <=  8'h00;      memory[27875] <=  8'h00;      memory[27876] <=  8'h00;      memory[27877] <=  8'h00;      memory[27878] <=  8'h00;      memory[27879] <=  8'h00;      memory[27880] <=  8'h00;      memory[27881] <=  8'h00;      memory[27882] <=  8'h00;      memory[27883] <=  8'h00;      memory[27884] <=  8'h00;      memory[27885] <=  8'h00;      memory[27886] <=  8'h00;      memory[27887] <=  8'h00;      memory[27888] <=  8'h00;      memory[27889] <=  8'h00;      memory[27890] <=  8'h00;      memory[27891] <=  8'h00;      memory[27892] <=  8'h00;      memory[27893] <=  8'h00;      memory[27894] <=  8'h00;      memory[27895] <=  8'h00;      memory[27896] <=  8'h00;      memory[27897] <=  8'h00;      memory[27898] <=  8'h00;      memory[27899] <=  8'h00;      memory[27900] <=  8'h00;      memory[27901] <=  8'h00;      memory[27902] <=  8'h00;      memory[27903] <=  8'h00;      memory[27904] <=  8'h00;      memory[27905] <=  8'h00;      memory[27906] <=  8'h00;      memory[27907] <=  8'h00;      memory[27908] <=  8'h00;      memory[27909] <=  8'h00;      memory[27910] <=  8'h00;      memory[27911] <=  8'h00;      memory[27912] <=  8'h00;      memory[27913] <=  8'h00;      memory[27914] <=  8'h00;      memory[27915] <=  8'h00;      memory[27916] <=  8'h00;      memory[27917] <=  8'h00;      memory[27918] <=  8'h00;      memory[27919] <=  8'h00;      memory[27920] <=  8'h00;      memory[27921] <=  8'h00;      memory[27922] <=  8'h00;      memory[27923] <=  8'h00;      memory[27924] <=  8'h00;      memory[27925] <=  8'h00;      memory[27926] <=  8'h00;      memory[27927] <=  8'h00;      memory[27928] <=  8'h00;      memory[27929] <=  8'h00;      memory[27930] <=  8'h00;      memory[27931] <=  8'h00;      memory[27932] <=  8'h00;      memory[27933] <=  8'h00;      memory[27934] <=  8'h00;      memory[27935] <=  8'h00;      memory[27936] <=  8'h00;      memory[27937] <=  8'h00;      memory[27938] <=  8'h00;      memory[27939] <=  8'h00;      memory[27940] <=  8'h00;      memory[27941] <=  8'h00;      memory[27942] <=  8'h00;      memory[27943] <=  8'h00;      memory[27944] <=  8'h00;      memory[27945] <=  8'h00;      memory[27946] <=  8'h00;      memory[27947] <=  8'h00;      memory[27948] <=  8'h00;      memory[27949] <=  8'h00;      memory[27950] <=  8'h00;      memory[27951] <=  8'h00;      memory[27952] <=  8'h00;      memory[27953] <=  8'h00;      memory[27954] <=  8'h00;      memory[27955] <=  8'h00;      memory[27956] <=  8'h00;      memory[27957] <=  8'h00;      memory[27958] <=  8'h00;      memory[27959] <=  8'h00;      memory[27960] <=  8'h00;      memory[27961] <=  8'h00;      memory[27962] <=  8'h00;      memory[27963] <=  8'h00;      memory[27964] <=  8'h00;      memory[27965] <=  8'h00;      memory[27966] <=  8'h00;      memory[27967] <=  8'h00;      memory[27968] <=  8'h00;      memory[27969] <=  8'h00;      memory[27970] <=  8'h00;      memory[27971] <=  8'h00;      memory[27972] <=  8'h00;      memory[27973] <=  8'h00;      memory[27974] <=  8'h00;      memory[27975] <=  8'h00;      memory[27976] <=  8'h00;      memory[27977] <=  8'h00;      memory[27978] <=  8'h00;      memory[27979] <=  8'h00;      memory[27980] <=  8'h00;      memory[27981] <=  8'h00;      memory[27982] <=  8'h00;      memory[27983] <=  8'h00;      memory[27984] <=  8'h00;      memory[27985] <=  8'h00;      memory[27986] <=  8'h00;      memory[27987] <=  8'h00;      memory[27988] <=  8'h00;      memory[27989] <=  8'h00;      memory[27990] <=  8'h00;      memory[27991] <=  8'h00;      memory[27992] <=  8'h00;      memory[27993] <=  8'h00;      memory[27994] <=  8'h00;      memory[27995] <=  8'h00;      memory[27996] <=  8'h00;      memory[27997] <=  8'h00;      memory[27998] <=  8'h00;      memory[27999] <=  8'h00;      memory[28000] <=  8'h00;      memory[28001] <=  8'h00;      memory[28002] <=  8'h00;      memory[28003] <=  8'h00;      memory[28004] <=  8'h00;      memory[28005] <=  8'h00;      memory[28006] <=  8'h00;      memory[28007] <=  8'h00;      memory[28008] <=  8'h00;      memory[28009] <=  8'h00;      memory[28010] <=  8'h00;      memory[28011] <=  8'h00;      memory[28012] <=  8'h00;      memory[28013] <=  8'h00;      memory[28014] <=  8'h00;      memory[28015] <=  8'h00;      memory[28016] <=  8'h00;      memory[28017] <=  8'h00;      memory[28018] <=  8'h00;      memory[28019] <=  8'h00;      memory[28020] <=  8'h00;      memory[28021] <=  8'h00;      memory[28022] <=  8'h00;      memory[28023] <=  8'h00;      memory[28024] <=  8'h00;      memory[28025] <=  8'h00;      memory[28026] <=  8'h00;      memory[28027] <=  8'h00;      memory[28028] <=  8'h00;      memory[28029] <=  8'h00;      memory[28030] <=  8'h00;      memory[28031] <=  8'h00;      memory[28032] <=  8'h00;      memory[28033] <=  8'h00;      memory[28034] <=  8'h00;      memory[28035] <=  8'h00;      memory[28036] <=  8'h00;      memory[28037] <=  8'h00;      memory[28038] <=  8'h00;      memory[28039] <=  8'h00;      memory[28040] <=  8'h00;      memory[28041] <=  8'h00;      memory[28042] <=  8'h00;      memory[28043] <=  8'h00;      memory[28044] <=  8'h00;      memory[28045] <=  8'h00;      memory[28046] <=  8'h00;      memory[28047] <=  8'h00;      memory[28048] <=  8'h00;      memory[28049] <=  8'h00;      memory[28050] <=  8'h00;      memory[28051] <=  8'h00;      memory[28052] <=  8'h00;      memory[28053] <=  8'h00;      memory[28054] <=  8'h00;      memory[28055] <=  8'h00;      memory[28056] <=  8'h00;      memory[28057] <=  8'h00;      memory[28058] <=  8'h00;      memory[28059] <=  8'h00;      memory[28060] <=  8'h00;      memory[28061] <=  8'h00;      memory[28062] <=  8'h00;      memory[28063] <=  8'h00;      memory[28064] <=  8'h00;      memory[28065] <=  8'h00;      memory[28066] <=  8'h00;      memory[28067] <=  8'h00;      memory[28068] <=  8'h00;      memory[28069] <=  8'h00;      memory[28070] <=  8'h00;      memory[28071] <=  8'h00;      memory[28072] <=  8'h00;      memory[28073] <=  8'h00;      memory[28074] <=  8'h00;      memory[28075] <=  8'h00;      memory[28076] <=  8'h00;      memory[28077] <=  8'h00;      memory[28078] <=  8'h00;      memory[28079] <=  8'h00;      memory[28080] <=  8'h00;      memory[28081] <=  8'h00;      memory[28082] <=  8'h00;      memory[28083] <=  8'h00;      memory[28084] <=  8'h00;      memory[28085] <=  8'h00;      memory[28086] <=  8'h00;      memory[28087] <=  8'h00;      memory[28088] <=  8'h00;      memory[28089] <=  8'h00;      memory[28090] <=  8'h00;      memory[28091] <=  8'h00;      memory[28092] <=  8'h00;      memory[28093] <=  8'h00;      memory[28094] <=  8'h00;      memory[28095] <=  8'h00;      memory[28096] <=  8'h00;      memory[28097] <=  8'h00;      memory[28098] <=  8'h00;      memory[28099] <=  8'h00;      memory[28100] <=  8'h00;      memory[28101] <=  8'h00;      memory[28102] <=  8'h00;      memory[28103] <=  8'h00;      memory[28104] <=  8'h00;      memory[28105] <=  8'h00;      memory[28106] <=  8'h00;      memory[28107] <=  8'h00;      memory[28108] <=  8'h00;      memory[28109] <=  8'h00;      memory[28110] <=  8'h00;      memory[28111] <=  8'h00;      memory[28112] <=  8'h00;      memory[28113] <=  8'h00;      memory[28114] <=  8'h00;      memory[28115] <=  8'h00;      memory[28116] <=  8'h00;      memory[28117] <=  8'h00;      memory[28118] <=  8'h00;      memory[28119] <=  8'h00;      memory[28120] <=  8'h00;      memory[28121] <=  8'h00;      memory[28122] <=  8'h00;      memory[28123] <=  8'h00;      memory[28124] <=  8'h00;      memory[28125] <=  8'h00;      memory[28126] <=  8'h00;      memory[28127] <=  8'h00;      memory[28128] <=  8'h00;      memory[28129] <=  8'h00;      memory[28130] <=  8'h00;      memory[28131] <=  8'h00;      memory[28132] <=  8'h00;      memory[28133] <=  8'h00;      memory[28134] <=  8'h00;      memory[28135] <=  8'h00;      memory[28136] <=  8'h00;      memory[28137] <=  8'h00;      memory[28138] <=  8'h00;      memory[28139] <=  8'h00;      memory[28140] <=  8'h00;      memory[28141] <=  8'h00;      memory[28142] <=  8'h00;      memory[28143] <=  8'h00;      memory[28144] <=  8'h00;      memory[28145] <=  8'h00;      memory[28146] <=  8'h00;      memory[28147] <=  8'h00;      memory[28148] <=  8'h00;      memory[28149] <=  8'h00;      memory[28150] <=  8'h00;      memory[28151] <=  8'h00;      memory[28152] <=  8'h00;      memory[28153] <=  8'h00;      memory[28154] <=  8'h00;      memory[28155] <=  8'h00;      memory[28156] <=  8'h00;      memory[28157] <=  8'h00;      memory[28158] <=  8'h00;      memory[28159] <=  8'h00;      memory[28160] <=  8'h00;      memory[28161] <=  8'h00;      memory[28162] <=  8'h00;      memory[28163] <=  8'h00;      memory[28164] <=  8'h00;      memory[28165] <=  8'h00;      memory[28166] <=  8'h00;      memory[28167] <=  8'h00;      memory[28168] <=  8'h00;      memory[28169] <=  8'h00;      memory[28170] <=  8'h00;      memory[28171] <=  8'h00;      memory[28172] <=  8'h00;      memory[28173] <=  8'h00;      memory[28174] <=  8'h00;      memory[28175] <=  8'h00;      memory[28176] <=  8'h00;      memory[28177] <=  8'h00;      memory[28178] <=  8'h00;      memory[28179] <=  8'h00;      memory[28180] <=  8'h00;      memory[28181] <=  8'h00;      memory[28182] <=  8'h00;      memory[28183] <=  8'h00;      memory[28184] <=  8'h00;      memory[28185] <=  8'h00;      memory[28186] <=  8'h00;      memory[28187] <=  8'h00;      memory[28188] <=  8'h00;      memory[28189] <=  8'h00;      memory[28190] <=  8'h00;      memory[28191] <=  8'h00;      memory[28192] <=  8'h00;      memory[28193] <=  8'h00;      memory[28194] <=  8'h00;      memory[28195] <=  8'h00;      memory[28196] <=  8'h00;      memory[28197] <=  8'h00;      memory[28198] <=  8'h00;      memory[28199] <=  8'h00;      memory[28200] <=  8'h00;      memory[28201] <=  8'h00;      memory[28202] <=  8'h00;      memory[28203] <=  8'h00;      memory[28204] <=  8'h00;      memory[28205] <=  8'h00;      memory[28206] <=  8'h00;      memory[28207] <=  8'h00;      memory[28208] <=  8'h00;      memory[28209] <=  8'h00;      memory[28210] <=  8'h00;      memory[28211] <=  8'h00;      memory[28212] <=  8'h00;      memory[28213] <=  8'h00;      memory[28214] <=  8'h00;      memory[28215] <=  8'h00;      memory[28216] <=  8'h00;      memory[28217] <=  8'h00;      memory[28218] <=  8'h00;      memory[28219] <=  8'h00;      memory[28220] <=  8'h00;      memory[28221] <=  8'h00;      memory[28222] <=  8'h00;      memory[28223] <=  8'h00;      memory[28224] <=  8'h00;      memory[28225] <=  8'h00;      memory[28226] <=  8'h00;      memory[28227] <=  8'h00;      memory[28228] <=  8'h00;      memory[28229] <=  8'h00;      memory[28230] <=  8'h00;      memory[28231] <=  8'h00;      memory[28232] <=  8'h00;      memory[28233] <=  8'h00;      memory[28234] <=  8'h00;      memory[28235] <=  8'h00;      memory[28236] <=  8'h00;      memory[28237] <=  8'h00;      memory[28238] <=  8'h00;      memory[28239] <=  8'h00;      memory[28240] <=  8'h00;      memory[28241] <=  8'h00;      memory[28242] <=  8'h00;      memory[28243] <=  8'h00;      memory[28244] <=  8'h00;      memory[28245] <=  8'h00;      memory[28246] <=  8'h00;      memory[28247] <=  8'h00;      memory[28248] <=  8'h00;      memory[28249] <=  8'h00;      memory[28250] <=  8'h00;      memory[28251] <=  8'h00;      memory[28252] <=  8'h00;      memory[28253] <=  8'h00;      memory[28254] <=  8'h00;      memory[28255] <=  8'h00;      memory[28256] <=  8'h00;      memory[28257] <=  8'h00;      memory[28258] <=  8'h00;      memory[28259] <=  8'h00;      memory[28260] <=  8'h00;      memory[28261] <=  8'h00;      memory[28262] <=  8'h00;      memory[28263] <=  8'h00;      memory[28264] <=  8'h00;      memory[28265] <=  8'h00;      memory[28266] <=  8'h00;      memory[28267] <=  8'h00;      memory[28268] <=  8'h00;      memory[28269] <=  8'h00;      memory[28270] <=  8'h00;      memory[28271] <=  8'h00;      memory[28272] <=  8'h00;      memory[28273] <=  8'h00;      memory[28274] <=  8'h00;      memory[28275] <=  8'h00;      memory[28276] <=  8'h00;      memory[28277] <=  8'h00;      memory[28278] <=  8'h00;      memory[28279] <=  8'h00;      memory[28280] <=  8'h00;      memory[28281] <=  8'h00;      memory[28282] <=  8'h00;      memory[28283] <=  8'h00;      memory[28284] <=  8'h00;      memory[28285] <=  8'h00;      memory[28286] <=  8'h00;      memory[28287] <=  8'h00;      memory[28288] <=  8'h00;      memory[28289] <=  8'h00;      memory[28290] <=  8'h00;      memory[28291] <=  8'h00;      memory[28292] <=  8'h00;      memory[28293] <=  8'h00;      memory[28294] <=  8'h00;      memory[28295] <=  8'h00;      memory[28296] <=  8'h00;      memory[28297] <=  8'h00;      memory[28298] <=  8'h00;      memory[28299] <=  8'h00;      memory[28300] <=  8'h00;      memory[28301] <=  8'h00;      memory[28302] <=  8'h00;      memory[28303] <=  8'h00;      memory[28304] <=  8'h00;      memory[28305] <=  8'h00;      memory[28306] <=  8'h00;      memory[28307] <=  8'h00;      memory[28308] <=  8'h00;      memory[28309] <=  8'h00;      memory[28310] <=  8'h00;      memory[28311] <=  8'h00;      memory[28312] <=  8'h00;      memory[28313] <=  8'h00;      memory[28314] <=  8'h00;      memory[28315] <=  8'h00;      memory[28316] <=  8'h00;      memory[28317] <=  8'h00;      memory[28318] <=  8'h00;      memory[28319] <=  8'h00;      memory[28320] <=  8'h00;      memory[28321] <=  8'h00;      memory[28322] <=  8'h00;      memory[28323] <=  8'h00;      memory[28324] <=  8'h00;      memory[28325] <=  8'h00;      memory[28326] <=  8'h00;      memory[28327] <=  8'h00;      memory[28328] <=  8'h00;      memory[28329] <=  8'h00;      memory[28330] <=  8'h00;      memory[28331] <=  8'h00;      memory[28332] <=  8'h00;      memory[28333] <=  8'h00;      memory[28334] <=  8'h00;      memory[28335] <=  8'h00;      memory[28336] <=  8'h00;      memory[28337] <=  8'h00;      memory[28338] <=  8'h00;      memory[28339] <=  8'h00;      memory[28340] <=  8'h00;      memory[28341] <=  8'h00;      memory[28342] <=  8'h00;      memory[28343] <=  8'h00;      memory[28344] <=  8'h00;      memory[28345] <=  8'h00;      memory[28346] <=  8'h00;      memory[28347] <=  8'h00;      memory[28348] <=  8'h00;      memory[28349] <=  8'h00;      memory[28350] <=  8'h00;      memory[28351] <=  8'h00;      memory[28352] <=  8'h00;      memory[28353] <=  8'h00;      memory[28354] <=  8'h00;      memory[28355] <=  8'h00;      memory[28356] <=  8'h00;      memory[28357] <=  8'h00;      memory[28358] <=  8'h00;      memory[28359] <=  8'h00;      memory[28360] <=  8'h00;      memory[28361] <=  8'h00;      memory[28362] <=  8'h00;      memory[28363] <=  8'h00;      memory[28364] <=  8'h00;      memory[28365] <=  8'h00;      memory[28366] <=  8'h00;      memory[28367] <=  8'h00;      memory[28368] <=  8'h00;      memory[28369] <=  8'h00;      memory[28370] <=  8'h00;      memory[28371] <=  8'h00;      memory[28372] <=  8'h00;      memory[28373] <=  8'h00;      memory[28374] <=  8'h00;      memory[28375] <=  8'h00;      memory[28376] <=  8'h00;      memory[28377] <=  8'h00;      memory[28378] <=  8'h00;      memory[28379] <=  8'h00;      memory[28380] <=  8'h00;      memory[28381] <=  8'h00;      memory[28382] <=  8'h00;      memory[28383] <=  8'h00;      memory[28384] <=  8'h00;      memory[28385] <=  8'h00;      memory[28386] <=  8'h00;      memory[28387] <=  8'h00;      memory[28388] <=  8'h00;      memory[28389] <=  8'h00;      memory[28390] <=  8'h00;      memory[28391] <=  8'h00;      memory[28392] <=  8'h00;      memory[28393] <=  8'h00;      memory[28394] <=  8'h00;      memory[28395] <=  8'h00;      memory[28396] <=  8'h00;      memory[28397] <=  8'h00;      memory[28398] <=  8'h00;      memory[28399] <=  8'h00;      memory[28400] <=  8'h00;      memory[28401] <=  8'h00;      memory[28402] <=  8'h00;      memory[28403] <=  8'h00;      memory[28404] <=  8'h00;      memory[28405] <=  8'h00;      memory[28406] <=  8'h00;      memory[28407] <=  8'h00;      memory[28408] <=  8'h00;      memory[28409] <=  8'h00;      memory[28410] <=  8'h00;      memory[28411] <=  8'h00;      memory[28412] <=  8'h00;      memory[28413] <=  8'h00;      memory[28414] <=  8'h00;      memory[28415] <=  8'h00;      memory[28416] <=  8'h00;      memory[28417] <=  8'h00;      memory[28418] <=  8'h00;      memory[28419] <=  8'h00;      memory[28420] <=  8'h00;      memory[28421] <=  8'h00;      memory[28422] <=  8'h00;      memory[28423] <=  8'h00;      memory[28424] <=  8'h00;      memory[28425] <=  8'h00;      memory[28426] <=  8'h00;      memory[28427] <=  8'h00;      memory[28428] <=  8'h00;      memory[28429] <=  8'h00;      memory[28430] <=  8'h00;      memory[28431] <=  8'h00;      memory[28432] <=  8'h00;      memory[28433] <=  8'h00;      memory[28434] <=  8'h00;      memory[28435] <=  8'h00;      memory[28436] <=  8'h00;      memory[28437] <=  8'h00;      memory[28438] <=  8'h00;      memory[28439] <=  8'h00;      memory[28440] <=  8'h00;      memory[28441] <=  8'h00;      memory[28442] <=  8'h00;      memory[28443] <=  8'h00;      memory[28444] <=  8'h00;      memory[28445] <=  8'h00;      memory[28446] <=  8'h00;      memory[28447] <=  8'h00;      memory[28448] <=  8'h00;      memory[28449] <=  8'h00;      memory[28450] <=  8'h00;      memory[28451] <=  8'h00;      memory[28452] <=  8'h00;      memory[28453] <=  8'h00;      memory[28454] <=  8'h00;      memory[28455] <=  8'h00;      memory[28456] <=  8'h00;      memory[28457] <=  8'h00;      memory[28458] <=  8'h00;      memory[28459] <=  8'h00;      memory[28460] <=  8'h00;      memory[28461] <=  8'h00;      memory[28462] <=  8'h00;      memory[28463] <=  8'h00;      memory[28464] <=  8'h00;      memory[28465] <=  8'h00;      memory[28466] <=  8'h00;      memory[28467] <=  8'h00;      memory[28468] <=  8'h00;      memory[28469] <=  8'h00;      memory[28470] <=  8'h00;      memory[28471] <=  8'h00;      memory[28472] <=  8'h00;      memory[28473] <=  8'h00;      memory[28474] <=  8'h00;      memory[28475] <=  8'h00;      memory[28476] <=  8'h00;      memory[28477] <=  8'h00;      memory[28478] <=  8'h00;      memory[28479] <=  8'h00;      memory[28480] <=  8'h00;      memory[28481] <=  8'h00;      memory[28482] <=  8'h00;      memory[28483] <=  8'h00;      memory[28484] <=  8'h00;      memory[28485] <=  8'h00;      memory[28486] <=  8'h00;      memory[28487] <=  8'h00;      memory[28488] <=  8'h00;      memory[28489] <=  8'h00;      memory[28490] <=  8'h00;      memory[28491] <=  8'h00;      memory[28492] <=  8'h00;      memory[28493] <=  8'h00;      memory[28494] <=  8'h00;      memory[28495] <=  8'h00;      memory[28496] <=  8'h00;      memory[28497] <=  8'h00;      memory[28498] <=  8'h00;      memory[28499] <=  8'h00;      memory[28500] <=  8'h00;      memory[28501] <=  8'h00;      memory[28502] <=  8'h00;      memory[28503] <=  8'h00;      memory[28504] <=  8'h00;      memory[28505] <=  8'h00;      memory[28506] <=  8'h00;      memory[28507] <=  8'h00;      memory[28508] <=  8'h00;      memory[28509] <=  8'h00;      memory[28510] <=  8'h00;      memory[28511] <=  8'h00;      memory[28512] <=  8'h00;      memory[28513] <=  8'h00;      memory[28514] <=  8'h00;      memory[28515] <=  8'h00;      memory[28516] <=  8'h00;      memory[28517] <=  8'h00;      memory[28518] <=  8'h00;      memory[28519] <=  8'h00;      memory[28520] <=  8'h00;      memory[28521] <=  8'h00;      memory[28522] <=  8'h00;      memory[28523] <=  8'h00;      memory[28524] <=  8'h00;      memory[28525] <=  8'h00;      memory[28526] <=  8'h00;      memory[28527] <=  8'h00;      memory[28528] <=  8'h00;      memory[28529] <=  8'h00;      memory[28530] <=  8'h00;      memory[28531] <=  8'h00;      memory[28532] <=  8'h00;      memory[28533] <=  8'h00;      memory[28534] <=  8'h00;      memory[28535] <=  8'h00;      memory[28536] <=  8'h00;      memory[28537] <=  8'h00;      memory[28538] <=  8'h00;      memory[28539] <=  8'h00;      memory[28540] <=  8'h00;      memory[28541] <=  8'h00;      memory[28542] <=  8'h00;      memory[28543] <=  8'h00;      memory[28544] <=  8'h00;      memory[28545] <=  8'h00;      memory[28546] <=  8'h00;      memory[28547] <=  8'h00;      memory[28548] <=  8'h00;      memory[28549] <=  8'h00;      memory[28550] <=  8'h00;      memory[28551] <=  8'h00;      memory[28552] <=  8'h00;      memory[28553] <=  8'h00;      memory[28554] <=  8'h00;      memory[28555] <=  8'h00;      memory[28556] <=  8'h00;      memory[28557] <=  8'h00;      memory[28558] <=  8'h00;      memory[28559] <=  8'h00;      memory[28560] <=  8'h00;      memory[28561] <=  8'h00;      memory[28562] <=  8'h00;      memory[28563] <=  8'h00;      memory[28564] <=  8'h00;      memory[28565] <=  8'h00;      memory[28566] <=  8'h00;      memory[28567] <=  8'h00;      memory[28568] <=  8'h00;      memory[28569] <=  8'h00;      memory[28570] <=  8'h00;      memory[28571] <=  8'h00;      memory[28572] <=  8'h00;      memory[28573] <=  8'h00;      memory[28574] <=  8'h00;      memory[28575] <=  8'h00;      memory[28576] <=  8'h00;      memory[28577] <=  8'h00;      memory[28578] <=  8'h00;      memory[28579] <=  8'h00;      memory[28580] <=  8'h00;      memory[28581] <=  8'h00;      memory[28582] <=  8'h00;      memory[28583] <=  8'h00;      memory[28584] <=  8'h00;      memory[28585] <=  8'h00;      memory[28586] <=  8'h00;      memory[28587] <=  8'h00;      memory[28588] <=  8'h00;      memory[28589] <=  8'h00;      memory[28590] <=  8'h00;      memory[28591] <=  8'h00;      memory[28592] <=  8'h00;      memory[28593] <=  8'h00;      memory[28594] <=  8'h00;      memory[28595] <=  8'h00;      memory[28596] <=  8'h00;      memory[28597] <=  8'h00;      memory[28598] <=  8'h00;      memory[28599] <=  8'h00;      memory[28600] <=  8'h00;      memory[28601] <=  8'h00;      memory[28602] <=  8'h00;      memory[28603] <=  8'h00;      memory[28604] <=  8'h00;      memory[28605] <=  8'h00;      memory[28606] <=  8'h00;      memory[28607] <=  8'h00;      memory[28608] <=  8'h00;      memory[28609] <=  8'h00;      memory[28610] <=  8'h00;      memory[28611] <=  8'h00;      memory[28612] <=  8'h00;      memory[28613] <=  8'h00;      memory[28614] <=  8'h00;      memory[28615] <=  8'h00;      memory[28616] <=  8'h00;      memory[28617] <=  8'h00;      memory[28618] <=  8'h00;      memory[28619] <=  8'h00;      memory[28620] <=  8'h00;      memory[28621] <=  8'h00;      memory[28622] <=  8'h00;      memory[28623] <=  8'h00;      memory[28624] <=  8'h00;      memory[28625] <=  8'h00;      memory[28626] <=  8'h00;      memory[28627] <=  8'h00;      memory[28628] <=  8'h00;      memory[28629] <=  8'h00;      memory[28630] <=  8'h00;      memory[28631] <=  8'h00;      memory[28632] <=  8'h00;      memory[28633] <=  8'h00;      memory[28634] <=  8'h00;      memory[28635] <=  8'h00;      memory[28636] <=  8'h00;      memory[28637] <=  8'h00;      memory[28638] <=  8'h00;      memory[28639] <=  8'h00;      memory[28640] <=  8'h00;      memory[28641] <=  8'h00;      memory[28642] <=  8'h00;      memory[28643] <=  8'h00;      memory[28644] <=  8'h00;      memory[28645] <=  8'h00;      memory[28646] <=  8'h00;      memory[28647] <=  8'h00;      memory[28648] <=  8'h00;      memory[28649] <=  8'h00;      memory[28650] <=  8'h00;      memory[28651] <=  8'h00;      memory[28652] <=  8'h00;      memory[28653] <=  8'h00;      memory[28654] <=  8'h00;      memory[28655] <=  8'h00;      memory[28656] <=  8'h00;      memory[28657] <=  8'h00;      memory[28658] <=  8'h00;      memory[28659] <=  8'h00;      memory[28660] <=  8'h00;      memory[28661] <=  8'h00;      memory[28662] <=  8'h00;      memory[28663] <=  8'h00;      memory[28664] <=  8'h00;      memory[28665] <=  8'h00;      memory[28666] <=  8'h00;      memory[28667] <=  8'h00;      memory[28668] <=  8'h00;      memory[28669] <=  8'h00;      memory[28670] <=  8'h00;      memory[28671] <=  8'h00;      memory[28672] <=  8'h00;      memory[28673] <=  8'h00;      memory[28674] <=  8'h00;      memory[28675] <=  8'h00;      memory[28676] <=  8'h00;      memory[28677] <=  8'h00;      memory[28678] <=  8'h00;      memory[28679] <=  8'h00;      memory[28680] <=  8'h00;      memory[28681] <=  8'h00;      memory[28682] <=  8'h00;      memory[28683] <=  8'h00;      memory[28684] <=  8'h00;      memory[28685] <=  8'h00;      memory[28686] <=  8'h00;      memory[28687] <=  8'h00;      memory[28688] <=  8'h00;      memory[28689] <=  8'h00;      memory[28690] <=  8'h00;      memory[28691] <=  8'h00;      memory[28692] <=  8'h00;      memory[28693] <=  8'h00;      memory[28694] <=  8'h00;      memory[28695] <=  8'h00;      memory[28696] <=  8'h00;      memory[28697] <=  8'h00;      memory[28698] <=  8'h00;      memory[28699] <=  8'h00;      memory[28700] <=  8'h00;      memory[28701] <=  8'h00;      memory[28702] <=  8'h00;      memory[28703] <=  8'h00;      memory[28704] <=  8'h00;      memory[28705] <=  8'h00;      memory[28706] <=  8'h00;      memory[28707] <=  8'h00;      memory[28708] <=  8'h00;      memory[28709] <=  8'h00;      memory[28710] <=  8'h00;      memory[28711] <=  8'h00;      memory[28712] <=  8'h00;      memory[28713] <=  8'h00;      memory[28714] <=  8'h00;      memory[28715] <=  8'h00;      memory[28716] <=  8'h00;      memory[28717] <=  8'h00;      memory[28718] <=  8'h00;      memory[28719] <=  8'h00;      memory[28720] <=  8'h00;      memory[28721] <=  8'h00;      memory[28722] <=  8'h00;      memory[28723] <=  8'h00;      memory[28724] <=  8'h00;      memory[28725] <=  8'h00;      memory[28726] <=  8'h00;      memory[28727] <=  8'h00;      memory[28728] <=  8'h00;      memory[28729] <=  8'h00;      memory[28730] <=  8'h00;      memory[28731] <=  8'h00;      memory[28732] <=  8'h00;      memory[28733] <=  8'h00;      memory[28734] <=  8'h00;      memory[28735] <=  8'h00;      memory[28736] <=  8'h00;      memory[28737] <=  8'h00;      memory[28738] <=  8'h00;      memory[28739] <=  8'h00;      memory[28740] <=  8'h00;      memory[28741] <=  8'h00;      memory[28742] <=  8'h00;      memory[28743] <=  8'h00;      memory[28744] <=  8'h00;      memory[28745] <=  8'h00;      memory[28746] <=  8'h00;      memory[28747] <=  8'h00;      memory[28748] <=  8'h00;      memory[28749] <=  8'h00;      memory[28750] <=  8'h00;      memory[28751] <=  8'h00;      memory[28752] <=  8'h00;      memory[28753] <=  8'h00;      memory[28754] <=  8'h00;      memory[28755] <=  8'h00;      memory[28756] <=  8'h00;      memory[28757] <=  8'h00;      memory[28758] <=  8'h00;      memory[28759] <=  8'h00;      memory[28760] <=  8'h00;      memory[28761] <=  8'h00;      memory[28762] <=  8'h00;      memory[28763] <=  8'h00;      memory[28764] <=  8'h00;      memory[28765] <=  8'h00;      memory[28766] <=  8'h00;      memory[28767] <=  8'h00;      memory[28768] <=  8'h00;      memory[28769] <=  8'h00;      memory[28770] <=  8'h00;      memory[28771] <=  8'h00;      memory[28772] <=  8'h00;      memory[28773] <=  8'h00;      memory[28774] <=  8'h00;      memory[28775] <=  8'h00;      memory[28776] <=  8'h00;      memory[28777] <=  8'h00;      memory[28778] <=  8'h00;      memory[28779] <=  8'h00;      memory[28780] <=  8'h00;      memory[28781] <=  8'h00;      memory[28782] <=  8'h00;      memory[28783] <=  8'h00;      memory[28784] <=  8'h00;      memory[28785] <=  8'h00;      memory[28786] <=  8'h00;      memory[28787] <=  8'h00;      memory[28788] <=  8'h00;      memory[28789] <=  8'h00;      memory[28790] <=  8'h00;      memory[28791] <=  8'h00;      memory[28792] <=  8'h00;      memory[28793] <=  8'h00;      memory[28794] <=  8'h00;      memory[28795] <=  8'h00;      memory[28796] <=  8'h00;      memory[28797] <=  8'h00;      memory[28798] <=  8'h00;      memory[28799] <=  8'h00;      memory[28800] <=  8'h00;      memory[28801] <=  8'h00;      memory[28802] <=  8'h00;      memory[28803] <=  8'h00;      memory[28804] <=  8'h00;      memory[28805] <=  8'h00;      memory[28806] <=  8'h00;      memory[28807] <=  8'h00;      memory[28808] <=  8'h00;      memory[28809] <=  8'h00;      memory[28810] <=  8'h00;      memory[28811] <=  8'h00;      memory[28812] <=  8'h00;      memory[28813] <=  8'h00;      memory[28814] <=  8'h00;      memory[28815] <=  8'h00;      memory[28816] <=  8'h00;      memory[28817] <=  8'h00;      memory[28818] <=  8'h00;      memory[28819] <=  8'h00;      memory[28820] <=  8'h00;      memory[28821] <=  8'h00;      memory[28822] <=  8'h00;      memory[28823] <=  8'h00;      memory[28824] <=  8'h00;      memory[28825] <=  8'h00;      memory[28826] <=  8'h00;      memory[28827] <=  8'h00;      memory[28828] <=  8'h00;      memory[28829] <=  8'h00;      memory[28830] <=  8'h00;      memory[28831] <=  8'h00;      memory[28832] <=  8'h00;      memory[28833] <=  8'h00;      memory[28834] <=  8'h00;      memory[28835] <=  8'h00;      memory[28836] <=  8'h00;      memory[28837] <=  8'h00;      memory[28838] <=  8'h00;      memory[28839] <=  8'h00;      memory[28840] <=  8'h00;      memory[28841] <=  8'h00;      memory[28842] <=  8'h00;      memory[28843] <=  8'h00;      memory[28844] <=  8'h00;      memory[28845] <=  8'h00;      memory[28846] <=  8'h00;      memory[28847] <=  8'h00;      memory[28848] <=  8'h00;      memory[28849] <=  8'h00;      memory[28850] <=  8'h00;      memory[28851] <=  8'h00;      memory[28852] <=  8'h00;      memory[28853] <=  8'h00;      memory[28854] <=  8'h00;      memory[28855] <=  8'h00;      memory[28856] <=  8'h00;      memory[28857] <=  8'h00;      memory[28858] <=  8'h00;      memory[28859] <=  8'h00;      memory[28860] <=  8'h00;      memory[28861] <=  8'h00;      memory[28862] <=  8'h00;      memory[28863] <=  8'h00;      memory[28864] <=  8'h00;      memory[28865] <=  8'h00;      memory[28866] <=  8'h00;      memory[28867] <=  8'h00;      memory[28868] <=  8'h00;      memory[28869] <=  8'h00;      memory[28870] <=  8'h00;      memory[28871] <=  8'h00;      memory[28872] <=  8'h00;      memory[28873] <=  8'h00;      memory[28874] <=  8'h00;      memory[28875] <=  8'h00;      memory[28876] <=  8'h00;      memory[28877] <=  8'h00;      memory[28878] <=  8'h00;      memory[28879] <=  8'h00;      memory[28880] <=  8'h00;      memory[28881] <=  8'h00;      memory[28882] <=  8'h00;      memory[28883] <=  8'h00;      memory[28884] <=  8'h00;      memory[28885] <=  8'h00;      memory[28886] <=  8'h00;      memory[28887] <=  8'h00;      memory[28888] <=  8'h00;      memory[28889] <=  8'h00;      memory[28890] <=  8'h00;      memory[28891] <=  8'h00;      memory[28892] <=  8'h00;      memory[28893] <=  8'h00;      memory[28894] <=  8'h00;      memory[28895] <=  8'h00;      memory[28896] <=  8'h00;      memory[28897] <=  8'h00;      memory[28898] <=  8'h00;      memory[28899] <=  8'h00;      memory[28900] <=  8'h00;      memory[28901] <=  8'h00;      memory[28902] <=  8'h00;      memory[28903] <=  8'h00;      memory[28904] <=  8'h00;      memory[28905] <=  8'h00;      memory[28906] <=  8'h00;      memory[28907] <=  8'h00;      memory[28908] <=  8'h00;      memory[28909] <=  8'h00;      memory[28910] <=  8'h00;      memory[28911] <=  8'h00;      memory[28912] <=  8'h00;      memory[28913] <=  8'h00;      memory[28914] <=  8'h00;      memory[28915] <=  8'h00;      memory[28916] <=  8'h00;      memory[28917] <=  8'h00;      memory[28918] <=  8'h00;      memory[28919] <=  8'h00;      memory[28920] <=  8'h00;      memory[28921] <=  8'h00;      memory[28922] <=  8'h00;      memory[28923] <=  8'h00;      memory[28924] <=  8'h00;      memory[28925] <=  8'h00;      memory[28926] <=  8'h00;      memory[28927] <=  8'h00;      memory[28928] <=  8'h00;      memory[28929] <=  8'h00;      memory[28930] <=  8'h00;      memory[28931] <=  8'h00;      memory[28932] <=  8'h00;      memory[28933] <=  8'h00;      memory[28934] <=  8'h00;      memory[28935] <=  8'h00;      memory[28936] <=  8'h00;      memory[28937] <=  8'h00;      memory[28938] <=  8'h00;      memory[28939] <=  8'h00;      memory[28940] <=  8'h00;      memory[28941] <=  8'h00;      memory[28942] <=  8'h00;      memory[28943] <=  8'h00;      memory[28944] <=  8'h00;      memory[28945] <=  8'h00;      memory[28946] <=  8'h00;      memory[28947] <=  8'h00;      memory[28948] <=  8'h00;      memory[28949] <=  8'h00;      memory[28950] <=  8'h00;      memory[28951] <=  8'h00;      memory[28952] <=  8'h00;      memory[28953] <=  8'h00;      memory[28954] <=  8'h00;      memory[28955] <=  8'h00;      memory[28956] <=  8'h00;      memory[28957] <=  8'h00;      memory[28958] <=  8'h00;      memory[28959] <=  8'h00;      memory[28960] <=  8'h00;      memory[28961] <=  8'h00;      memory[28962] <=  8'h00;      memory[28963] <=  8'h00;      memory[28964] <=  8'h00;      memory[28965] <=  8'h00;      memory[28966] <=  8'h00;      memory[28967] <=  8'h00;      memory[28968] <=  8'h00;      memory[28969] <=  8'h00;      memory[28970] <=  8'h00;      memory[28971] <=  8'h00;      memory[28972] <=  8'h00;      memory[28973] <=  8'h00;      memory[28974] <=  8'h00;      memory[28975] <=  8'h00;      memory[28976] <=  8'h00;      memory[28977] <=  8'h00;      memory[28978] <=  8'h00;      memory[28979] <=  8'h00;      memory[28980] <=  8'h00;      memory[28981] <=  8'h00;      memory[28982] <=  8'h00;      memory[28983] <=  8'h00;      memory[28984] <=  8'h00;      memory[28985] <=  8'h00;      memory[28986] <=  8'h00;      memory[28987] <=  8'h00;      memory[28988] <=  8'h00;      memory[28989] <=  8'h00;      memory[28990] <=  8'h00;      memory[28991] <=  8'h00;      memory[28992] <=  8'h00;      memory[28993] <=  8'h00;      memory[28994] <=  8'h00;      memory[28995] <=  8'h00;      memory[28996] <=  8'h00;      memory[28997] <=  8'h00;      memory[28998] <=  8'h00;      memory[28999] <=  8'h00;      memory[29000] <=  8'h00;      memory[29001] <=  8'h00;      memory[29002] <=  8'h00;      memory[29003] <=  8'h00;      memory[29004] <=  8'h00;      memory[29005] <=  8'h00;      memory[29006] <=  8'h00;      memory[29007] <=  8'h00;      memory[29008] <=  8'h00;      memory[29009] <=  8'h00;      memory[29010] <=  8'h00;      memory[29011] <=  8'h00;      memory[29012] <=  8'h00;      memory[29013] <=  8'h00;      memory[29014] <=  8'h00;      memory[29015] <=  8'h00;      memory[29016] <=  8'h00;      memory[29017] <=  8'h00;      memory[29018] <=  8'h00;      memory[29019] <=  8'h00;      memory[29020] <=  8'h00;      memory[29021] <=  8'h00;      memory[29022] <=  8'h00;      memory[29023] <=  8'h00;      memory[29024] <=  8'h00;      memory[29025] <=  8'h00;      memory[29026] <=  8'h00;      memory[29027] <=  8'h00;      memory[29028] <=  8'h00;      memory[29029] <=  8'h00;      memory[29030] <=  8'h00;      memory[29031] <=  8'h00;      memory[29032] <=  8'h00;      memory[29033] <=  8'h00;      memory[29034] <=  8'h00;      memory[29035] <=  8'h00;      memory[29036] <=  8'h00;      memory[29037] <=  8'h00;      memory[29038] <=  8'h00;      memory[29039] <=  8'h00;      memory[29040] <=  8'h00;      memory[29041] <=  8'h00;      memory[29042] <=  8'h00;      memory[29043] <=  8'h00;      memory[29044] <=  8'h00;      memory[29045] <=  8'h00;      memory[29046] <=  8'h00;      memory[29047] <=  8'h00;      memory[29048] <=  8'h00;      memory[29049] <=  8'h00;      memory[29050] <=  8'h00;      memory[29051] <=  8'h00;      memory[29052] <=  8'h00;      memory[29053] <=  8'h00;      memory[29054] <=  8'h00;      memory[29055] <=  8'h00;      memory[29056] <=  8'h00;      memory[29057] <=  8'h00;      memory[29058] <=  8'h00;      memory[29059] <=  8'h00;      memory[29060] <=  8'h00;      memory[29061] <=  8'h00;      memory[29062] <=  8'h00;      memory[29063] <=  8'h00;      memory[29064] <=  8'h00;      memory[29065] <=  8'h00;      memory[29066] <=  8'h00;      memory[29067] <=  8'h00;      memory[29068] <=  8'h00;      memory[29069] <=  8'h00;      memory[29070] <=  8'h00;      memory[29071] <=  8'h00;      memory[29072] <=  8'h00;      memory[29073] <=  8'h00;      memory[29074] <=  8'h00;      memory[29075] <=  8'h00;      memory[29076] <=  8'h00;      memory[29077] <=  8'h00;      memory[29078] <=  8'h00;      memory[29079] <=  8'h00;      memory[29080] <=  8'h00;      memory[29081] <=  8'h00;      memory[29082] <=  8'h00;      memory[29083] <=  8'h00;      memory[29084] <=  8'h00;      memory[29085] <=  8'h00;      memory[29086] <=  8'h00;      memory[29087] <=  8'h00;      memory[29088] <=  8'h00;      memory[29089] <=  8'h00;      memory[29090] <=  8'h00;      memory[29091] <=  8'h00;      memory[29092] <=  8'h00;      memory[29093] <=  8'h00;      memory[29094] <=  8'h00;      memory[29095] <=  8'h00;      memory[29096] <=  8'h00;      memory[29097] <=  8'h00;      memory[29098] <=  8'h00;      memory[29099] <=  8'h00;      memory[29100] <=  8'h00;      memory[29101] <=  8'h00;      memory[29102] <=  8'h00;      memory[29103] <=  8'h00;      memory[29104] <=  8'h00;      memory[29105] <=  8'h00;      memory[29106] <=  8'h00;      memory[29107] <=  8'h00;      memory[29108] <=  8'h00;      memory[29109] <=  8'h00;      memory[29110] <=  8'h00;      memory[29111] <=  8'h00;      memory[29112] <=  8'h00;      memory[29113] <=  8'h00;      memory[29114] <=  8'h00;      memory[29115] <=  8'h00;      memory[29116] <=  8'h00;      memory[29117] <=  8'h00;      memory[29118] <=  8'h00;      memory[29119] <=  8'h00;      memory[29120] <=  8'h00;      memory[29121] <=  8'h00;      memory[29122] <=  8'h00;      memory[29123] <=  8'h00;      memory[29124] <=  8'h00;      memory[29125] <=  8'h00;      memory[29126] <=  8'h00;      memory[29127] <=  8'h00;      memory[29128] <=  8'h00;      memory[29129] <=  8'h00;      memory[29130] <=  8'h00;      memory[29131] <=  8'h00;      memory[29132] <=  8'h00;      memory[29133] <=  8'h00;      memory[29134] <=  8'h00;      memory[29135] <=  8'h00;      memory[29136] <=  8'h00;      memory[29137] <=  8'h00;      memory[29138] <=  8'h00;      memory[29139] <=  8'h00;      memory[29140] <=  8'h00;      memory[29141] <=  8'h00;      memory[29142] <=  8'h00;      memory[29143] <=  8'h00;      memory[29144] <=  8'h00;      memory[29145] <=  8'h00;      memory[29146] <=  8'h00;      memory[29147] <=  8'h00;      memory[29148] <=  8'h00;      memory[29149] <=  8'h00;      memory[29150] <=  8'h00;      memory[29151] <=  8'h00;      memory[29152] <=  8'h00;      memory[29153] <=  8'h00;      memory[29154] <=  8'h00;      memory[29155] <=  8'h00;      memory[29156] <=  8'h00;      memory[29157] <=  8'h00;      memory[29158] <=  8'h00;      memory[29159] <=  8'h00;      memory[29160] <=  8'h00;      memory[29161] <=  8'h00;      memory[29162] <=  8'h00;      memory[29163] <=  8'h00;      memory[29164] <=  8'h00;      memory[29165] <=  8'h00;      memory[29166] <=  8'h00;      memory[29167] <=  8'h00;      memory[29168] <=  8'h00;      memory[29169] <=  8'h00;      memory[29170] <=  8'h00;      memory[29171] <=  8'h00;      memory[29172] <=  8'h00;      memory[29173] <=  8'h00;      memory[29174] <=  8'h00;      memory[29175] <=  8'h00;      memory[29176] <=  8'h00;      memory[29177] <=  8'h00;      memory[29178] <=  8'h00;      memory[29179] <=  8'h00;      memory[29180] <=  8'h00;      memory[29181] <=  8'h00;      memory[29182] <=  8'h00;      memory[29183] <=  8'h00;      memory[29184] <=  8'h00;      memory[29185] <=  8'h00;      memory[29186] <=  8'h00;      memory[29187] <=  8'h00;      memory[29188] <=  8'h00;      memory[29189] <=  8'h00;      memory[29190] <=  8'h00;      memory[29191] <=  8'h00;      memory[29192] <=  8'h00;      memory[29193] <=  8'h00;      memory[29194] <=  8'h00;      memory[29195] <=  8'h00;      memory[29196] <=  8'h00;      memory[29197] <=  8'h00;      memory[29198] <=  8'h00;      memory[29199] <=  8'h00;      memory[29200] <=  8'h00;      memory[29201] <=  8'h00;      memory[29202] <=  8'h00;      memory[29203] <=  8'h00;      memory[29204] <=  8'h00;      memory[29205] <=  8'h00;      memory[29206] <=  8'h00;      memory[29207] <=  8'h00;      memory[29208] <=  8'h00;      memory[29209] <=  8'h00;      memory[29210] <=  8'h00;      memory[29211] <=  8'h00;      memory[29212] <=  8'h00;      memory[29213] <=  8'h00;      memory[29214] <=  8'h00;      memory[29215] <=  8'h00;      memory[29216] <=  8'h00;      memory[29217] <=  8'h00;      memory[29218] <=  8'h00;      memory[29219] <=  8'h00;      memory[29220] <=  8'h00;      memory[29221] <=  8'h00;      memory[29222] <=  8'h00;      memory[29223] <=  8'h00;      memory[29224] <=  8'h00;      memory[29225] <=  8'h00;      memory[29226] <=  8'h00;      memory[29227] <=  8'h00;      memory[29228] <=  8'h00;      memory[29229] <=  8'h00;      memory[29230] <=  8'h00;      memory[29231] <=  8'h00;      memory[29232] <=  8'h00;      memory[29233] <=  8'h00;      memory[29234] <=  8'h00;      memory[29235] <=  8'h00;      memory[29236] <=  8'h00;      memory[29237] <=  8'h00;      memory[29238] <=  8'h00;      memory[29239] <=  8'h00;      memory[29240] <=  8'h00;      memory[29241] <=  8'h00;      memory[29242] <=  8'h00;      memory[29243] <=  8'h00;      memory[29244] <=  8'h00;      memory[29245] <=  8'h00;      memory[29246] <=  8'h00;      memory[29247] <=  8'h00;      memory[29248] <=  8'h00;      memory[29249] <=  8'h00;      memory[29250] <=  8'h00;      memory[29251] <=  8'h00;      memory[29252] <=  8'h00;      memory[29253] <=  8'h00;      memory[29254] <=  8'h00;      memory[29255] <=  8'h00;      memory[29256] <=  8'h00;      memory[29257] <=  8'h00;      memory[29258] <=  8'h00;      memory[29259] <=  8'h00;      memory[29260] <=  8'h00;      memory[29261] <=  8'h00;      memory[29262] <=  8'h00;      memory[29263] <=  8'h00;      memory[29264] <=  8'h00;      memory[29265] <=  8'h00;      memory[29266] <=  8'h00;      memory[29267] <=  8'h00;      memory[29268] <=  8'h00;      memory[29269] <=  8'h00;      memory[29270] <=  8'h00;      memory[29271] <=  8'h00;      memory[29272] <=  8'h00;      memory[29273] <=  8'h00;      memory[29274] <=  8'h00;      memory[29275] <=  8'h00;      memory[29276] <=  8'h00;      memory[29277] <=  8'h00;      memory[29278] <=  8'h00;      memory[29279] <=  8'h00;      memory[29280] <=  8'h00;      memory[29281] <=  8'h00;      memory[29282] <=  8'h00;      memory[29283] <=  8'h00;      memory[29284] <=  8'h00;      memory[29285] <=  8'h00;      memory[29286] <=  8'h00;      memory[29287] <=  8'h00;      memory[29288] <=  8'h00;      memory[29289] <=  8'h00;      memory[29290] <=  8'h00;      memory[29291] <=  8'h00;      memory[29292] <=  8'h00;      memory[29293] <=  8'h00;      memory[29294] <=  8'h00;      memory[29295] <=  8'h00;      memory[29296] <=  8'h00;      memory[29297] <=  8'h00;      memory[29298] <=  8'h00;      memory[29299] <=  8'h00;      memory[29300] <=  8'h00;      memory[29301] <=  8'h00;      memory[29302] <=  8'h00;      memory[29303] <=  8'h00;      memory[29304] <=  8'h00;      memory[29305] <=  8'h00;      memory[29306] <=  8'h00;      memory[29307] <=  8'h00;      memory[29308] <=  8'h00;      memory[29309] <=  8'h00;      memory[29310] <=  8'h00;      memory[29311] <=  8'h00;      memory[29312] <=  8'h00;      memory[29313] <=  8'h00;      memory[29314] <=  8'h00;      memory[29315] <=  8'h00;      memory[29316] <=  8'h00;      memory[29317] <=  8'h00;      memory[29318] <=  8'h00;      memory[29319] <=  8'h00;      memory[29320] <=  8'h00;      memory[29321] <=  8'h00;      memory[29322] <=  8'h00;      memory[29323] <=  8'h00;      memory[29324] <=  8'h00;      memory[29325] <=  8'h00;      memory[29326] <=  8'h00;      memory[29327] <=  8'h00;      memory[29328] <=  8'h00;      memory[29329] <=  8'h00;      memory[29330] <=  8'h00;      memory[29331] <=  8'h00;      memory[29332] <=  8'h00;      memory[29333] <=  8'h00;      memory[29334] <=  8'h00;      memory[29335] <=  8'h00;      memory[29336] <=  8'h00;      memory[29337] <=  8'h00;      memory[29338] <=  8'h00;      memory[29339] <=  8'h00;      memory[29340] <=  8'h00;      memory[29341] <=  8'h00;      memory[29342] <=  8'h00;      memory[29343] <=  8'h00;      memory[29344] <=  8'h00;      memory[29345] <=  8'h00;      memory[29346] <=  8'h00;      memory[29347] <=  8'h00;      memory[29348] <=  8'h00;      memory[29349] <=  8'h00;      memory[29350] <=  8'h00;      memory[29351] <=  8'h00;      memory[29352] <=  8'h00;      memory[29353] <=  8'h00;      memory[29354] <=  8'h00;      memory[29355] <=  8'h00;      memory[29356] <=  8'h00;      memory[29357] <=  8'h00;      memory[29358] <=  8'h00;      memory[29359] <=  8'h00;      memory[29360] <=  8'h00;      memory[29361] <=  8'h00;      memory[29362] <=  8'h00;      memory[29363] <=  8'h00;      memory[29364] <=  8'h00;      memory[29365] <=  8'h00;      memory[29366] <=  8'h00;      memory[29367] <=  8'h00;      memory[29368] <=  8'h00;      memory[29369] <=  8'h00;      memory[29370] <=  8'h00;      memory[29371] <=  8'h00;      memory[29372] <=  8'h00;      memory[29373] <=  8'h00;      memory[29374] <=  8'h00;      memory[29375] <=  8'h00;      memory[29376] <=  8'h00;      memory[29377] <=  8'h00;      memory[29378] <=  8'h00;      memory[29379] <=  8'h00;      memory[29380] <=  8'h00;      memory[29381] <=  8'h00;      memory[29382] <=  8'h00;      memory[29383] <=  8'h00;      memory[29384] <=  8'h00;      memory[29385] <=  8'h00;      memory[29386] <=  8'h00;      memory[29387] <=  8'h00;      memory[29388] <=  8'h00;      memory[29389] <=  8'h00;      memory[29390] <=  8'h00;      memory[29391] <=  8'h00;      memory[29392] <=  8'h00;      memory[29393] <=  8'h00;      memory[29394] <=  8'h00;      memory[29395] <=  8'h00;      memory[29396] <=  8'h00;      memory[29397] <=  8'h00;      memory[29398] <=  8'h00;      memory[29399] <=  8'h00;      memory[29400] <=  8'h00;      memory[29401] <=  8'h00;      memory[29402] <=  8'h00;      memory[29403] <=  8'h00;      memory[29404] <=  8'h00;      memory[29405] <=  8'h00;      memory[29406] <=  8'h00;      memory[29407] <=  8'h00;      memory[29408] <=  8'h00;      memory[29409] <=  8'h00;      memory[29410] <=  8'h00;      memory[29411] <=  8'h00;      memory[29412] <=  8'h00;      memory[29413] <=  8'h00;      memory[29414] <=  8'h00;      memory[29415] <=  8'h00;      memory[29416] <=  8'h00;      memory[29417] <=  8'h00;      memory[29418] <=  8'h00;      memory[29419] <=  8'h00;      memory[29420] <=  8'h00;      memory[29421] <=  8'h00;      memory[29422] <=  8'h00;      memory[29423] <=  8'h00;      memory[29424] <=  8'h00;      memory[29425] <=  8'h00;      memory[29426] <=  8'h00;      memory[29427] <=  8'h00;      memory[29428] <=  8'h00;      memory[29429] <=  8'h00;      memory[29430] <=  8'h00;      memory[29431] <=  8'h00;      memory[29432] <=  8'h00;      memory[29433] <=  8'h00;      memory[29434] <=  8'h00;      memory[29435] <=  8'h00;      memory[29436] <=  8'h00;      memory[29437] <=  8'h00;      memory[29438] <=  8'h00;      memory[29439] <=  8'h00;      memory[29440] <=  8'h00;      memory[29441] <=  8'h00;      memory[29442] <=  8'h00;      memory[29443] <=  8'h00;      memory[29444] <=  8'h00;      memory[29445] <=  8'h00;      memory[29446] <=  8'h00;      memory[29447] <=  8'h00;      memory[29448] <=  8'h00;      memory[29449] <=  8'h00;      memory[29450] <=  8'h00;      memory[29451] <=  8'h00;      memory[29452] <=  8'h00;      memory[29453] <=  8'h00;      memory[29454] <=  8'h00;      memory[29455] <=  8'h00;      memory[29456] <=  8'h00;      memory[29457] <=  8'h00;      memory[29458] <=  8'h00;      memory[29459] <=  8'h00;      memory[29460] <=  8'h00;      memory[29461] <=  8'h00;      memory[29462] <=  8'h00;      memory[29463] <=  8'h00;      memory[29464] <=  8'h00;      memory[29465] <=  8'h00;      memory[29466] <=  8'h00;      memory[29467] <=  8'h00;      memory[29468] <=  8'h00;      memory[29469] <=  8'h00;      memory[29470] <=  8'h00;      memory[29471] <=  8'h00;      memory[29472] <=  8'h00;      memory[29473] <=  8'h00;      memory[29474] <=  8'h00;      memory[29475] <=  8'h00;      memory[29476] <=  8'h00;      memory[29477] <=  8'h00;      memory[29478] <=  8'h00;      memory[29479] <=  8'h00;      memory[29480] <=  8'h00;      memory[29481] <=  8'h00;      memory[29482] <=  8'h00;      memory[29483] <=  8'h00;      memory[29484] <=  8'h00;      memory[29485] <=  8'h00;      memory[29486] <=  8'h00;      memory[29487] <=  8'h00;      memory[29488] <=  8'h00;      memory[29489] <=  8'h00;      memory[29490] <=  8'h00;      memory[29491] <=  8'h00;      memory[29492] <=  8'h00;      memory[29493] <=  8'h00;      memory[29494] <=  8'h00;      memory[29495] <=  8'h00;      memory[29496] <=  8'h00;      memory[29497] <=  8'h00;      memory[29498] <=  8'h00;      memory[29499] <=  8'h00;      memory[29500] <=  8'h00;      memory[29501] <=  8'h00;      memory[29502] <=  8'h00;      memory[29503] <=  8'h00;      memory[29504] <=  8'h00;      memory[29505] <=  8'h00;      memory[29506] <=  8'h00;      memory[29507] <=  8'h00;      memory[29508] <=  8'h00;      memory[29509] <=  8'h00;      memory[29510] <=  8'h00;      memory[29511] <=  8'h00;      memory[29512] <=  8'h00;      memory[29513] <=  8'h00;      memory[29514] <=  8'h00;      memory[29515] <=  8'h00;      memory[29516] <=  8'h00;      memory[29517] <=  8'h00;      memory[29518] <=  8'h00;      memory[29519] <=  8'h00;      memory[29520] <=  8'h00;      memory[29521] <=  8'h00;      memory[29522] <=  8'h00;      memory[29523] <=  8'h00;      memory[29524] <=  8'h00;      memory[29525] <=  8'h00;      memory[29526] <=  8'h00;      memory[29527] <=  8'h00;      memory[29528] <=  8'h00;      memory[29529] <=  8'h00;      memory[29530] <=  8'h00;      memory[29531] <=  8'h00;      memory[29532] <=  8'h00;      memory[29533] <=  8'h00;      memory[29534] <=  8'h00;      memory[29535] <=  8'h00;      memory[29536] <=  8'h00;      memory[29537] <=  8'h00;      memory[29538] <=  8'h00;      memory[29539] <=  8'h00;      memory[29540] <=  8'h00;      memory[29541] <=  8'h00;      memory[29542] <=  8'h00;      memory[29543] <=  8'h00;      memory[29544] <=  8'h00;      memory[29545] <=  8'h00;      memory[29546] <=  8'h00;      memory[29547] <=  8'h00;      memory[29548] <=  8'h00;      memory[29549] <=  8'h00;      memory[29550] <=  8'h00;      memory[29551] <=  8'h00;      memory[29552] <=  8'h00;      memory[29553] <=  8'h00;      memory[29554] <=  8'h00;      memory[29555] <=  8'h00;      memory[29556] <=  8'h00;      memory[29557] <=  8'h00;      memory[29558] <=  8'h00;      memory[29559] <=  8'h00;      memory[29560] <=  8'h00;      memory[29561] <=  8'h00;      memory[29562] <=  8'h00;      memory[29563] <=  8'h00;      memory[29564] <=  8'h00;      memory[29565] <=  8'h00;      memory[29566] <=  8'h00;      memory[29567] <=  8'h00;      memory[29568] <=  8'h00;      memory[29569] <=  8'h00;      memory[29570] <=  8'h00;      memory[29571] <=  8'h00;      memory[29572] <=  8'h00;      memory[29573] <=  8'h00;      memory[29574] <=  8'h00;      memory[29575] <=  8'h00;      memory[29576] <=  8'h00;      memory[29577] <=  8'h00;      memory[29578] <=  8'h00;      memory[29579] <=  8'h00;      memory[29580] <=  8'h00;      memory[29581] <=  8'h00;      memory[29582] <=  8'h00;      memory[29583] <=  8'h00;      memory[29584] <=  8'h00;      memory[29585] <=  8'h00;      memory[29586] <=  8'h00;      memory[29587] <=  8'h00;      memory[29588] <=  8'h00;      memory[29589] <=  8'h00;      memory[29590] <=  8'h00;      memory[29591] <=  8'h00;      memory[29592] <=  8'h00;      memory[29593] <=  8'h00;      memory[29594] <=  8'h00;      memory[29595] <=  8'h00;      memory[29596] <=  8'h00;      memory[29597] <=  8'h00;      memory[29598] <=  8'h00;      memory[29599] <=  8'h00;      memory[29600] <=  8'h00;      memory[29601] <=  8'h00;      memory[29602] <=  8'h00;      memory[29603] <=  8'h00;      memory[29604] <=  8'h00;      memory[29605] <=  8'h00;      memory[29606] <=  8'h00;      memory[29607] <=  8'h00;      memory[29608] <=  8'h00;      memory[29609] <=  8'h00;      memory[29610] <=  8'h00;      memory[29611] <=  8'h00;      memory[29612] <=  8'h00;      memory[29613] <=  8'h00;      memory[29614] <=  8'h00;      memory[29615] <=  8'h00;      memory[29616] <=  8'h00;      memory[29617] <=  8'h00;      memory[29618] <=  8'h00;      memory[29619] <=  8'h00;      memory[29620] <=  8'h00;      memory[29621] <=  8'h00;      memory[29622] <=  8'h00;      memory[29623] <=  8'h00;      memory[29624] <=  8'h00;      memory[29625] <=  8'h00;      memory[29626] <=  8'h00;      memory[29627] <=  8'h00;      memory[29628] <=  8'h00;      memory[29629] <=  8'h00;      memory[29630] <=  8'h00;      memory[29631] <=  8'h00;      memory[29632] <=  8'h00;      memory[29633] <=  8'h00;      memory[29634] <=  8'h00;      memory[29635] <=  8'h00;      memory[29636] <=  8'h00;      memory[29637] <=  8'h00;      memory[29638] <=  8'h00;      memory[29639] <=  8'h00;      memory[29640] <=  8'h00;      memory[29641] <=  8'h00;      memory[29642] <=  8'h00;      memory[29643] <=  8'h00;      memory[29644] <=  8'h00;      memory[29645] <=  8'h00;      memory[29646] <=  8'h00;      memory[29647] <=  8'h00;      memory[29648] <=  8'h00;      memory[29649] <=  8'h00;      memory[29650] <=  8'h00;      memory[29651] <=  8'h00;      memory[29652] <=  8'h00;      memory[29653] <=  8'h00;      memory[29654] <=  8'h00;      memory[29655] <=  8'h00;      memory[29656] <=  8'h00;      memory[29657] <=  8'h00;      memory[29658] <=  8'h00;      memory[29659] <=  8'h00;      memory[29660] <=  8'h00;      memory[29661] <=  8'h00;      memory[29662] <=  8'h00;      memory[29663] <=  8'h00;      memory[29664] <=  8'h00;      memory[29665] <=  8'h00;      memory[29666] <=  8'h00;      memory[29667] <=  8'h00;      memory[29668] <=  8'h00;      memory[29669] <=  8'h00;      memory[29670] <=  8'h00;      memory[29671] <=  8'h00;      memory[29672] <=  8'h00;      memory[29673] <=  8'h00;      memory[29674] <=  8'h00;      memory[29675] <=  8'h00;      memory[29676] <=  8'h00;      memory[29677] <=  8'h00;      memory[29678] <=  8'h00;      memory[29679] <=  8'h00;      memory[29680] <=  8'h00;      memory[29681] <=  8'h00;      memory[29682] <=  8'h00;      memory[29683] <=  8'h00;      memory[29684] <=  8'h00;      memory[29685] <=  8'h00;      memory[29686] <=  8'h00;      memory[29687] <=  8'h00;      memory[29688] <=  8'h00;      memory[29689] <=  8'h00;      memory[29690] <=  8'h00;      memory[29691] <=  8'h00;      memory[29692] <=  8'h00;      memory[29693] <=  8'h00;      memory[29694] <=  8'h00;      memory[29695] <=  8'h00;      memory[29696] <=  8'h00;      memory[29697] <=  8'h00;      memory[29698] <=  8'h00;      memory[29699] <=  8'h00;      memory[29700] <=  8'h00;      memory[29701] <=  8'h00;      memory[29702] <=  8'h00;      memory[29703] <=  8'h00;      memory[29704] <=  8'h00;      memory[29705] <=  8'h00;      memory[29706] <=  8'h00;      memory[29707] <=  8'h00;      memory[29708] <=  8'h00;      memory[29709] <=  8'h00;      memory[29710] <=  8'h00;      memory[29711] <=  8'h00;      memory[29712] <=  8'h00;      memory[29713] <=  8'h00;      memory[29714] <=  8'h00;      memory[29715] <=  8'h00;      memory[29716] <=  8'h00;      memory[29717] <=  8'h00;      memory[29718] <=  8'h00;      memory[29719] <=  8'h00;      memory[29720] <=  8'h00;      memory[29721] <=  8'h00;      memory[29722] <=  8'h00;      memory[29723] <=  8'h00;      memory[29724] <=  8'h00;      memory[29725] <=  8'h00;      memory[29726] <=  8'h00;      memory[29727] <=  8'h00;      memory[29728] <=  8'h00;      memory[29729] <=  8'h00;      memory[29730] <=  8'h00;      memory[29731] <=  8'h00;      memory[29732] <=  8'h00;      memory[29733] <=  8'h00;      memory[29734] <=  8'h00;      memory[29735] <=  8'h00;      memory[29736] <=  8'h00;      memory[29737] <=  8'h00;      memory[29738] <=  8'h00;      memory[29739] <=  8'h00;      memory[29740] <=  8'h00;      memory[29741] <=  8'h00;      memory[29742] <=  8'h00;      memory[29743] <=  8'h00;      memory[29744] <=  8'h00;      memory[29745] <=  8'h00;      memory[29746] <=  8'h00;      memory[29747] <=  8'h00;      memory[29748] <=  8'h00;      memory[29749] <=  8'h00;      memory[29750] <=  8'h00;      memory[29751] <=  8'h00;      memory[29752] <=  8'h00;      memory[29753] <=  8'h00;      memory[29754] <=  8'h00;      memory[29755] <=  8'h00;      memory[29756] <=  8'h00;      memory[29757] <=  8'h00;      memory[29758] <=  8'h00;      memory[29759] <=  8'h00;      memory[29760] <=  8'h00;      memory[29761] <=  8'h00;      memory[29762] <=  8'h00;      memory[29763] <=  8'h00;      memory[29764] <=  8'h00;      memory[29765] <=  8'h00;      memory[29766] <=  8'h00;      memory[29767] <=  8'h00;      memory[29768] <=  8'h00;      memory[29769] <=  8'h00;      memory[29770] <=  8'h00;      memory[29771] <=  8'h00;      memory[29772] <=  8'h00;      memory[29773] <=  8'h00;      memory[29774] <=  8'h00;      memory[29775] <=  8'h00;      memory[29776] <=  8'h00;      memory[29777] <=  8'h00;      memory[29778] <=  8'h00;      memory[29779] <=  8'h00;      memory[29780] <=  8'h00;      memory[29781] <=  8'h00;      memory[29782] <=  8'h00;      memory[29783] <=  8'h00;      memory[29784] <=  8'h00;      memory[29785] <=  8'h00;      memory[29786] <=  8'h00;      memory[29787] <=  8'h00;      memory[29788] <=  8'h00;      memory[29789] <=  8'h00;      memory[29790] <=  8'h00;      memory[29791] <=  8'h00;      memory[29792] <=  8'h00;      memory[29793] <=  8'h00;      memory[29794] <=  8'h00;      memory[29795] <=  8'h00;      memory[29796] <=  8'h00;      memory[29797] <=  8'h00;      memory[29798] <=  8'h00;      memory[29799] <=  8'h00;      memory[29800] <=  8'h00;      memory[29801] <=  8'h00;      memory[29802] <=  8'h00;      memory[29803] <=  8'h00;      memory[29804] <=  8'h00;      memory[29805] <=  8'h00;      memory[29806] <=  8'h00;      memory[29807] <=  8'h00;      memory[29808] <=  8'h00;      memory[29809] <=  8'h00;      memory[29810] <=  8'h00;      memory[29811] <=  8'h00;      memory[29812] <=  8'h00;      memory[29813] <=  8'h00;      memory[29814] <=  8'h00;      memory[29815] <=  8'h00;      memory[29816] <=  8'h00;      memory[29817] <=  8'h00;      memory[29818] <=  8'h00;      memory[29819] <=  8'h00;      memory[29820] <=  8'h00;      memory[29821] <=  8'h00;      memory[29822] <=  8'h00;      memory[29823] <=  8'h00;      memory[29824] <=  8'h00;      memory[29825] <=  8'h00;      memory[29826] <=  8'h00;      memory[29827] <=  8'h00;      memory[29828] <=  8'h00;      memory[29829] <=  8'h00;      memory[29830] <=  8'h00;      memory[29831] <=  8'h00;      memory[29832] <=  8'h00;      memory[29833] <=  8'h00;      memory[29834] <=  8'h00;      memory[29835] <=  8'h00;      memory[29836] <=  8'h00;      memory[29837] <=  8'h00;      memory[29838] <=  8'h00;      memory[29839] <=  8'h00;      memory[29840] <=  8'h00;      memory[29841] <=  8'h00;      memory[29842] <=  8'h00;      memory[29843] <=  8'h00;      memory[29844] <=  8'h00;      memory[29845] <=  8'h00;      memory[29846] <=  8'h00;      memory[29847] <=  8'h00;      memory[29848] <=  8'h00;      memory[29849] <=  8'h00;      memory[29850] <=  8'h00;      memory[29851] <=  8'h00;      memory[29852] <=  8'h00;      memory[29853] <=  8'h00;      memory[29854] <=  8'h00;      memory[29855] <=  8'h00;      memory[29856] <=  8'h00;      memory[29857] <=  8'h00;      memory[29858] <=  8'h00;      memory[29859] <=  8'h00;      memory[29860] <=  8'h00;      memory[29861] <=  8'h00;      memory[29862] <=  8'h00;      memory[29863] <=  8'h00;      memory[29864] <=  8'h00;      memory[29865] <=  8'h00;      memory[29866] <=  8'h00;      memory[29867] <=  8'h00;      memory[29868] <=  8'h00;      memory[29869] <=  8'h00;      memory[29870] <=  8'h00;      memory[29871] <=  8'h00;      memory[29872] <=  8'h00;      memory[29873] <=  8'h00;      memory[29874] <=  8'h00;      memory[29875] <=  8'h00;      memory[29876] <=  8'h00;      memory[29877] <=  8'h00;      memory[29878] <=  8'h00;      memory[29879] <=  8'h00;      memory[29880] <=  8'h00;      memory[29881] <=  8'h00;      memory[29882] <=  8'h00;      memory[29883] <=  8'h00;      memory[29884] <=  8'h00;      memory[29885] <=  8'h00;      memory[29886] <=  8'h00;      memory[29887] <=  8'h00;      memory[29888] <=  8'h00;      memory[29889] <=  8'h00;      memory[29890] <=  8'h00;      memory[29891] <=  8'h00;      memory[29892] <=  8'h00;      memory[29893] <=  8'h00;      memory[29894] <=  8'h00;      memory[29895] <=  8'h00;      memory[29896] <=  8'h00;      memory[29897] <=  8'h00;      memory[29898] <=  8'h00;      memory[29899] <=  8'h00;      memory[29900] <=  8'h00;      memory[29901] <=  8'h00;      memory[29902] <=  8'h00;      memory[29903] <=  8'h00;      memory[29904] <=  8'h00;      memory[29905] <=  8'h00;      memory[29906] <=  8'h00;      memory[29907] <=  8'h00;      memory[29908] <=  8'h00;      memory[29909] <=  8'h00;      memory[29910] <=  8'h00;      memory[29911] <=  8'h00;      memory[29912] <=  8'h00;      memory[29913] <=  8'h00;      memory[29914] <=  8'h00;      memory[29915] <=  8'h00;      memory[29916] <=  8'h00;      memory[29917] <=  8'h00;      memory[29918] <=  8'h00;      memory[29919] <=  8'h00;      memory[29920] <=  8'h00;      memory[29921] <=  8'h00;      memory[29922] <=  8'h00;      memory[29923] <=  8'h00;      memory[29924] <=  8'h00;      memory[29925] <=  8'h00;      memory[29926] <=  8'h00;      memory[29927] <=  8'h00;      memory[29928] <=  8'h00;      memory[29929] <=  8'h00;      memory[29930] <=  8'h00;      memory[29931] <=  8'h00;      memory[29932] <=  8'h00;      memory[29933] <=  8'h00;      memory[29934] <=  8'h00;      memory[29935] <=  8'h00;      memory[29936] <=  8'h00;      memory[29937] <=  8'h00;      memory[29938] <=  8'h00;      memory[29939] <=  8'h00;      memory[29940] <=  8'h00;      memory[29941] <=  8'h00;      memory[29942] <=  8'h00;      memory[29943] <=  8'h00;      memory[29944] <=  8'h00;      memory[29945] <=  8'h00;      memory[29946] <=  8'h00;      memory[29947] <=  8'h00;      memory[29948] <=  8'h00;      memory[29949] <=  8'h00;      memory[29950] <=  8'h00;      memory[29951] <=  8'h00;      memory[29952] <=  8'h00;      memory[29953] <=  8'h00;      memory[29954] <=  8'h00;      memory[29955] <=  8'h00;      memory[29956] <=  8'h00;      memory[29957] <=  8'h00;      memory[29958] <=  8'h00;      memory[29959] <=  8'h00;      memory[29960] <=  8'h00;      memory[29961] <=  8'h00;      memory[29962] <=  8'h00;      memory[29963] <=  8'h00;      memory[29964] <=  8'h00;      memory[29965] <=  8'h00;      memory[29966] <=  8'h00;      memory[29967] <=  8'h00;      memory[29968] <=  8'h00;      memory[29969] <=  8'h00;      memory[29970] <=  8'h00;      memory[29971] <=  8'h00;      memory[29972] <=  8'h00;      memory[29973] <=  8'h00;      memory[29974] <=  8'h00;      memory[29975] <=  8'h00;      memory[29976] <=  8'h00;      memory[29977] <=  8'h00;      memory[29978] <=  8'h00;      memory[29979] <=  8'h00;      memory[29980] <=  8'h00;      memory[29981] <=  8'h00;      memory[29982] <=  8'h00;      memory[29983] <=  8'h00;      memory[29984] <=  8'h00;      memory[29985] <=  8'h00;      memory[29986] <=  8'h00;      memory[29987] <=  8'h00;      memory[29988] <=  8'h00;      memory[29989] <=  8'h00;      memory[29990] <=  8'h00;      memory[29991] <=  8'h00;      memory[29992] <=  8'h00;      memory[29993] <=  8'h00;      memory[29994] <=  8'h00;      memory[29995] <=  8'h00;      memory[29996] <=  8'h00;      memory[29997] <=  8'h00;      memory[29998] <=  8'h00;      memory[29999] <=  8'h00;      memory[30000] <=  8'h00;      memory[30001] <=  8'h00;      memory[30002] <=  8'h00;      memory[30003] <=  8'h00;      memory[30004] <=  8'h00;      memory[30005] <=  8'h00;      memory[30006] <=  8'h00;      memory[30007] <=  8'h00;      memory[30008] <=  8'h00;      memory[30009] <=  8'h00;      memory[30010] <=  8'h00;      memory[30011] <=  8'h00;      memory[30012] <=  8'h00;      memory[30013] <=  8'h00;      memory[30014] <=  8'h00;      memory[30015] <=  8'h00;      memory[30016] <=  8'h00;      memory[30017] <=  8'h00;      memory[30018] <=  8'h00;      memory[30019] <=  8'h00;      memory[30020] <=  8'h00;      memory[30021] <=  8'h00;      memory[30022] <=  8'h00;      memory[30023] <=  8'h00;      memory[30024] <=  8'h00;      memory[30025] <=  8'h00;      memory[30026] <=  8'h00;      memory[30027] <=  8'h00;      memory[30028] <=  8'h00;      memory[30029] <=  8'h00;      memory[30030] <=  8'h00;      memory[30031] <=  8'h00;      memory[30032] <=  8'h00;      memory[30033] <=  8'h00;      memory[30034] <=  8'h00;      memory[30035] <=  8'h00;      memory[30036] <=  8'h00;      memory[30037] <=  8'h00;      memory[30038] <=  8'h00;      memory[30039] <=  8'h00;      memory[30040] <=  8'h00;      memory[30041] <=  8'h00;      memory[30042] <=  8'h00;      memory[30043] <=  8'h00;      memory[30044] <=  8'h00;      memory[30045] <=  8'h00;      memory[30046] <=  8'h00;      memory[30047] <=  8'h00;      memory[30048] <=  8'h00;      memory[30049] <=  8'h00;      memory[30050] <=  8'h00;      memory[30051] <=  8'h00;      memory[30052] <=  8'h00;      memory[30053] <=  8'h00;      memory[30054] <=  8'h00;      memory[30055] <=  8'h00;      memory[30056] <=  8'h00;      memory[30057] <=  8'h00;      memory[30058] <=  8'h00;      memory[30059] <=  8'h00;      memory[30060] <=  8'h00;      memory[30061] <=  8'h00;      memory[30062] <=  8'h00;      memory[30063] <=  8'h00;      memory[30064] <=  8'h00;      memory[30065] <=  8'h00;      memory[30066] <=  8'h00;      memory[30067] <=  8'h00;      memory[30068] <=  8'h00;      memory[30069] <=  8'h00;      memory[30070] <=  8'h00;      memory[30071] <=  8'h00;      memory[30072] <=  8'h00;      memory[30073] <=  8'h00;      memory[30074] <=  8'h00;      memory[30075] <=  8'h00;      memory[30076] <=  8'h00;      memory[30077] <=  8'h00;      memory[30078] <=  8'h00;      memory[30079] <=  8'h00;      memory[30080] <=  8'h00;      memory[30081] <=  8'h00;      memory[30082] <=  8'h00;      memory[30083] <=  8'h00;      memory[30084] <=  8'h00;      memory[30085] <=  8'h00;      memory[30086] <=  8'h00;      memory[30087] <=  8'h00;      memory[30088] <=  8'h00;      memory[30089] <=  8'h00;      memory[30090] <=  8'h00;      memory[30091] <=  8'h00;      memory[30092] <=  8'h00;      memory[30093] <=  8'h00;      memory[30094] <=  8'h00;      memory[30095] <=  8'h00;      memory[30096] <=  8'h00;      memory[30097] <=  8'h00;      memory[30098] <=  8'h00;      memory[30099] <=  8'h00;      memory[30100] <=  8'h00;      memory[30101] <=  8'h00;      memory[30102] <=  8'h00;      memory[30103] <=  8'h00;      memory[30104] <=  8'h00;      memory[30105] <=  8'h00;      memory[30106] <=  8'h00;      memory[30107] <=  8'h00;      memory[30108] <=  8'h00;      memory[30109] <=  8'h00;      memory[30110] <=  8'h00;      memory[30111] <=  8'h00;      memory[30112] <=  8'h00;      memory[30113] <=  8'h00;      memory[30114] <=  8'h00;      memory[30115] <=  8'h00;      memory[30116] <=  8'h00;      memory[30117] <=  8'h00;      memory[30118] <=  8'h00;      memory[30119] <=  8'h00;      memory[30120] <=  8'h00;      memory[30121] <=  8'h00;      memory[30122] <=  8'h00;      memory[30123] <=  8'h00;      memory[30124] <=  8'h00;      memory[30125] <=  8'h00;      memory[30126] <=  8'h00;      memory[30127] <=  8'h00;      memory[30128] <=  8'h00;      memory[30129] <=  8'h00;      memory[30130] <=  8'h00;      memory[30131] <=  8'h00;      memory[30132] <=  8'h00;      memory[30133] <=  8'h00;      memory[30134] <=  8'h00;      memory[30135] <=  8'h00;      memory[30136] <=  8'h00;      memory[30137] <=  8'h00;      memory[30138] <=  8'h00;      memory[30139] <=  8'h00;      memory[30140] <=  8'h00;      memory[30141] <=  8'h00;      memory[30142] <=  8'h00;      memory[30143] <=  8'h00;      memory[30144] <=  8'h00;      memory[30145] <=  8'h00;      memory[30146] <=  8'h00;      memory[30147] <=  8'h00;      memory[30148] <=  8'h00;      memory[30149] <=  8'h00;      memory[30150] <=  8'h00;      memory[30151] <=  8'h00;      memory[30152] <=  8'h00;      memory[30153] <=  8'h00;      memory[30154] <=  8'h00;      memory[30155] <=  8'h00;      memory[30156] <=  8'h00;      memory[30157] <=  8'h00;      memory[30158] <=  8'h00;      memory[30159] <=  8'h00;      memory[30160] <=  8'h00;      memory[30161] <=  8'h00;      memory[30162] <=  8'h00;      memory[30163] <=  8'h00;      memory[30164] <=  8'h00;      memory[30165] <=  8'h00;      memory[30166] <=  8'h00;      memory[30167] <=  8'h00;      memory[30168] <=  8'h00;      memory[30169] <=  8'h00;      memory[30170] <=  8'h00;      memory[30171] <=  8'h00;      memory[30172] <=  8'h00;      memory[30173] <=  8'h00;      memory[30174] <=  8'h00;      memory[30175] <=  8'h00;      memory[30176] <=  8'h00;      memory[30177] <=  8'h00;      memory[30178] <=  8'h00;      memory[30179] <=  8'h00;      memory[30180] <=  8'h00;      memory[30181] <=  8'h00;      memory[30182] <=  8'h00;      memory[30183] <=  8'h00;      memory[30184] <=  8'h00;      memory[30185] <=  8'h00;      memory[30186] <=  8'h00;      memory[30187] <=  8'h00;      memory[30188] <=  8'h00;      memory[30189] <=  8'h00;      memory[30190] <=  8'h00;      memory[30191] <=  8'h00;      memory[30192] <=  8'h00;      memory[30193] <=  8'h00;      memory[30194] <=  8'h00;      memory[30195] <=  8'h00;      memory[30196] <=  8'h00;      memory[30197] <=  8'h00;      memory[30198] <=  8'h00;      memory[30199] <=  8'h00;      memory[30200] <=  8'h00;      memory[30201] <=  8'h00;      memory[30202] <=  8'h00;      memory[30203] <=  8'h00;      memory[30204] <=  8'h00;      memory[30205] <=  8'h00;      memory[30206] <=  8'h00;      memory[30207] <=  8'h00;      memory[30208] <=  8'h00;      memory[30209] <=  8'h00;      memory[30210] <=  8'h00;      memory[30211] <=  8'h00;      memory[30212] <=  8'h00;      memory[30213] <=  8'h00;      memory[30214] <=  8'h00;      memory[30215] <=  8'h00;      memory[30216] <=  8'h00;      memory[30217] <=  8'h00;      memory[30218] <=  8'h00;      memory[30219] <=  8'h00;      memory[30220] <=  8'h00;      memory[30221] <=  8'h00;      memory[30222] <=  8'h00;      memory[30223] <=  8'h00;      memory[30224] <=  8'h00;      memory[30225] <=  8'h00;      memory[30226] <=  8'h00;      memory[30227] <=  8'h00;      memory[30228] <=  8'h00;      memory[30229] <=  8'h00;      memory[30230] <=  8'h00;      memory[30231] <=  8'h00;      memory[30232] <=  8'h00;      memory[30233] <=  8'h00;      memory[30234] <=  8'h00;      memory[30235] <=  8'h00;      memory[30236] <=  8'h00;      memory[30237] <=  8'h00;      memory[30238] <=  8'h00;      memory[30239] <=  8'h00;      memory[30240] <=  8'h00;      memory[30241] <=  8'h00;      memory[30242] <=  8'h00;      memory[30243] <=  8'h00;      memory[30244] <=  8'h00;      memory[30245] <=  8'h00;      memory[30246] <=  8'h00;      memory[30247] <=  8'h00;      memory[30248] <=  8'h00;      memory[30249] <=  8'h00;      memory[30250] <=  8'h00;      memory[30251] <=  8'h00;      memory[30252] <=  8'h00;      memory[30253] <=  8'h00;      memory[30254] <=  8'h00;      memory[30255] <=  8'h00;      memory[30256] <=  8'h00;      memory[30257] <=  8'h00;      memory[30258] <=  8'h00;      memory[30259] <=  8'h00;      memory[30260] <=  8'h00;      memory[30261] <=  8'h00;      memory[30262] <=  8'h00;      memory[30263] <=  8'h00;      memory[30264] <=  8'h00;      memory[30265] <=  8'h00;      memory[30266] <=  8'h00;      memory[30267] <=  8'h00;      memory[30268] <=  8'h00;      memory[30269] <=  8'h00;      memory[30270] <=  8'h00;      memory[30271] <=  8'h00;      memory[30272] <=  8'h00;      memory[30273] <=  8'h00;      memory[30274] <=  8'h00;      memory[30275] <=  8'h00;      memory[30276] <=  8'h00;      memory[30277] <=  8'h00;      memory[30278] <=  8'h00;      memory[30279] <=  8'h00;      memory[30280] <=  8'h00;      memory[30281] <=  8'h00;      memory[30282] <=  8'h00;      memory[30283] <=  8'h00;      memory[30284] <=  8'h00;      memory[30285] <=  8'h00;      memory[30286] <=  8'h00;      memory[30287] <=  8'h00;      memory[30288] <=  8'h00;      memory[30289] <=  8'h00;      memory[30290] <=  8'h00;      memory[30291] <=  8'h00;      memory[30292] <=  8'h00;      memory[30293] <=  8'h00;      memory[30294] <=  8'h00;      memory[30295] <=  8'h00;      memory[30296] <=  8'h00;      memory[30297] <=  8'h00;      memory[30298] <=  8'h00;      memory[30299] <=  8'h00;      memory[30300] <=  8'h00;      memory[30301] <=  8'h00;      memory[30302] <=  8'h00;      memory[30303] <=  8'h00;      memory[30304] <=  8'h00;      memory[30305] <=  8'h00;      memory[30306] <=  8'h00;      memory[30307] <=  8'h00;      memory[30308] <=  8'h00;      memory[30309] <=  8'h00;      memory[30310] <=  8'h00;      memory[30311] <=  8'h00;      memory[30312] <=  8'h00;      memory[30313] <=  8'h00;      memory[30314] <=  8'h00;      memory[30315] <=  8'h00;      memory[30316] <=  8'h00;      memory[30317] <=  8'h00;      memory[30318] <=  8'h00;      memory[30319] <=  8'h00;      memory[30320] <=  8'h00;      memory[30321] <=  8'h00;      memory[30322] <=  8'h00;      memory[30323] <=  8'h00;      memory[30324] <=  8'h00;      memory[30325] <=  8'h00;      memory[30326] <=  8'h00;      memory[30327] <=  8'h00;      memory[30328] <=  8'h00;      memory[30329] <=  8'h00;      memory[30330] <=  8'h00;      memory[30331] <=  8'h00;      memory[30332] <=  8'h00;      memory[30333] <=  8'h00;      memory[30334] <=  8'h00;      memory[30335] <=  8'h00;      memory[30336] <=  8'h00;      memory[30337] <=  8'h00;      memory[30338] <=  8'h00;      memory[30339] <=  8'h00;      memory[30340] <=  8'h00;      memory[30341] <=  8'h00;      memory[30342] <=  8'h00;      memory[30343] <=  8'h00;      memory[30344] <=  8'h00;      memory[30345] <=  8'h00;      memory[30346] <=  8'h00;      memory[30347] <=  8'h00;      memory[30348] <=  8'h00;      memory[30349] <=  8'h00;      memory[30350] <=  8'h00;      memory[30351] <=  8'h00;      memory[30352] <=  8'h00;      memory[30353] <=  8'h00;      memory[30354] <=  8'h00;      memory[30355] <=  8'h00;      memory[30356] <=  8'h00;      memory[30357] <=  8'h00;      memory[30358] <=  8'h00;      memory[30359] <=  8'h00;      memory[30360] <=  8'h00;      memory[30361] <=  8'h00;      memory[30362] <=  8'h00;      memory[30363] <=  8'h00;      memory[30364] <=  8'h00;      memory[30365] <=  8'h00;      memory[30366] <=  8'h00;      memory[30367] <=  8'h00;      memory[30368] <=  8'h00;      memory[30369] <=  8'h00;      memory[30370] <=  8'h00;      memory[30371] <=  8'h00;      memory[30372] <=  8'h00;      memory[30373] <=  8'h00;      memory[30374] <=  8'h00;      memory[30375] <=  8'h00;      memory[30376] <=  8'h00;      memory[30377] <=  8'h00;      memory[30378] <=  8'h00;      memory[30379] <=  8'h00;      memory[30380] <=  8'h00;      memory[30381] <=  8'h00;      memory[30382] <=  8'h00;      memory[30383] <=  8'h00;      memory[30384] <=  8'h00;      memory[30385] <=  8'h00;      memory[30386] <=  8'h00;      memory[30387] <=  8'h00;      memory[30388] <=  8'h00;      memory[30389] <=  8'h00;      memory[30390] <=  8'h00;      memory[30391] <=  8'h00;      memory[30392] <=  8'h00;      memory[30393] <=  8'h00;      memory[30394] <=  8'h00;      memory[30395] <=  8'h00;      memory[30396] <=  8'h00;      memory[30397] <=  8'h00;      memory[30398] <=  8'h00;      memory[30399] <=  8'h00;      memory[30400] <=  8'h00;      memory[30401] <=  8'h00;      memory[30402] <=  8'h00;      memory[30403] <=  8'h00;      memory[30404] <=  8'h00;      memory[30405] <=  8'h00;      memory[30406] <=  8'h00;      memory[30407] <=  8'h00;      memory[30408] <=  8'h00;      memory[30409] <=  8'h00;      memory[30410] <=  8'h00;      memory[30411] <=  8'h00;      memory[30412] <=  8'h00;      memory[30413] <=  8'h00;      memory[30414] <=  8'h00;      memory[30415] <=  8'h00;      memory[30416] <=  8'h00;      memory[30417] <=  8'h00;      memory[30418] <=  8'h00;      memory[30419] <=  8'h00;      memory[30420] <=  8'h00;      memory[30421] <=  8'h00;      memory[30422] <=  8'h00;      memory[30423] <=  8'h00;      memory[30424] <=  8'h00;      memory[30425] <=  8'h00;      memory[30426] <=  8'h00;      memory[30427] <=  8'h00;      memory[30428] <=  8'h00;      memory[30429] <=  8'h00;      memory[30430] <=  8'h00;      memory[30431] <=  8'h00;      memory[30432] <=  8'h00;      memory[30433] <=  8'h00;      memory[30434] <=  8'h00;      memory[30435] <=  8'h00;      memory[30436] <=  8'h00;      memory[30437] <=  8'h00;      memory[30438] <=  8'h00;      memory[30439] <=  8'h00;      memory[30440] <=  8'h00;      memory[30441] <=  8'h00;      memory[30442] <=  8'h00;      memory[30443] <=  8'h00;      memory[30444] <=  8'h00;      memory[30445] <=  8'h00;      memory[30446] <=  8'h00;      memory[30447] <=  8'h00;      memory[30448] <=  8'h00;      memory[30449] <=  8'h00;      memory[30450] <=  8'h00;      memory[30451] <=  8'h00;      memory[30452] <=  8'h00;      memory[30453] <=  8'h00;      memory[30454] <=  8'h00;      memory[30455] <=  8'h00;      memory[30456] <=  8'h00;      memory[30457] <=  8'h00;      memory[30458] <=  8'h00;      memory[30459] <=  8'h00;      memory[30460] <=  8'h00;      memory[30461] <=  8'h00;      memory[30462] <=  8'h00;      memory[30463] <=  8'h00;      memory[30464] <=  8'h00;      memory[30465] <=  8'h00;      memory[30466] <=  8'h00;      memory[30467] <=  8'h00;      memory[30468] <=  8'h00;      memory[30469] <=  8'h00;      memory[30470] <=  8'h00;      memory[30471] <=  8'h00;      memory[30472] <=  8'h00;      memory[30473] <=  8'h00;      memory[30474] <=  8'h00;      memory[30475] <=  8'h00;      memory[30476] <=  8'h00;      memory[30477] <=  8'h00;      memory[30478] <=  8'h00;      memory[30479] <=  8'h00;      memory[30480] <=  8'h00;      memory[30481] <=  8'h00;      memory[30482] <=  8'h00;      memory[30483] <=  8'h00;      memory[30484] <=  8'h00;      memory[30485] <=  8'h00;      memory[30486] <=  8'h00;      memory[30487] <=  8'h00;      memory[30488] <=  8'h00;      memory[30489] <=  8'h00;      memory[30490] <=  8'h00;      memory[30491] <=  8'h00;      memory[30492] <=  8'h00;      memory[30493] <=  8'h00;      memory[30494] <=  8'h00;      memory[30495] <=  8'h00;      memory[30496] <=  8'h00;      memory[30497] <=  8'h00;      memory[30498] <=  8'h00;      memory[30499] <=  8'h00;      memory[30500] <=  8'h00;      memory[30501] <=  8'h00;      memory[30502] <=  8'h00;      memory[30503] <=  8'h00;      memory[30504] <=  8'h00;      memory[30505] <=  8'h00;      memory[30506] <=  8'h00;      memory[30507] <=  8'h00;      memory[30508] <=  8'h00;      memory[30509] <=  8'h00;      memory[30510] <=  8'h00;      memory[30511] <=  8'h00;      memory[30512] <=  8'h00;      memory[30513] <=  8'h00;      memory[30514] <=  8'h00;      memory[30515] <=  8'h00;      memory[30516] <=  8'h00;      memory[30517] <=  8'h00;      memory[30518] <=  8'h00;      memory[30519] <=  8'h00;      memory[30520] <=  8'h00;      memory[30521] <=  8'h00;      memory[30522] <=  8'h00;      memory[30523] <=  8'h00;      memory[30524] <=  8'h00;      memory[30525] <=  8'h00;      memory[30526] <=  8'h00;      memory[30527] <=  8'h00;      memory[30528] <=  8'h00;      memory[30529] <=  8'h00;      memory[30530] <=  8'h00;      memory[30531] <=  8'h00;      memory[30532] <=  8'h00;      memory[30533] <=  8'h00;      memory[30534] <=  8'h00;      memory[30535] <=  8'h00;      memory[30536] <=  8'h00;      memory[30537] <=  8'h00;      memory[30538] <=  8'h00;      memory[30539] <=  8'h00;      memory[30540] <=  8'h00;      memory[30541] <=  8'h00;      memory[30542] <=  8'h00;      memory[30543] <=  8'h00;      memory[30544] <=  8'h00;      memory[30545] <=  8'h00;      memory[30546] <=  8'h00;      memory[30547] <=  8'h00;      memory[30548] <=  8'h00;      memory[30549] <=  8'h00;      memory[30550] <=  8'h00;      memory[30551] <=  8'h00;      memory[30552] <=  8'h00;      memory[30553] <=  8'h00;      memory[30554] <=  8'h00;      memory[30555] <=  8'h00;      memory[30556] <=  8'h00;      memory[30557] <=  8'h00;      memory[30558] <=  8'h00;      memory[30559] <=  8'h00;      memory[30560] <=  8'h00;      memory[30561] <=  8'h00;      memory[30562] <=  8'h00;      memory[30563] <=  8'h00;      memory[30564] <=  8'h00;      memory[30565] <=  8'h00;      memory[30566] <=  8'h00;      memory[30567] <=  8'h00;      memory[30568] <=  8'h00;      memory[30569] <=  8'h00;      memory[30570] <=  8'h00;      memory[30571] <=  8'h00;      memory[30572] <=  8'h00;      memory[30573] <=  8'h00;      memory[30574] <=  8'h00;      memory[30575] <=  8'h00;      memory[30576] <=  8'h00;      memory[30577] <=  8'h00;      memory[30578] <=  8'h00;      memory[30579] <=  8'h00;      memory[30580] <=  8'h00;      memory[30581] <=  8'h00;      memory[30582] <=  8'h00;      memory[30583] <=  8'h00;      memory[30584] <=  8'h00;      memory[30585] <=  8'h00;      memory[30586] <=  8'h00;      memory[30587] <=  8'h00;      memory[30588] <=  8'h00;      memory[30589] <=  8'h00;      memory[30590] <=  8'h00;      memory[30591] <=  8'h00;      memory[30592] <=  8'h00;      memory[30593] <=  8'h00;      memory[30594] <=  8'h00;      memory[30595] <=  8'h00;      memory[30596] <=  8'h00;      memory[30597] <=  8'h00;      memory[30598] <=  8'h00;      memory[30599] <=  8'h00;      memory[30600] <=  8'h00;      memory[30601] <=  8'h00;      memory[30602] <=  8'h00;      memory[30603] <=  8'h00;      memory[30604] <=  8'h00;      memory[30605] <=  8'h00;      memory[30606] <=  8'h00;      memory[30607] <=  8'h00;      memory[30608] <=  8'h00;      memory[30609] <=  8'h00;      memory[30610] <=  8'h00;      memory[30611] <=  8'h00;      memory[30612] <=  8'h00;      memory[30613] <=  8'h00;      memory[30614] <=  8'h00;      memory[30615] <=  8'h00;      memory[30616] <=  8'h00;      memory[30617] <=  8'h00;      memory[30618] <=  8'h00;      memory[30619] <=  8'h00;      memory[30620] <=  8'h00;      memory[30621] <=  8'h00;      memory[30622] <=  8'h00;      memory[30623] <=  8'h00;      memory[30624] <=  8'h00;      memory[30625] <=  8'h00;      memory[30626] <=  8'h00;      memory[30627] <=  8'h00;      memory[30628] <=  8'h00;      memory[30629] <=  8'h00;      memory[30630] <=  8'h00;      memory[30631] <=  8'h00;      memory[30632] <=  8'h00;      memory[30633] <=  8'h00;      memory[30634] <=  8'h00;      memory[30635] <=  8'h00;      memory[30636] <=  8'h00;      memory[30637] <=  8'h00;      memory[30638] <=  8'h00;      memory[30639] <=  8'h00;      memory[30640] <=  8'h00;      memory[30641] <=  8'h00;      memory[30642] <=  8'h00;      memory[30643] <=  8'h00;      memory[30644] <=  8'h00;      memory[30645] <=  8'h00;      memory[30646] <=  8'h00;      memory[30647] <=  8'h00;      memory[30648] <=  8'h00;      memory[30649] <=  8'h00;      memory[30650] <=  8'h00;      memory[30651] <=  8'h00;      memory[30652] <=  8'h00;      memory[30653] <=  8'h00;      memory[30654] <=  8'h00;      memory[30655] <=  8'h00;      memory[30656] <=  8'h00;      memory[30657] <=  8'h00;      memory[30658] <=  8'h00;      memory[30659] <=  8'h00;      memory[30660] <=  8'h00;      memory[30661] <=  8'h00;      memory[30662] <=  8'h00;      memory[30663] <=  8'h00;      memory[30664] <=  8'h00;      memory[30665] <=  8'h00;      memory[30666] <=  8'h00;      memory[30667] <=  8'h00;      memory[30668] <=  8'h00;      memory[30669] <=  8'h00;      memory[30670] <=  8'h00;      memory[30671] <=  8'h00;      memory[30672] <=  8'h00;      memory[30673] <=  8'h00;      memory[30674] <=  8'h00;      memory[30675] <=  8'h00;      memory[30676] <=  8'h00;      memory[30677] <=  8'h00;      memory[30678] <=  8'h00;      memory[30679] <=  8'h00;      memory[30680] <=  8'h00;      memory[30681] <=  8'h00;      memory[30682] <=  8'h00;      memory[30683] <=  8'h00;      memory[30684] <=  8'h00;      memory[30685] <=  8'h00;      memory[30686] <=  8'h00;      memory[30687] <=  8'h00;      memory[30688] <=  8'h00;      memory[30689] <=  8'h00;      memory[30690] <=  8'h00;      memory[30691] <=  8'h00;      memory[30692] <=  8'h00;      memory[30693] <=  8'h00;      memory[30694] <=  8'h00;      memory[30695] <=  8'h00;      memory[30696] <=  8'h00;      memory[30697] <=  8'h00;      memory[30698] <=  8'h00;      memory[30699] <=  8'h00;      memory[30700] <=  8'h00;      memory[30701] <=  8'h00;      memory[30702] <=  8'h00;      memory[30703] <=  8'h00;      memory[30704] <=  8'h00;      memory[30705] <=  8'h00;      memory[30706] <=  8'h00;      memory[30707] <=  8'h00;      memory[30708] <=  8'h00;      memory[30709] <=  8'h00;      memory[30710] <=  8'h00;      memory[30711] <=  8'h00;      memory[30712] <=  8'h00;      memory[30713] <=  8'h00;      memory[30714] <=  8'h00;      memory[30715] <=  8'h00;      memory[30716] <=  8'h00;      memory[30717] <=  8'h00;      memory[30718] <=  8'h00;      memory[30719] <=  8'h00;      memory[30720] <=  8'h00;      memory[30721] <=  8'h00;      memory[30722] <=  8'h00;      memory[30723] <=  8'h00;      memory[30724] <=  8'h00;      memory[30725] <=  8'h00;      memory[30726] <=  8'h00;      memory[30727] <=  8'h00;      memory[30728] <=  8'h00;      memory[30729] <=  8'h00;      memory[30730] <=  8'h00;      memory[30731] <=  8'h00;      memory[30732] <=  8'h00;      memory[30733] <=  8'h00;      memory[30734] <=  8'h00;      memory[30735] <=  8'h00;      memory[30736] <=  8'h00;      memory[30737] <=  8'h00;      memory[30738] <=  8'h00;      memory[30739] <=  8'h00;      memory[30740] <=  8'h00;      memory[30741] <=  8'h00;      memory[30742] <=  8'h00;      memory[30743] <=  8'h00;      memory[30744] <=  8'h00;      memory[30745] <=  8'h00;      memory[30746] <=  8'h00;      memory[30747] <=  8'h00;      memory[30748] <=  8'h00;      memory[30749] <=  8'h00;      memory[30750] <=  8'h00;      memory[30751] <=  8'h00;      memory[30752] <=  8'h00;      memory[30753] <=  8'h00;      memory[30754] <=  8'h00;      memory[30755] <=  8'h00;      memory[30756] <=  8'h00;      memory[30757] <=  8'h00;      memory[30758] <=  8'h00;      memory[30759] <=  8'h00;      memory[30760] <=  8'h00;      memory[30761] <=  8'h00;      memory[30762] <=  8'h00;      memory[30763] <=  8'h00;      memory[30764] <=  8'h00;      memory[30765] <=  8'h00;      memory[30766] <=  8'h00;      memory[30767] <=  8'h00;      memory[30768] <=  8'h00;      memory[30769] <=  8'h00;      memory[30770] <=  8'h00;      memory[30771] <=  8'h00;      memory[30772] <=  8'h00;      memory[30773] <=  8'h00;      memory[30774] <=  8'h00;      memory[30775] <=  8'h00;      memory[30776] <=  8'h00;      memory[30777] <=  8'h00;      memory[30778] <=  8'h00;      memory[30779] <=  8'h00;      memory[30780] <=  8'h00;      memory[30781] <=  8'h00;      memory[30782] <=  8'h00;      memory[30783] <=  8'h00;      memory[30784] <=  8'h00;      memory[30785] <=  8'h00;      memory[30786] <=  8'h00;      memory[30787] <=  8'h00;      memory[30788] <=  8'h00;      memory[30789] <=  8'h00;      memory[30790] <=  8'h00;      memory[30791] <=  8'h00;      memory[30792] <=  8'h00;      memory[30793] <=  8'h00;      memory[30794] <=  8'h00;      memory[30795] <=  8'h00;      memory[30796] <=  8'h00;      memory[30797] <=  8'h00;      memory[30798] <=  8'h00;      memory[30799] <=  8'h00;      memory[30800] <=  8'h00;      memory[30801] <=  8'h00;      memory[30802] <=  8'h00;      memory[30803] <=  8'h00;      memory[30804] <=  8'h00;      memory[30805] <=  8'h00;      memory[30806] <=  8'h00;      memory[30807] <=  8'h00;      memory[30808] <=  8'h00;      memory[30809] <=  8'h00;      memory[30810] <=  8'h00;      memory[30811] <=  8'h00;      memory[30812] <=  8'h00;      memory[30813] <=  8'h00;      memory[30814] <=  8'h00;      memory[30815] <=  8'h00;      memory[30816] <=  8'h00;      memory[30817] <=  8'h00;      memory[30818] <=  8'h00;      memory[30819] <=  8'h00;      memory[30820] <=  8'h00;      memory[30821] <=  8'h00;      memory[30822] <=  8'h00;      memory[30823] <=  8'h00;      memory[30824] <=  8'h00;      memory[30825] <=  8'h00;      memory[30826] <=  8'h00;      memory[30827] <=  8'h00;      memory[30828] <=  8'h00;      memory[30829] <=  8'h00;      memory[30830] <=  8'h00;      memory[30831] <=  8'h00;      memory[30832] <=  8'h00;      memory[30833] <=  8'h00;      memory[30834] <=  8'h00;      memory[30835] <=  8'h00;      memory[30836] <=  8'h00;      memory[30837] <=  8'h00;      memory[30838] <=  8'h00;      memory[30839] <=  8'h00;      memory[30840] <=  8'h00;      memory[30841] <=  8'h00;      memory[30842] <=  8'h00;      memory[30843] <=  8'h00;      memory[30844] <=  8'h00;      memory[30845] <=  8'h00;      memory[30846] <=  8'h00;      memory[30847] <=  8'h00;      memory[30848] <=  8'h00;      memory[30849] <=  8'h00;      memory[30850] <=  8'h00;      memory[30851] <=  8'h00;      memory[30852] <=  8'h00;      memory[30853] <=  8'h00;      memory[30854] <=  8'h00;      memory[30855] <=  8'h00;      memory[30856] <=  8'h00;      memory[30857] <=  8'h00;      memory[30858] <=  8'h00;      memory[30859] <=  8'h00;      memory[30860] <=  8'h00;      memory[30861] <=  8'h00;      memory[30862] <=  8'h00;      memory[30863] <=  8'h00;      memory[30864] <=  8'h00;      memory[30865] <=  8'h00;      memory[30866] <=  8'h00;      memory[30867] <=  8'h00;      memory[30868] <=  8'h00;      memory[30869] <=  8'h00;      memory[30870] <=  8'h00;      memory[30871] <=  8'h00;      memory[30872] <=  8'h00;      memory[30873] <=  8'h00;      memory[30874] <=  8'h00;      memory[30875] <=  8'h00;      memory[30876] <=  8'h00;      memory[30877] <=  8'h00;      memory[30878] <=  8'h00;      memory[30879] <=  8'h00;      memory[30880] <=  8'h00;      memory[30881] <=  8'h00;      memory[30882] <=  8'h00;      memory[30883] <=  8'h00;      memory[30884] <=  8'h00;      memory[30885] <=  8'h00;      memory[30886] <=  8'h00;      memory[30887] <=  8'h00;      memory[30888] <=  8'h00;      memory[30889] <=  8'h00;      memory[30890] <=  8'h00;      memory[30891] <=  8'h00;      memory[30892] <=  8'h00;      memory[30893] <=  8'h00;      memory[30894] <=  8'h00;      memory[30895] <=  8'h00;      memory[30896] <=  8'h00;      memory[30897] <=  8'h00;      memory[30898] <=  8'h00;      memory[30899] <=  8'h00;      memory[30900] <=  8'h00;      memory[30901] <=  8'h00;      memory[30902] <=  8'h00;      memory[30903] <=  8'h00;      memory[30904] <=  8'h00;      memory[30905] <=  8'h00;      memory[30906] <=  8'h00;      memory[30907] <=  8'h00;      memory[30908] <=  8'h00;      memory[30909] <=  8'h00;      memory[30910] <=  8'h00;      memory[30911] <=  8'h00;      memory[30912] <=  8'h00;      memory[30913] <=  8'h00;      memory[30914] <=  8'h00;      memory[30915] <=  8'h00;      memory[30916] <=  8'h00;      memory[30917] <=  8'h00;      memory[30918] <=  8'h00;      memory[30919] <=  8'h00;      memory[30920] <=  8'h00;      memory[30921] <=  8'h00;      memory[30922] <=  8'h00;      memory[30923] <=  8'h00;      memory[30924] <=  8'h00;      memory[30925] <=  8'h00;      memory[30926] <=  8'h00;      memory[30927] <=  8'h00;      memory[30928] <=  8'h00;      memory[30929] <=  8'h00;      memory[30930] <=  8'h00;      memory[30931] <=  8'h00;      memory[30932] <=  8'h00;      memory[30933] <=  8'h00;      memory[30934] <=  8'h00;      memory[30935] <=  8'h00;      memory[30936] <=  8'h00;      memory[30937] <=  8'h00;      memory[30938] <=  8'h00;      memory[30939] <=  8'h00;      memory[30940] <=  8'h00;      memory[30941] <=  8'h00;      memory[30942] <=  8'h00;      memory[30943] <=  8'h00;      memory[30944] <=  8'h00;      memory[30945] <=  8'h00;      memory[30946] <=  8'h00;      memory[30947] <=  8'h00;      memory[30948] <=  8'h00;      memory[30949] <=  8'h00;      memory[30950] <=  8'h00;      memory[30951] <=  8'h00;      memory[30952] <=  8'h00;      memory[30953] <=  8'h00;      memory[30954] <=  8'h00;      memory[30955] <=  8'h00;      memory[30956] <=  8'h00;      memory[30957] <=  8'h00;      memory[30958] <=  8'h00;      memory[30959] <=  8'h00;      memory[30960] <=  8'h00;      memory[30961] <=  8'h00;      memory[30962] <=  8'h00;      memory[30963] <=  8'h00;      memory[30964] <=  8'h00;      memory[30965] <=  8'h00;      memory[30966] <=  8'h00;      memory[30967] <=  8'h00;      memory[30968] <=  8'h00;      memory[30969] <=  8'h00;      memory[30970] <=  8'h00;      memory[30971] <=  8'h00;      memory[30972] <=  8'h00;      memory[30973] <=  8'h00;      memory[30974] <=  8'h00;      memory[30975] <=  8'h00;      memory[30976] <=  8'h00;      memory[30977] <=  8'h00;      memory[30978] <=  8'h00;      memory[30979] <=  8'h00;      memory[30980] <=  8'h00;      memory[30981] <=  8'h00;      memory[30982] <=  8'h00;      memory[30983] <=  8'h00;      memory[30984] <=  8'h00;      memory[30985] <=  8'h00;      memory[30986] <=  8'h00;      memory[30987] <=  8'h00;      memory[30988] <=  8'h00;      memory[30989] <=  8'h00;      memory[30990] <=  8'h00;      memory[30991] <=  8'h00;      memory[30992] <=  8'h00;      memory[30993] <=  8'h00;      memory[30994] <=  8'h00;      memory[30995] <=  8'h00;      memory[30996] <=  8'h00;      memory[30997] <=  8'h00;      memory[30998] <=  8'h00;      memory[30999] <=  8'h00;      memory[31000] <=  8'h00;      memory[31001] <=  8'h00;      memory[31002] <=  8'h00;      memory[31003] <=  8'h00;      memory[31004] <=  8'h00;      memory[31005] <=  8'h00;      memory[31006] <=  8'h00;      memory[31007] <=  8'h00;      memory[31008] <=  8'h00;      memory[31009] <=  8'h00;      memory[31010] <=  8'h00;      memory[31011] <=  8'h00;      memory[31012] <=  8'h00;      memory[31013] <=  8'h00;      memory[31014] <=  8'h00;      memory[31015] <=  8'h00;      memory[31016] <=  8'h00;      memory[31017] <=  8'h00;      memory[31018] <=  8'h00;      memory[31019] <=  8'h00;      memory[31020] <=  8'h00;      memory[31021] <=  8'h00;      memory[31022] <=  8'h00;      memory[31023] <=  8'h00;      memory[31024] <=  8'h00;      memory[31025] <=  8'h00;      memory[31026] <=  8'h00;      memory[31027] <=  8'h00;      memory[31028] <=  8'h00;      memory[31029] <=  8'h00;      memory[31030] <=  8'h00;      memory[31031] <=  8'h00;      memory[31032] <=  8'h00;      memory[31033] <=  8'h00;      memory[31034] <=  8'h00;      memory[31035] <=  8'h00;      memory[31036] <=  8'h00;      memory[31037] <=  8'h00;      memory[31038] <=  8'h00;      memory[31039] <=  8'h00;      memory[31040] <=  8'h00;      memory[31041] <=  8'h00;      memory[31042] <=  8'h00;      memory[31043] <=  8'h00;      memory[31044] <=  8'h00;      memory[31045] <=  8'h00;      memory[31046] <=  8'h00;      memory[31047] <=  8'h00;      memory[31048] <=  8'h00;      memory[31049] <=  8'h00;      memory[31050] <=  8'h00;      memory[31051] <=  8'h00;      memory[31052] <=  8'h00;      memory[31053] <=  8'h00;      memory[31054] <=  8'h00;      memory[31055] <=  8'h00;      memory[31056] <=  8'h00;      memory[31057] <=  8'h00;      memory[31058] <=  8'h00;      memory[31059] <=  8'h00;      memory[31060] <=  8'h00;      memory[31061] <=  8'h00;      memory[31062] <=  8'h00;      memory[31063] <=  8'h00;      memory[31064] <=  8'h00;      memory[31065] <=  8'h00;      memory[31066] <=  8'h00;      memory[31067] <=  8'h00;      memory[31068] <=  8'h00;      memory[31069] <=  8'h00;      memory[31070] <=  8'h00;      memory[31071] <=  8'h00;      memory[31072] <=  8'h00;      memory[31073] <=  8'h00;      memory[31074] <=  8'h00;      memory[31075] <=  8'h00;      memory[31076] <=  8'h00;      memory[31077] <=  8'h00;      memory[31078] <=  8'h00;      memory[31079] <=  8'h00;      memory[31080] <=  8'h00;      memory[31081] <=  8'h00;      memory[31082] <=  8'h00;      memory[31083] <=  8'h00;      memory[31084] <=  8'h00;      memory[31085] <=  8'h00;      memory[31086] <=  8'h00;      memory[31087] <=  8'h00;      memory[31088] <=  8'h00;      memory[31089] <=  8'h00;      memory[31090] <=  8'h00;      memory[31091] <=  8'h00;      memory[31092] <=  8'h00;      memory[31093] <=  8'h00;      memory[31094] <=  8'h00;      memory[31095] <=  8'h00;      memory[31096] <=  8'h00;      memory[31097] <=  8'h00;      memory[31098] <=  8'h00;      memory[31099] <=  8'h00;      memory[31100] <=  8'h00;      memory[31101] <=  8'h00;      memory[31102] <=  8'h00;      memory[31103] <=  8'h00;      memory[31104] <=  8'h00;      memory[31105] <=  8'h00;      memory[31106] <=  8'h00;      memory[31107] <=  8'h00;      memory[31108] <=  8'h00;      memory[31109] <=  8'h00;      memory[31110] <=  8'h00;      memory[31111] <=  8'h00;      memory[31112] <=  8'h00;      memory[31113] <=  8'h00;      memory[31114] <=  8'h00;      memory[31115] <=  8'h00;      memory[31116] <=  8'h00;      memory[31117] <=  8'h00;      memory[31118] <=  8'h00;      memory[31119] <=  8'h00;      memory[31120] <=  8'h00;      memory[31121] <=  8'h00;      memory[31122] <=  8'h00;      memory[31123] <=  8'h00;      memory[31124] <=  8'h00;      memory[31125] <=  8'h00;      memory[31126] <=  8'h00;      memory[31127] <=  8'h00;      memory[31128] <=  8'h00;      memory[31129] <=  8'h00;      memory[31130] <=  8'h00;      memory[31131] <=  8'h00;      memory[31132] <=  8'h00;      memory[31133] <=  8'h00;      memory[31134] <=  8'h00;      memory[31135] <=  8'h00;      memory[31136] <=  8'h00;      memory[31137] <=  8'h00;      memory[31138] <=  8'h00;      memory[31139] <=  8'h00;      memory[31140] <=  8'h00;      memory[31141] <=  8'h00;      memory[31142] <=  8'h00;      memory[31143] <=  8'h00;      memory[31144] <=  8'h00;      memory[31145] <=  8'h00;      memory[31146] <=  8'h00;      memory[31147] <=  8'h00;      memory[31148] <=  8'h00;      memory[31149] <=  8'h00;      memory[31150] <=  8'h00;      memory[31151] <=  8'h00;      memory[31152] <=  8'h00;      memory[31153] <=  8'h00;      memory[31154] <=  8'h00;      memory[31155] <=  8'h00;      memory[31156] <=  8'h00;      memory[31157] <=  8'h00;      memory[31158] <=  8'h00;      memory[31159] <=  8'h00;      memory[31160] <=  8'h00;      memory[31161] <=  8'h00;      memory[31162] <=  8'h00;      memory[31163] <=  8'h00;      memory[31164] <=  8'h00;      memory[31165] <=  8'h00;      memory[31166] <=  8'h00;      memory[31167] <=  8'h00;      memory[31168] <=  8'h00;      memory[31169] <=  8'h00;      memory[31170] <=  8'h00;      memory[31171] <=  8'h00;      memory[31172] <=  8'h00;      memory[31173] <=  8'h00;      memory[31174] <=  8'h00;      memory[31175] <=  8'h00;      memory[31176] <=  8'h00;      memory[31177] <=  8'h00;      memory[31178] <=  8'h00;      memory[31179] <=  8'h00;      memory[31180] <=  8'h00;      memory[31181] <=  8'h00;      memory[31182] <=  8'h00;      memory[31183] <=  8'h00;      memory[31184] <=  8'h00;      memory[31185] <=  8'h00;      memory[31186] <=  8'h00;      memory[31187] <=  8'h00;      memory[31188] <=  8'h00;      memory[31189] <=  8'h00;      memory[31190] <=  8'h00;      memory[31191] <=  8'h00;      memory[31192] <=  8'h00;      memory[31193] <=  8'h00;      memory[31194] <=  8'h00;      memory[31195] <=  8'h00;      memory[31196] <=  8'h00;      memory[31197] <=  8'h00;      memory[31198] <=  8'h00;      memory[31199] <=  8'h00;      memory[31200] <=  8'h00;      memory[31201] <=  8'h00;      memory[31202] <=  8'h00;      memory[31203] <=  8'h00;      memory[31204] <=  8'h00;      memory[31205] <=  8'h00;      memory[31206] <=  8'h00;      memory[31207] <=  8'h00;      memory[31208] <=  8'h00;      memory[31209] <=  8'h00;      memory[31210] <=  8'h00;      memory[31211] <=  8'h00;      memory[31212] <=  8'h00;      memory[31213] <=  8'h00;      memory[31214] <=  8'h00;      memory[31215] <=  8'h00;      memory[31216] <=  8'h00;      memory[31217] <=  8'h00;      memory[31218] <=  8'h00;      memory[31219] <=  8'h00;      memory[31220] <=  8'h00;      memory[31221] <=  8'h00;      memory[31222] <=  8'h00;      memory[31223] <=  8'h00;      memory[31224] <=  8'h00;      memory[31225] <=  8'h00;      memory[31226] <=  8'h00;      memory[31227] <=  8'h00;      memory[31228] <=  8'h00;      memory[31229] <=  8'h00;      memory[31230] <=  8'h00;      memory[31231] <=  8'h00;      memory[31232] <=  8'h00;      memory[31233] <=  8'h00;      memory[31234] <=  8'h00;      memory[31235] <=  8'h00;      memory[31236] <=  8'h00;      memory[31237] <=  8'h00;      memory[31238] <=  8'h00;      memory[31239] <=  8'h00;      memory[31240] <=  8'h00;      memory[31241] <=  8'h00;      memory[31242] <=  8'h00;      memory[31243] <=  8'h00;      memory[31244] <=  8'h00;      memory[31245] <=  8'h00;      memory[31246] <=  8'h00;      memory[31247] <=  8'h00;      memory[31248] <=  8'h00;      memory[31249] <=  8'h00;      memory[31250] <=  8'h00;      memory[31251] <=  8'h00;      memory[31252] <=  8'h00;      memory[31253] <=  8'h00;      memory[31254] <=  8'h00;      memory[31255] <=  8'h00;      memory[31256] <=  8'h00;      memory[31257] <=  8'h00;      memory[31258] <=  8'h00;      memory[31259] <=  8'h00;      memory[31260] <=  8'h00;      memory[31261] <=  8'h00;      memory[31262] <=  8'h00;      memory[31263] <=  8'h00;      memory[31264] <=  8'h00;      memory[31265] <=  8'h00;      memory[31266] <=  8'h00;      memory[31267] <=  8'h00;      memory[31268] <=  8'h00;      memory[31269] <=  8'h00;      memory[31270] <=  8'h00;      memory[31271] <=  8'h00;      memory[31272] <=  8'h00;      memory[31273] <=  8'h00;      memory[31274] <=  8'h00;      memory[31275] <=  8'h00;      memory[31276] <=  8'h00;      memory[31277] <=  8'h00;      memory[31278] <=  8'h00;      memory[31279] <=  8'h00;      memory[31280] <=  8'h00;      memory[31281] <=  8'h00;      memory[31282] <=  8'h00;      memory[31283] <=  8'h00;      memory[31284] <=  8'h00;      memory[31285] <=  8'h00;      memory[31286] <=  8'h00;      memory[31287] <=  8'h00;      memory[31288] <=  8'h00;      memory[31289] <=  8'h00;      memory[31290] <=  8'h00;      memory[31291] <=  8'h00;      memory[31292] <=  8'h00;      memory[31293] <=  8'h00;      memory[31294] <=  8'h00;      memory[31295] <=  8'h00;      memory[31296] <=  8'h00;      memory[31297] <=  8'h00;      memory[31298] <=  8'h00;      memory[31299] <=  8'h00;      memory[31300] <=  8'h00;      memory[31301] <=  8'h00;      memory[31302] <=  8'h00;      memory[31303] <=  8'h00;      memory[31304] <=  8'h00;      memory[31305] <=  8'h00;      memory[31306] <=  8'h00;      memory[31307] <=  8'h00;      memory[31308] <=  8'h00;      memory[31309] <=  8'h00;      memory[31310] <=  8'h00;      memory[31311] <=  8'h00;      memory[31312] <=  8'h00;      memory[31313] <=  8'h00;      memory[31314] <=  8'h00;      memory[31315] <=  8'h00;      memory[31316] <=  8'h00;      memory[31317] <=  8'h00;      memory[31318] <=  8'h00;      memory[31319] <=  8'h00;      memory[31320] <=  8'h00;      memory[31321] <=  8'h00;      memory[31322] <=  8'h00;      memory[31323] <=  8'h00;      memory[31324] <=  8'h00;      memory[31325] <=  8'h00;      memory[31326] <=  8'h00;      memory[31327] <=  8'h00;      memory[31328] <=  8'h00;      memory[31329] <=  8'h00;      memory[31330] <=  8'h00;      memory[31331] <=  8'h00;      memory[31332] <=  8'h00;      memory[31333] <=  8'h00;      memory[31334] <=  8'h00;      memory[31335] <=  8'h00;      memory[31336] <=  8'h00;      memory[31337] <=  8'h00;      memory[31338] <=  8'h00;      memory[31339] <=  8'h00;      memory[31340] <=  8'h00;      memory[31341] <=  8'h00;      memory[31342] <=  8'h00;      memory[31343] <=  8'h00;      memory[31344] <=  8'h00;      memory[31345] <=  8'h00;      memory[31346] <=  8'h00;      memory[31347] <=  8'h00;      memory[31348] <=  8'h00;      memory[31349] <=  8'h00;      memory[31350] <=  8'h00;      memory[31351] <=  8'h00;      memory[31352] <=  8'h00;      memory[31353] <=  8'h00;      memory[31354] <=  8'h00;      memory[31355] <=  8'h00;      memory[31356] <=  8'h00;      memory[31357] <=  8'h00;      memory[31358] <=  8'h00;      memory[31359] <=  8'h00;      memory[31360] <=  8'h00;      memory[31361] <=  8'h00;      memory[31362] <=  8'h00;      memory[31363] <=  8'h00;      memory[31364] <=  8'h00;      memory[31365] <=  8'h00;      memory[31366] <=  8'h00;      memory[31367] <=  8'h00;      memory[31368] <=  8'h00;      memory[31369] <=  8'h00;      memory[31370] <=  8'h00;      memory[31371] <=  8'h00;      memory[31372] <=  8'h00;      memory[31373] <=  8'h00;      memory[31374] <=  8'h00;      memory[31375] <=  8'h00;      memory[31376] <=  8'h00;      memory[31377] <=  8'h00;      memory[31378] <=  8'h00;      memory[31379] <=  8'h00;      memory[31380] <=  8'h00;      memory[31381] <=  8'h00;      memory[31382] <=  8'h00;      memory[31383] <=  8'h00;      memory[31384] <=  8'h00;      memory[31385] <=  8'h00;      memory[31386] <=  8'h00;      memory[31387] <=  8'h00;      memory[31388] <=  8'h00;      memory[31389] <=  8'h00;      memory[31390] <=  8'h00;      memory[31391] <=  8'h00;      memory[31392] <=  8'h00;      memory[31393] <=  8'h00;      memory[31394] <=  8'h00;      memory[31395] <=  8'h00;      memory[31396] <=  8'h00;      memory[31397] <=  8'h00;      memory[31398] <=  8'h00;      memory[31399] <=  8'h00;      memory[31400] <=  8'h00;      memory[31401] <=  8'h00;      memory[31402] <=  8'h00;      memory[31403] <=  8'h00;      memory[31404] <=  8'h00;      memory[31405] <=  8'h00;      memory[31406] <=  8'h00;      memory[31407] <=  8'h00;      memory[31408] <=  8'h00;      memory[31409] <=  8'h00;      memory[31410] <=  8'h00;      memory[31411] <=  8'h00;      memory[31412] <=  8'h00;      memory[31413] <=  8'h00;      memory[31414] <=  8'h00;      memory[31415] <=  8'h00;      memory[31416] <=  8'h00;      memory[31417] <=  8'h00;      memory[31418] <=  8'h00;      memory[31419] <=  8'h00;      memory[31420] <=  8'h00;      memory[31421] <=  8'h00;      memory[31422] <=  8'h00;      memory[31423] <=  8'h00;      memory[31424] <=  8'h00;      memory[31425] <=  8'h00;      memory[31426] <=  8'h00;      memory[31427] <=  8'h00;      memory[31428] <=  8'h00;      memory[31429] <=  8'h00;      memory[31430] <=  8'h00;      memory[31431] <=  8'h00;      memory[31432] <=  8'h00;      memory[31433] <=  8'h00;      memory[31434] <=  8'h00;      memory[31435] <=  8'h00;      memory[31436] <=  8'h00;      memory[31437] <=  8'h00;      memory[31438] <=  8'h00;      memory[31439] <=  8'h00;      memory[31440] <=  8'h00;      memory[31441] <=  8'h00;      memory[31442] <=  8'h00;      memory[31443] <=  8'h00;      memory[31444] <=  8'h00;      memory[31445] <=  8'h00;      memory[31446] <=  8'h00;      memory[31447] <=  8'h00;      memory[31448] <=  8'h00;      memory[31449] <=  8'h00;      memory[31450] <=  8'h00;      memory[31451] <=  8'h00;      memory[31452] <=  8'h00;      memory[31453] <=  8'h00;      memory[31454] <=  8'h00;      memory[31455] <=  8'h00;      memory[31456] <=  8'h00;      memory[31457] <=  8'h00;      memory[31458] <=  8'h00;      memory[31459] <=  8'h00;      memory[31460] <=  8'h00;      memory[31461] <=  8'h00;      memory[31462] <=  8'h00;      memory[31463] <=  8'h00;      memory[31464] <=  8'h00;      memory[31465] <=  8'h00;      memory[31466] <=  8'h00;      memory[31467] <=  8'h00;      memory[31468] <=  8'h00;      memory[31469] <=  8'h00;      memory[31470] <=  8'h00;      memory[31471] <=  8'h00;      memory[31472] <=  8'h00;      memory[31473] <=  8'h00;      memory[31474] <=  8'h00;      memory[31475] <=  8'h00;      memory[31476] <=  8'h00;      memory[31477] <=  8'h00;      memory[31478] <=  8'h00;      memory[31479] <=  8'h00;      memory[31480] <=  8'h00;      memory[31481] <=  8'h00;      memory[31482] <=  8'h00;      memory[31483] <=  8'h00;      memory[31484] <=  8'h00;      memory[31485] <=  8'h00;      memory[31486] <=  8'h00;      memory[31487] <=  8'h00;      memory[31488] <=  8'h00;      memory[31489] <=  8'h00;      memory[31490] <=  8'h00;      memory[31491] <=  8'h00;      memory[31492] <=  8'h00;      memory[31493] <=  8'h00;      memory[31494] <=  8'h00;      memory[31495] <=  8'h00;      memory[31496] <=  8'h00;      memory[31497] <=  8'h00;      memory[31498] <=  8'h00;      memory[31499] <=  8'h00;      memory[31500] <=  8'h00;      memory[31501] <=  8'h00;      memory[31502] <=  8'h00;      memory[31503] <=  8'h00;      memory[31504] <=  8'h00;      memory[31505] <=  8'h00;      memory[31506] <=  8'h00;      memory[31507] <=  8'h00;      memory[31508] <=  8'h00;      memory[31509] <=  8'h00;      memory[31510] <=  8'h00;      memory[31511] <=  8'h00;      memory[31512] <=  8'h00;      memory[31513] <=  8'h00;      memory[31514] <=  8'h00;      memory[31515] <=  8'h00;      memory[31516] <=  8'h00;      memory[31517] <=  8'h00;      memory[31518] <=  8'h00;      memory[31519] <=  8'h00;      memory[31520] <=  8'h00;      memory[31521] <=  8'h00;      memory[31522] <=  8'h00;      memory[31523] <=  8'h00;      memory[31524] <=  8'h00;      memory[31525] <=  8'h00;      memory[31526] <=  8'h00;      memory[31527] <=  8'h00;      memory[31528] <=  8'h00;      memory[31529] <=  8'h00;      memory[31530] <=  8'h00;      memory[31531] <=  8'h00;      memory[31532] <=  8'h00;      memory[31533] <=  8'h00;      memory[31534] <=  8'h00;      memory[31535] <=  8'h00;      memory[31536] <=  8'h00;      memory[31537] <=  8'h00;      memory[31538] <=  8'h00;      memory[31539] <=  8'h00;      memory[31540] <=  8'h00;      memory[31541] <=  8'h00;      memory[31542] <=  8'h00;      memory[31543] <=  8'h00;      memory[31544] <=  8'h00;      memory[31545] <=  8'h00;      memory[31546] <=  8'h00;      memory[31547] <=  8'h00;      memory[31548] <=  8'h00;      memory[31549] <=  8'h00;      memory[31550] <=  8'h00;      memory[31551] <=  8'h00;      memory[31552] <=  8'h00;      memory[31553] <=  8'h00;      memory[31554] <=  8'h00;      memory[31555] <=  8'h00;      memory[31556] <=  8'h00;      memory[31557] <=  8'h00;      memory[31558] <=  8'h00;      memory[31559] <=  8'h00;      memory[31560] <=  8'h00;      memory[31561] <=  8'h00;      memory[31562] <=  8'h00;      memory[31563] <=  8'h00;      memory[31564] <=  8'h00;      memory[31565] <=  8'h00;      memory[31566] <=  8'h00;      memory[31567] <=  8'h00;      memory[31568] <=  8'h00;      memory[31569] <=  8'h00;      memory[31570] <=  8'h00;      memory[31571] <=  8'h00;      memory[31572] <=  8'h00;      memory[31573] <=  8'h00;      memory[31574] <=  8'h00;      memory[31575] <=  8'h00;      memory[31576] <=  8'h00;      memory[31577] <=  8'h00;      memory[31578] <=  8'h00;      memory[31579] <=  8'h00;      memory[31580] <=  8'h00;      memory[31581] <=  8'h00;      memory[31582] <=  8'h00;      memory[31583] <=  8'h00;      memory[31584] <=  8'h00;      memory[31585] <=  8'h00;      memory[31586] <=  8'h00;      memory[31587] <=  8'h00;      memory[31588] <=  8'h00;      memory[31589] <=  8'h00;      memory[31590] <=  8'h00;      memory[31591] <=  8'h00;      memory[31592] <=  8'h00;      memory[31593] <=  8'h00;      memory[31594] <=  8'h00;      memory[31595] <=  8'h00;      memory[31596] <=  8'h00;      memory[31597] <=  8'h00;      memory[31598] <=  8'h00;      memory[31599] <=  8'h00;      memory[31600] <=  8'h00;      memory[31601] <=  8'h00;      memory[31602] <=  8'h00;      memory[31603] <=  8'h00;      memory[31604] <=  8'h00;      memory[31605] <=  8'h00;      memory[31606] <=  8'h00;      memory[31607] <=  8'h00;      memory[31608] <=  8'h00;      memory[31609] <=  8'h00;      memory[31610] <=  8'h00;      memory[31611] <=  8'h00;      memory[31612] <=  8'h00;      memory[31613] <=  8'h00;      memory[31614] <=  8'h00;      memory[31615] <=  8'h00;      memory[31616] <=  8'h00;      memory[31617] <=  8'h00;      memory[31618] <=  8'h00;      memory[31619] <=  8'h00;      memory[31620] <=  8'h00;      memory[31621] <=  8'h00;      memory[31622] <=  8'h00;      memory[31623] <=  8'h00;      memory[31624] <=  8'h00;      memory[31625] <=  8'h00;      memory[31626] <=  8'h00;      memory[31627] <=  8'h00;      memory[31628] <=  8'h00;      memory[31629] <=  8'h00;      memory[31630] <=  8'h00;      memory[31631] <=  8'h00;      memory[31632] <=  8'h00;      memory[31633] <=  8'h00;      memory[31634] <=  8'h00;      memory[31635] <=  8'h00;      memory[31636] <=  8'h00;      memory[31637] <=  8'h00;      memory[31638] <=  8'h00;      memory[31639] <=  8'h00;      memory[31640] <=  8'h00;      memory[31641] <=  8'h00;      memory[31642] <=  8'h00;      memory[31643] <=  8'h00;      memory[31644] <=  8'h00;      memory[31645] <=  8'h00;      memory[31646] <=  8'h00;      memory[31647] <=  8'h00;      memory[31648] <=  8'h00;      memory[31649] <=  8'h00;      memory[31650] <=  8'h00;      memory[31651] <=  8'h00;      memory[31652] <=  8'h00;      memory[31653] <=  8'h00;      memory[31654] <=  8'h00;      memory[31655] <=  8'h00;      memory[31656] <=  8'h00;      memory[31657] <=  8'h00;      memory[31658] <=  8'h00;      memory[31659] <=  8'h00;      memory[31660] <=  8'h00;      memory[31661] <=  8'h00;      memory[31662] <=  8'h00;      memory[31663] <=  8'h00;      memory[31664] <=  8'h00;      memory[31665] <=  8'h00;      memory[31666] <=  8'h00;      memory[31667] <=  8'h00;      memory[31668] <=  8'h00;      memory[31669] <=  8'h00;      memory[31670] <=  8'h00;      memory[31671] <=  8'h00;      memory[31672] <=  8'h00;      memory[31673] <=  8'h00;      memory[31674] <=  8'h00;      memory[31675] <=  8'h00;      memory[31676] <=  8'h00;      memory[31677] <=  8'h00;      memory[31678] <=  8'h00;      memory[31679] <=  8'h00;      memory[31680] <=  8'h00;      memory[31681] <=  8'h00;      memory[31682] <=  8'h00;      memory[31683] <=  8'h00;      memory[31684] <=  8'h00;      memory[31685] <=  8'h00;      memory[31686] <=  8'h00;      memory[31687] <=  8'h00;      memory[31688] <=  8'h00;      memory[31689] <=  8'h00;      memory[31690] <=  8'h00;      memory[31691] <=  8'h00;      memory[31692] <=  8'h00;      memory[31693] <=  8'h00;      memory[31694] <=  8'h00;      memory[31695] <=  8'h00;      memory[31696] <=  8'h00;      memory[31697] <=  8'h00;      memory[31698] <=  8'h00;      memory[31699] <=  8'h00;      memory[31700] <=  8'h00;      memory[31701] <=  8'h00;      memory[31702] <=  8'h00;      memory[31703] <=  8'h00;      memory[31704] <=  8'h00;      memory[31705] <=  8'h00;      memory[31706] <=  8'h00;      memory[31707] <=  8'h00;      memory[31708] <=  8'h00;      memory[31709] <=  8'h00;      memory[31710] <=  8'h00;      memory[31711] <=  8'h00;      memory[31712] <=  8'h00;      memory[31713] <=  8'h00;      memory[31714] <=  8'h00;      memory[31715] <=  8'h00;      memory[31716] <=  8'h00;      memory[31717] <=  8'h00;      memory[31718] <=  8'h00;      memory[31719] <=  8'h00;      memory[31720] <=  8'h00;      memory[31721] <=  8'h00;      memory[31722] <=  8'h00;      memory[31723] <=  8'h00;      memory[31724] <=  8'h00;      memory[31725] <=  8'h00;      memory[31726] <=  8'h00;      memory[31727] <=  8'h00;      memory[31728] <=  8'h00;      memory[31729] <=  8'h00;      memory[31730] <=  8'h00;      memory[31731] <=  8'h00;      memory[31732] <=  8'h00;      memory[31733] <=  8'h00;      memory[31734] <=  8'h00;      memory[31735] <=  8'h00;      memory[31736] <=  8'h00;      memory[31737] <=  8'h00;      memory[31738] <=  8'h00;      memory[31739] <=  8'h00;      memory[31740] <=  8'h00;      memory[31741] <=  8'h00;      memory[31742] <=  8'h00;      memory[31743] <=  8'h00;      memory[31744] <=  8'h00;      memory[31745] <=  8'h00;      memory[31746] <=  8'h00;      memory[31747] <=  8'h00;      memory[31748] <=  8'h00;      memory[31749] <=  8'h00;      memory[31750] <=  8'h00;      memory[31751] <=  8'h00;      memory[31752] <=  8'h00;      memory[31753] <=  8'h00;      memory[31754] <=  8'h00;      memory[31755] <=  8'h00;      memory[31756] <=  8'h00;      memory[31757] <=  8'h00;      memory[31758] <=  8'h00;      memory[31759] <=  8'h00;      memory[31760] <=  8'h00;      memory[31761] <=  8'h00;      memory[31762] <=  8'h00;      memory[31763] <=  8'h00;      memory[31764] <=  8'h00;      memory[31765] <=  8'h00;      memory[31766] <=  8'h00;      memory[31767] <=  8'h00;      memory[31768] <=  8'h00;      memory[31769] <=  8'h00;      memory[31770] <=  8'h00;      memory[31771] <=  8'h00;      memory[31772] <=  8'h00;      memory[31773] <=  8'h00;      memory[31774] <=  8'h00;      memory[31775] <=  8'h00;      memory[31776] <=  8'h00;      memory[31777] <=  8'h00;      memory[31778] <=  8'h00;      memory[31779] <=  8'h00;      memory[31780] <=  8'h00;      memory[31781] <=  8'h00;      memory[31782] <=  8'h00;      memory[31783] <=  8'h00;      memory[31784] <=  8'h00;      memory[31785] <=  8'h00;      memory[31786] <=  8'h00;      memory[31787] <=  8'h00;      memory[31788] <=  8'h00;      memory[31789] <=  8'h00;      memory[31790] <=  8'h00;      memory[31791] <=  8'h00;      memory[31792] <=  8'h00;      memory[31793] <=  8'h00;      memory[31794] <=  8'h00;      memory[31795] <=  8'h00;      memory[31796] <=  8'h00;      memory[31797] <=  8'h00;      memory[31798] <=  8'h00;      memory[31799] <=  8'h00;      memory[31800] <=  8'h00;      memory[31801] <=  8'h00;      memory[31802] <=  8'h00;      memory[31803] <=  8'h00;      memory[31804] <=  8'h00;      memory[31805] <=  8'h00;      memory[31806] <=  8'h00;      memory[31807] <=  8'h00;      memory[31808] <=  8'h00;      memory[31809] <=  8'h00;      memory[31810] <=  8'h00;      memory[31811] <=  8'h00;      memory[31812] <=  8'h00;      memory[31813] <=  8'h00;      memory[31814] <=  8'h00;      memory[31815] <=  8'h00;      memory[31816] <=  8'h00;      memory[31817] <=  8'h00;      memory[31818] <=  8'h00;      memory[31819] <=  8'h00;      memory[31820] <=  8'h00;      memory[31821] <=  8'h00;      memory[31822] <=  8'h00;      memory[31823] <=  8'h00;      memory[31824] <=  8'h00;      memory[31825] <=  8'h00;      memory[31826] <=  8'h00;      memory[31827] <=  8'h00;      memory[31828] <=  8'h00;      memory[31829] <=  8'h00;      memory[31830] <=  8'h00;      memory[31831] <=  8'h00;      memory[31832] <=  8'h00;      memory[31833] <=  8'h00;      memory[31834] <=  8'h00;      memory[31835] <=  8'h00;      memory[31836] <=  8'h00;      memory[31837] <=  8'h00;      memory[31838] <=  8'h00;      memory[31839] <=  8'h00;      memory[31840] <=  8'h00;      memory[31841] <=  8'h00;      memory[31842] <=  8'h00;      memory[31843] <=  8'h00;      memory[31844] <=  8'h00;      memory[31845] <=  8'h00;      memory[31846] <=  8'h00;      memory[31847] <=  8'h00;      memory[31848] <=  8'h00;      memory[31849] <=  8'h00;      memory[31850] <=  8'h00;      memory[31851] <=  8'h00;      memory[31852] <=  8'h00;      memory[31853] <=  8'h00;      memory[31854] <=  8'h00;      memory[31855] <=  8'h00;      memory[31856] <=  8'h00;      memory[31857] <=  8'h00;      memory[31858] <=  8'h00;      memory[31859] <=  8'h00;      memory[31860] <=  8'h00;      memory[31861] <=  8'h00;      memory[31862] <=  8'h00;      memory[31863] <=  8'h00;      memory[31864] <=  8'h00;      memory[31865] <=  8'h00;      memory[31866] <=  8'h00;      memory[31867] <=  8'h00;      memory[31868] <=  8'h00;      memory[31869] <=  8'h00;      memory[31870] <=  8'h00;      memory[31871] <=  8'h00;      memory[31872] <=  8'h00;      memory[31873] <=  8'h00;      memory[31874] <=  8'h00;      memory[31875] <=  8'h00;      memory[31876] <=  8'h00;      memory[31877] <=  8'h00;      memory[31878] <=  8'h00;      memory[31879] <=  8'h00;      memory[31880] <=  8'h00;      memory[31881] <=  8'h00;      memory[31882] <=  8'h00;      memory[31883] <=  8'h00;      memory[31884] <=  8'h00;      memory[31885] <=  8'h00;      memory[31886] <=  8'h00;      memory[31887] <=  8'h00;      memory[31888] <=  8'h00;      memory[31889] <=  8'h00;      memory[31890] <=  8'h00;      memory[31891] <=  8'h00;      memory[31892] <=  8'h00;      memory[31893] <=  8'h00;      memory[31894] <=  8'h00;      memory[31895] <=  8'h00;      memory[31896] <=  8'h00;      memory[31897] <=  8'h00;      memory[31898] <=  8'h00;      memory[31899] <=  8'h00;      memory[31900] <=  8'h00;      memory[31901] <=  8'h00;      memory[31902] <=  8'h00;      memory[31903] <=  8'h00;      memory[31904] <=  8'h00;      memory[31905] <=  8'h00;      memory[31906] <=  8'h00;      memory[31907] <=  8'h00;      memory[31908] <=  8'h00;      memory[31909] <=  8'h00;      memory[31910] <=  8'h00;      memory[31911] <=  8'h00;      memory[31912] <=  8'h00;      memory[31913] <=  8'h00;      memory[31914] <=  8'h00;      memory[31915] <=  8'h00;      memory[31916] <=  8'h00;      memory[31917] <=  8'h00;      memory[31918] <=  8'h00;      memory[31919] <=  8'h00;      memory[31920] <=  8'h00;      memory[31921] <=  8'h00;      memory[31922] <=  8'h00;      memory[31923] <=  8'h00;      memory[31924] <=  8'h00;      memory[31925] <=  8'h00;      memory[31926] <=  8'h00;      memory[31927] <=  8'h00;      memory[31928] <=  8'h00;      memory[31929] <=  8'h00;      memory[31930] <=  8'h00;      memory[31931] <=  8'h00;      memory[31932] <=  8'h00;      memory[31933] <=  8'h00;      memory[31934] <=  8'h00;      memory[31935] <=  8'h00;      memory[31936] <=  8'h00;      memory[31937] <=  8'h00;      memory[31938] <=  8'h00;      memory[31939] <=  8'h00;      memory[31940] <=  8'h00;      memory[31941] <=  8'h00;      memory[31942] <=  8'h00;      memory[31943] <=  8'h00;      memory[31944] <=  8'h00;      memory[31945] <=  8'h00;      memory[31946] <=  8'h00;      memory[31947] <=  8'h00;      memory[31948] <=  8'h00;      memory[31949] <=  8'h00;      memory[31950] <=  8'h00;      memory[31951] <=  8'h00;      memory[31952] <=  8'h00;      memory[31953] <=  8'h00;      memory[31954] <=  8'h00;      memory[31955] <=  8'h00;      memory[31956] <=  8'h00;      memory[31957] <=  8'h00;      memory[31958] <=  8'h00;      memory[31959] <=  8'h00;      memory[31960] <=  8'h00;      memory[31961] <=  8'h00;      memory[31962] <=  8'h00;      memory[31963] <=  8'h00;      memory[31964] <=  8'h00;      memory[31965] <=  8'h00;      memory[31966] <=  8'h00;      memory[31967] <=  8'h00;      memory[31968] <=  8'h00;      memory[31969] <=  8'h00;      memory[31970] <=  8'h00;      memory[31971] <=  8'h00;      memory[31972] <=  8'h00;      memory[31973] <=  8'h00;      memory[31974] <=  8'h00;      memory[31975] <=  8'h00;      memory[31976] <=  8'h00;      memory[31977] <=  8'h00;      memory[31978] <=  8'h00;      memory[31979] <=  8'h00;      memory[31980] <=  8'h00;      memory[31981] <=  8'h00;      memory[31982] <=  8'h00;      memory[31983] <=  8'h00;      memory[31984] <=  8'h00;      memory[31985] <=  8'h00;      memory[31986] <=  8'h00;      memory[31987] <=  8'h00;      memory[31988] <=  8'h00;      memory[31989] <=  8'h00;      memory[31990] <=  8'h00;      memory[31991] <=  8'h00;      memory[31992] <=  8'h00;      memory[31993] <=  8'h00;      memory[31994] <=  8'h00;      memory[31995] <=  8'h00;      memory[31996] <=  8'h00;      memory[31997] <=  8'h00;      memory[31998] <=  8'h00;      memory[31999] <=  8'h00;      memory[32000] <=  8'h00;      memory[32001] <=  8'h00;      memory[32002] <=  8'h00;      memory[32003] <=  8'h00;      memory[32004] <=  8'h00;      memory[32005] <=  8'h00;      memory[32006] <=  8'h00;      memory[32007] <=  8'h00;      memory[32008] <=  8'h00;      memory[32009] <=  8'h00;      memory[32010] <=  8'h00;      memory[32011] <=  8'h00;      memory[32012] <=  8'h00;      memory[32013] <=  8'h00;      memory[32014] <=  8'h00;      memory[32015] <=  8'h00;      memory[32016] <=  8'h00;      memory[32017] <=  8'h00;      memory[32018] <=  8'h00;      memory[32019] <=  8'h00;      memory[32020] <=  8'h00;      memory[32021] <=  8'h00;      memory[32022] <=  8'h00;      memory[32023] <=  8'h00;      memory[32024] <=  8'h00;      memory[32025] <=  8'h00;      memory[32026] <=  8'h00;      memory[32027] <=  8'h00;      memory[32028] <=  8'h00;      memory[32029] <=  8'h00;      memory[32030] <=  8'h00;      memory[32031] <=  8'h00;      memory[32032] <=  8'h00;      memory[32033] <=  8'h00;      memory[32034] <=  8'h00;      memory[32035] <=  8'h00;      memory[32036] <=  8'h00;      memory[32037] <=  8'h00;      memory[32038] <=  8'h00;      memory[32039] <=  8'h00;      memory[32040] <=  8'h00;      memory[32041] <=  8'h00;      memory[32042] <=  8'h00;      memory[32043] <=  8'h00;      memory[32044] <=  8'h00;      memory[32045] <=  8'h00;      memory[32046] <=  8'h00;      memory[32047] <=  8'h00;      memory[32048] <=  8'h00;      memory[32049] <=  8'h00;      memory[32050] <=  8'h00;      memory[32051] <=  8'h00;      memory[32052] <=  8'h00;      memory[32053] <=  8'h00;      memory[32054] <=  8'h00;      memory[32055] <=  8'h00;      memory[32056] <=  8'h00;      memory[32057] <=  8'h00;      memory[32058] <=  8'h00;      memory[32059] <=  8'h00;      memory[32060] <=  8'h00;      memory[32061] <=  8'h00;      memory[32062] <=  8'h00;      memory[32063] <=  8'h00;      memory[32064] <=  8'h00;      memory[32065] <=  8'h00;      memory[32066] <=  8'h00;      memory[32067] <=  8'h00;      memory[32068] <=  8'h00;      memory[32069] <=  8'h00;      memory[32070] <=  8'h00;      memory[32071] <=  8'h00;      memory[32072] <=  8'h00;      memory[32073] <=  8'h00;      memory[32074] <=  8'h00;      memory[32075] <=  8'h00;      memory[32076] <=  8'h00;      memory[32077] <=  8'h00;      memory[32078] <=  8'h00;      memory[32079] <=  8'h00;      memory[32080] <=  8'h00;      memory[32081] <=  8'h00;      memory[32082] <=  8'h00;      memory[32083] <=  8'h00;      memory[32084] <=  8'h00;      memory[32085] <=  8'h00;      memory[32086] <=  8'h00;      memory[32087] <=  8'h00;      memory[32088] <=  8'h00;      memory[32089] <=  8'h00;      memory[32090] <=  8'h00;      memory[32091] <=  8'h00;      memory[32092] <=  8'h00;      memory[32093] <=  8'h00;      memory[32094] <=  8'h00;      memory[32095] <=  8'h00;      memory[32096] <=  8'h00;      memory[32097] <=  8'h00;      memory[32098] <=  8'h00;      memory[32099] <=  8'h00;      memory[32100] <=  8'h00;      memory[32101] <=  8'h00;      memory[32102] <=  8'h00;      memory[32103] <=  8'h00;      memory[32104] <=  8'h00;      memory[32105] <=  8'h00;      memory[32106] <=  8'h00;      memory[32107] <=  8'h00;      memory[32108] <=  8'h00;      memory[32109] <=  8'h00;      memory[32110] <=  8'h00;      memory[32111] <=  8'h00;      memory[32112] <=  8'h00;      memory[32113] <=  8'h00;      memory[32114] <=  8'h00;      memory[32115] <=  8'h00;      memory[32116] <=  8'h00;      memory[32117] <=  8'h00;      memory[32118] <=  8'h00;      memory[32119] <=  8'h00;      memory[32120] <=  8'h00;      memory[32121] <=  8'h00;      memory[32122] <=  8'h00;      memory[32123] <=  8'h00;      memory[32124] <=  8'h00;      memory[32125] <=  8'h00;      memory[32126] <=  8'h00;      memory[32127] <=  8'h00;      memory[32128] <=  8'h00;      memory[32129] <=  8'h00;      memory[32130] <=  8'h00;      memory[32131] <=  8'h00;      memory[32132] <=  8'h00;      memory[32133] <=  8'h00;      memory[32134] <=  8'h00;      memory[32135] <=  8'h00;      memory[32136] <=  8'h00;      memory[32137] <=  8'h00;      memory[32138] <=  8'h00;      memory[32139] <=  8'h00;      memory[32140] <=  8'h00;      memory[32141] <=  8'h00;      memory[32142] <=  8'h00;      memory[32143] <=  8'h00;      memory[32144] <=  8'h00;      memory[32145] <=  8'h00;      memory[32146] <=  8'h00;      memory[32147] <=  8'h00;      memory[32148] <=  8'h00;      memory[32149] <=  8'h00;      memory[32150] <=  8'h00;      memory[32151] <=  8'h00;      memory[32152] <=  8'h00;      memory[32153] <=  8'h00;      memory[32154] <=  8'h00;      memory[32155] <=  8'h00;      memory[32156] <=  8'h00;      memory[32157] <=  8'h00;      memory[32158] <=  8'h00;      memory[32159] <=  8'h00;      memory[32160] <=  8'h00;      memory[32161] <=  8'h00;      memory[32162] <=  8'h00;      memory[32163] <=  8'h00;      memory[32164] <=  8'h00;      memory[32165] <=  8'h00;      memory[32166] <=  8'h00;      memory[32167] <=  8'h00;      memory[32168] <=  8'h00;      memory[32169] <=  8'h00;      memory[32170] <=  8'h00;      memory[32171] <=  8'h00;      memory[32172] <=  8'h00;      memory[32173] <=  8'h00;      memory[32174] <=  8'h00;      memory[32175] <=  8'h00;      memory[32176] <=  8'h00;      memory[32177] <=  8'h00;      memory[32178] <=  8'h00;      memory[32179] <=  8'h00;      memory[32180] <=  8'h00;      memory[32181] <=  8'h00;      memory[32182] <=  8'h00;      memory[32183] <=  8'h00;      memory[32184] <=  8'h00;      memory[32185] <=  8'h00;      memory[32186] <=  8'h00;      memory[32187] <=  8'h00;      memory[32188] <=  8'h00;      memory[32189] <=  8'h00;      memory[32190] <=  8'h00;      memory[32191] <=  8'h00;      memory[32192] <=  8'h00;      memory[32193] <=  8'h00;      memory[32194] <=  8'h00;      memory[32195] <=  8'h00;      memory[32196] <=  8'h00;      memory[32197] <=  8'h00;      memory[32198] <=  8'h00;      memory[32199] <=  8'h00;      memory[32200] <=  8'h00;      memory[32201] <=  8'h00;      memory[32202] <=  8'h00;      memory[32203] <=  8'h00;      memory[32204] <=  8'h00;      memory[32205] <=  8'h00;      memory[32206] <=  8'h00;      memory[32207] <=  8'h00;      memory[32208] <=  8'h00;      memory[32209] <=  8'h00;      memory[32210] <=  8'h00;      memory[32211] <=  8'h00;      memory[32212] <=  8'h00;      memory[32213] <=  8'h00;      memory[32214] <=  8'h00;      memory[32215] <=  8'h00;      memory[32216] <=  8'h00;      memory[32217] <=  8'h00;      memory[32218] <=  8'h00;      memory[32219] <=  8'h00;      memory[32220] <=  8'h00;      memory[32221] <=  8'h00;      memory[32222] <=  8'h00;      memory[32223] <=  8'h00;      memory[32224] <=  8'h00;      memory[32225] <=  8'h00;      memory[32226] <=  8'h00;      memory[32227] <=  8'h00;      memory[32228] <=  8'h00;      memory[32229] <=  8'h00;      memory[32230] <=  8'h00;      memory[32231] <=  8'h00;      memory[32232] <=  8'h00;      memory[32233] <=  8'h00;      memory[32234] <=  8'h00;      memory[32235] <=  8'h00;      memory[32236] <=  8'h00;      memory[32237] <=  8'h00;      memory[32238] <=  8'h00;      memory[32239] <=  8'h00;      memory[32240] <=  8'h00;      memory[32241] <=  8'h00;      memory[32242] <=  8'h00;      memory[32243] <=  8'h00;      memory[32244] <=  8'h00;      memory[32245] <=  8'h00;      memory[32246] <=  8'h00;      memory[32247] <=  8'h00;      memory[32248] <=  8'h00;      memory[32249] <=  8'h00;      memory[32250] <=  8'h00;      memory[32251] <=  8'h00;      memory[32252] <=  8'h00;      memory[32253] <=  8'h00;      memory[32254] <=  8'h00;      memory[32255] <=  8'h00;      memory[32256] <=  8'h00;      memory[32257] <=  8'h00;      memory[32258] <=  8'h00;      memory[32259] <=  8'h00;      memory[32260] <=  8'h00;      memory[32261] <=  8'h00;      memory[32262] <=  8'h00;      memory[32263] <=  8'h00;      memory[32264] <=  8'h00;      memory[32265] <=  8'h00;      memory[32266] <=  8'h00;      memory[32267] <=  8'h00;      memory[32268] <=  8'h00;      memory[32269] <=  8'h00;      memory[32270] <=  8'h00;      memory[32271] <=  8'h00;      memory[32272] <=  8'h00;      memory[32273] <=  8'h00;      memory[32274] <=  8'h00;      memory[32275] <=  8'h00;      memory[32276] <=  8'h00;      memory[32277] <=  8'h00;      memory[32278] <=  8'h00;      memory[32279] <=  8'h00;      memory[32280] <=  8'h00;      memory[32281] <=  8'h00;      memory[32282] <=  8'h00;      memory[32283] <=  8'h00;      memory[32284] <=  8'h00;      memory[32285] <=  8'h00;      memory[32286] <=  8'h00;      memory[32287] <=  8'h00;      memory[32288] <=  8'h00;      memory[32289] <=  8'h00;      memory[32290] <=  8'h00;      memory[32291] <=  8'h00;      memory[32292] <=  8'h00;      memory[32293] <=  8'h00;      memory[32294] <=  8'h00;      memory[32295] <=  8'h00;      memory[32296] <=  8'h00;      memory[32297] <=  8'h00;      memory[32298] <=  8'h00;      memory[32299] <=  8'h00;      memory[32300] <=  8'h00;      memory[32301] <=  8'h00;      memory[32302] <=  8'h00;      memory[32303] <=  8'h00;      memory[32304] <=  8'h00;      memory[32305] <=  8'h00;      memory[32306] <=  8'h00;      memory[32307] <=  8'h00;      memory[32308] <=  8'h00;      memory[32309] <=  8'h00;      memory[32310] <=  8'h00;      memory[32311] <=  8'h00;      memory[32312] <=  8'h00;      memory[32313] <=  8'h00;      memory[32314] <=  8'h00;      memory[32315] <=  8'h00;      memory[32316] <=  8'h00;      memory[32317] <=  8'h00;      memory[32318] <=  8'h00;      memory[32319] <=  8'h00;      memory[32320] <=  8'h00;      memory[32321] <=  8'h00;      memory[32322] <=  8'h00;      memory[32323] <=  8'h00;      memory[32324] <=  8'h00;      memory[32325] <=  8'h00;      memory[32326] <=  8'h00;      memory[32327] <=  8'h00;      memory[32328] <=  8'h00;      memory[32329] <=  8'h00;      memory[32330] <=  8'h00;      memory[32331] <=  8'h00;      memory[32332] <=  8'h00;      memory[32333] <=  8'h00;      memory[32334] <=  8'h00;      memory[32335] <=  8'h00;      memory[32336] <=  8'h00;      memory[32337] <=  8'h00;      memory[32338] <=  8'h00;      memory[32339] <=  8'h00;      memory[32340] <=  8'h00;      memory[32341] <=  8'h00;      memory[32342] <=  8'h00;      memory[32343] <=  8'h00;      memory[32344] <=  8'h00;      memory[32345] <=  8'h00;      memory[32346] <=  8'h00;      memory[32347] <=  8'h00;      memory[32348] <=  8'h00;      memory[32349] <=  8'h00;      memory[32350] <=  8'h00;      memory[32351] <=  8'h00;      memory[32352] <=  8'h00;      memory[32353] <=  8'h00;      memory[32354] <=  8'h00;      memory[32355] <=  8'h00;      memory[32356] <=  8'h00;      memory[32357] <=  8'h00;      memory[32358] <=  8'h00;      memory[32359] <=  8'h00;      memory[32360] <=  8'h00;      memory[32361] <=  8'h00;      memory[32362] <=  8'h00;      memory[32363] <=  8'h00;      memory[32364] <=  8'h00;      memory[32365] <=  8'h00;      memory[32366] <=  8'h00;      memory[32367] <=  8'h00;      memory[32368] <=  8'h00;      memory[32369] <=  8'h00;      memory[32370] <=  8'h00;      memory[32371] <=  8'h00;      memory[32372] <=  8'h00;      memory[32373] <=  8'h00;      memory[32374] <=  8'h00;      memory[32375] <=  8'h00;      memory[32376] <=  8'h00;      memory[32377] <=  8'h00;      memory[32378] <=  8'h00;      memory[32379] <=  8'h00;      memory[32380] <=  8'h00;      memory[32381] <=  8'h00;      memory[32382] <=  8'h00;      memory[32383] <=  8'h00;      memory[32384] <=  8'h00;      memory[32385] <=  8'h00;      memory[32386] <=  8'h00;      memory[32387] <=  8'h00;      memory[32388] <=  8'h00;      memory[32389] <=  8'h00;      memory[32390] <=  8'h00;      memory[32391] <=  8'h00;      memory[32392] <=  8'h00;      memory[32393] <=  8'h00;      memory[32394] <=  8'h00;      memory[32395] <=  8'h00;      memory[32396] <=  8'h00;      memory[32397] <=  8'h00;      memory[32398] <=  8'h00;      memory[32399] <=  8'h00;      memory[32400] <=  8'h00;      memory[32401] <=  8'h00;      memory[32402] <=  8'h00;      memory[32403] <=  8'h00;      memory[32404] <=  8'h00;      memory[32405] <=  8'h00;      memory[32406] <=  8'h00;      memory[32407] <=  8'h00;      memory[32408] <=  8'h00;      memory[32409] <=  8'h00;      memory[32410] <=  8'h00;      memory[32411] <=  8'h00;      memory[32412] <=  8'h00;      memory[32413] <=  8'h00;      memory[32414] <=  8'h00;      memory[32415] <=  8'h00;      memory[32416] <=  8'h00;      memory[32417] <=  8'h00;      memory[32418] <=  8'h00;      memory[32419] <=  8'h00;      memory[32420] <=  8'h00;      memory[32421] <=  8'h00;      memory[32422] <=  8'h00;      memory[32423] <=  8'h00;      memory[32424] <=  8'h00;      memory[32425] <=  8'h00;      memory[32426] <=  8'h00;      memory[32427] <=  8'h00;      memory[32428] <=  8'h00;      memory[32429] <=  8'h00;      memory[32430] <=  8'h00;      memory[32431] <=  8'h00;      memory[32432] <=  8'h00;      memory[32433] <=  8'h00;      memory[32434] <=  8'h00;      memory[32435] <=  8'h00;      memory[32436] <=  8'h00;      memory[32437] <=  8'h00;      memory[32438] <=  8'h00;      memory[32439] <=  8'h00;      memory[32440] <=  8'h00;      memory[32441] <=  8'h00;      memory[32442] <=  8'h00;      memory[32443] <=  8'h00;      memory[32444] <=  8'h00;      memory[32445] <=  8'h00;      memory[32446] <=  8'h00;      memory[32447] <=  8'h00;      memory[32448] <=  8'h00;      memory[32449] <=  8'h00;      memory[32450] <=  8'h00;      memory[32451] <=  8'h00;      memory[32452] <=  8'h00;      memory[32453] <=  8'h00;      memory[32454] <=  8'h00;      memory[32455] <=  8'h00;      memory[32456] <=  8'h00;      memory[32457] <=  8'h00;      memory[32458] <=  8'h00;      memory[32459] <=  8'h00;      memory[32460] <=  8'h00;      memory[32461] <=  8'h00;      memory[32462] <=  8'h00;      memory[32463] <=  8'h00;      memory[32464] <=  8'h00;      memory[32465] <=  8'h00;      memory[32466] <=  8'h00;      memory[32467] <=  8'h00;      memory[32468] <=  8'h00;      memory[32469] <=  8'h00;      memory[32470] <=  8'h00;      memory[32471] <=  8'h00;      memory[32472] <=  8'h00;      memory[32473] <=  8'h00;      memory[32474] <=  8'h00;      memory[32475] <=  8'h00;      memory[32476] <=  8'h00;      memory[32477] <=  8'h00;      memory[32478] <=  8'h00;      memory[32479] <=  8'h00;      memory[32480] <=  8'h00;      memory[32481] <=  8'h00;      memory[32482] <=  8'h00;      memory[32483] <=  8'h00;      memory[32484] <=  8'h00;      memory[32485] <=  8'h00;      memory[32486] <=  8'h00;      memory[32487] <=  8'h00;      memory[32488] <=  8'h00;      memory[32489] <=  8'h00;      memory[32490] <=  8'h00;      memory[32491] <=  8'h00;      memory[32492] <=  8'h00;      memory[32493] <=  8'h00;      memory[32494] <=  8'h00;      memory[32495] <=  8'h00;      memory[32496] <=  8'h00;      memory[32497] <=  8'h00;      memory[32498] <=  8'h00;      memory[32499] <=  8'h00;      memory[32500] <=  8'h00;      memory[32501] <=  8'h00;      memory[32502] <=  8'h00;      memory[32503] <=  8'h00;      memory[32504] <=  8'h00;      memory[32505] <=  8'h00;      memory[32506] <=  8'h00;      memory[32507] <=  8'h00;      memory[32508] <=  8'h00;      memory[32509] <=  8'h00;      memory[32510] <=  8'h00;      memory[32511] <=  8'h00;      memory[32512] <=  8'h00;      memory[32513] <=  8'h00;      memory[32514] <=  8'h00;      memory[32515] <=  8'h00;      memory[32516] <=  8'h00;      memory[32517] <=  8'h00;      memory[32518] <=  8'h00;      memory[32519] <=  8'h00;      memory[32520] <=  8'h00;      memory[32521] <=  8'h00;      memory[32522] <=  8'h00;      memory[32523] <=  8'h00;      memory[32524] <=  8'h00;      memory[32525] <=  8'h00;      memory[32526] <=  8'h00;      memory[32527] <=  8'h00;      memory[32528] <=  8'h00;      memory[32529] <=  8'h00;      memory[32530] <=  8'h00;      memory[32531] <=  8'h00;      memory[32532] <=  8'h00;      memory[32533] <=  8'h00;      memory[32534] <=  8'h00;      memory[32535] <=  8'h00;      memory[32536] <=  8'h00;      memory[32537] <=  8'h00;      memory[32538] <=  8'h00;      memory[32539] <=  8'h00;      memory[32540] <=  8'h00;      memory[32541] <=  8'h00;      memory[32542] <=  8'h00;      memory[32543] <=  8'h00;      memory[32544] <=  8'h00;      memory[32545] <=  8'h00;      memory[32546] <=  8'h00;      memory[32547] <=  8'h00;      memory[32548] <=  8'h00;      memory[32549] <=  8'h00;      memory[32550] <=  8'h00;      memory[32551] <=  8'h00;      memory[32552] <=  8'h00;      memory[32553] <=  8'h00;      memory[32554] <=  8'h00;      memory[32555] <=  8'h00;      memory[32556] <=  8'h00;      memory[32557] <=  8'h00;      memory[32558] <=  8'h00;      memory[32559] <=  8'h00;      memory[32560] <=  8'h00;      memory[32561] <=  8'h00;      memory[32562] <=  8'h00;      memory[32563] <=  8'h00;      memory[32564] <=  8'h00;      memory[32565] <=  8'h00;      memory[32566] <=  8'h00;      memory[32567] <=  8'h00;      memory[32568] <=  8'h00;      memory[32569] <=  8'h00;      memory[32570] <=  8'h00;      memory[32571] <=  8'h00;      memory[32572] <=  8'h00;      memory[32573] <=  8'h00;      memory[32574] <=  8'h00;      memory[32575] <=  8'h00;      memory[32576] <=  8'h00;      memory[32577] <=  8'h00;      memory[32578] <=  8'h00;      memory[32579] <=  8'h00;      memory[32580] <=  8'h00;      memory[32581] <=  8'h00;      memory[32582] <=  8'h00;      memory[32583] <=  8'h00;      memory[32584] <=  8'h00;      memory[32585] <=  8'h00;      memory[32586] <=  8'h00;      memory[32587] <=  8'h00;      memory[32588] <=  8'h00;      memory[32589] <=  8'h00;      memory[32590] <=  8'h00;      memory[32591] <=  8'h00;      memory[32592] <=  8'h00;      memory[32593] <=  8'h00;      memory[32594] <=  8'h00;      memory[32595] <=  8'h00;      memory[32596] <=  8'h00;      memory[32597] <=  8'h00;      memory[32598] <=  8'h00;      memory[32599] <=  8'h00;      memory[32600] <=  8'h00;      memory[32601] <=  8'h00;      memory[32602] <=  8'h00;      memory[32603] <=  8'h00;      memory[32604] <=  8'h00;      memory[32605] <=  8'h00;      memory[32606] <=  8'h00;      memory[32607] <=  8'h00;      memory[32608] <=  8'h00;      memory[32609] <=  8'h00;      memory[32610] <=  8'h00;      memory[32611] <=  8'h00;      memory[32612] <=  8'h00;      memory[32613] <=  8'h00;      memory[32614] <=  8'h00;      memory[32615] <=  8'h00;      memory[32616] <=  8'h00;      memory[32617] <=  8'h00;      memory[32618] <=  8'h00;      memory[32619] <=  8'h00;      memory[32620] <=  8'h00;      memory[32621] <=  8'h00;      memory[32622] <=  8'h00;      memory[32623] <=  8'h00;      memory[32624] <=  8'h00;      memory[32625] <=  8'h00;      memory[32626] <=  8'h00;      memory[32627] <=  8'h00;      memory[32628] <=  8'h00;      memory[32629] <=  8'h00;      memory[32630] <=  8'h00;      memory[32631] <=  8'h00;      memory[32632] <=  8'h00;      memory[32633] <=  8'h00;      memory[32634] <=  8'h00;      memory[32635] <=  8'h00;      memory[32636] <=  8'h00;      memory[32637] <=  8'h00;      memory[32638] <=  8'h00;      memory[32639] <=  8'h00;      memory[32640] <=  8'h00;      memory[32641] <=  8'h00;      memory[32642] <=  8'h00;      memory[32643] <=  8'h00;      memory[32644] <=  8'h00;      memory[32645] <=  8'h00;      memory[32646] <=  8'h00;      memory[32647] <=  8'h00;      memory[32648] <=  8'h00;      memory[32649] <=  8'h00;      memory[32650] <=  8'h00;      memory[32651] <=  8'h00;      memory[32652] <=  8'h00;      memory[32653] <=  8'h00;      memory[32654] <=  8'h00;      memory[32655] <=  8'h00;      memory[32656] <=  8'h00;      memory[32657] <=  8'h00;      memory[32658] <=  8'h00;      memory[32659] <=  8'h00;      memory[32660] <=  8'h00;      memory[32661] <=  8'h00;      memory[32662] <=  8'h00;      memory[32663] <=  8'h00;      memory[32664] <=  8'h00;      memory[32665] <=  8'h00;      memory[32666] <=  8'h00;      memory[32667] <=  8'h00;      memory[32668] <=  8'h00;      memory[32669] <=  8'h00;      memory[32670] <=  8'h00;      memory[32671] <=  8'h00;      memory[32672] <=  8'h00;      memory[32673] <=  8'h00;      memory[32674] <=  8'h00;      memory[32675] <=  8'h00;      memory[32676] <=  8'h00;      memory[32677] <=  8'h00;      memory[32678] <=  8'h00;      memory[32679] <=  8'h00;      memory[32680] <=  8'h00;      memory[32681] <=  8'h00;      memory[32682] <=  8'h00;      memory[32683] <=  8'h00;      memory[32684] <=  8'h00;      memory[32685] <=  8'h00;      memory[32686] <=  8'h00;      memory[32687] <=  8'h00;      memory[32688] <=  8'h00;      memory[32689] <=  8'h00;      memory[32690] <=  8'h00;      memory[32691] <=  8'h00;      memory[32692] <=  8'h00;      memory[32693] <=  8'h00;      memory[32694] <=  8'h00;      memory[32695] <=  8'h00;      memory[32696] <=  8'h00;      memory[32697] <=  8'h00;      memory[32698] <=  8'h00;      memory[32699] <=  8'h00;      memory[32700] <=  8'h00;      memory[32701] <=  8'h00;      memory[32702] <=  8'h00;      memory[32703] <=  8'h00;      memory[32704] <=  8'h00;      memory[32705] <=  8'h00;      memory[32706] <=  8'h00;      memory[32707] <=  8'h00;      memory[32708] <=  8'h00;      memory[32709] <=  8'h00;      memory[32710] <=  8'h00;      memory[32711] <=  8'h00;      memory[32712] <=  8'h00;      memory[32713] <=  8'h00;      memory[32714] <=  8'h00;      memory[32715] <=  8'h00;      memory[32716] <=  8'h00;      memory[32717] <=  8'h00;      memory[32718] <=  8'h00;      memory[32719] <=  8'h00;      memory[32720] <=  8'h00;      memory[32721] <=  8'h00;      memory[32722] <=  8'h00;      memory[32723] <=  8'h00;      memory[32724] <=  8'h00;      memory[32725] <=  8'h00;      memory[32726] <=  8'h00;      memory[32727] <=  8'h00;      memory[32728] <=  8'h00;      memory[32729] <=  8'h00;      memory[32730] <=  8'h00;      memory[32731] <=  8'h00;      memory[32732] <=  8'h00;      memory[32733] <=  8'h00;      memory[32734] <=  8'h00;      memory[32735] <=  8'h00;      memory[32736] <=  8'h00;      memory[32737] <=  8'h00;      memory[32738] <=  8'h00;      memory[32739] <=  8'h00;      memory[32740] <=  8'h00;      memory[32741] <=  8'h00;      memory[32742] <=  8'h00;      memory[32743] <=  8'h00;      memory[32744] <=  8'h00;      memory[32745] <=  8'h00;      memory[32746] <=  8'h00;      memory[32747] <=  8'h00;      memory[32748] <=  8'h00;      memory[32749] <=  8'h00;      memory[32750] <=  8'h00;      memory[32751] <=  8'h00;      memory[32752] <=  8'h00;      memory[32753] <=  8'h00;      memory[32754] <=  8'h00;      memory[32755] <=  8'h00;      memory[32756] <=  8'h00;      memory[32757] <=  8'h00;      memory[32758] <=  8'h00;      memory[32759] <=  8'h00;      memory[32760] <=  8'h00;      memory[32761] <=  8'h00;      memory[32762] <=  8'h00;      memory[32763] <=  8'h00;      memory[32764] <=  8'h00;      memory[32765] <=  8'h00;      memory[32766] <=  8'h00;      memory[32767] <=  8'h00;      memory[32768] <=  8'h00;      memory[32769] <=  8'h00;      memory[32770] <=  8'h00;      memory[32771] <=  8'h00;      memory[32772] <=  8'h00;      memory[32773] <=  8'h00;      memory[32774] <=  8'h00;      memory[32775] <=  8'h00;      memory[32776] <=  8'h00;      memory[32777] <=  8'h00;      memory[32778] <=  8'h00;      memory[32779] <=  8'h00;      memory[32780] <=  8'h00;      memory[32781] <=  8'h00;      memory[32782] <=  8'h00;      memory[32783] <=  8'h00;      memory[32784] <=  8'h00;      memory[32785] <=  8'h00;      memory[32786] <=  8'h00;      memory[32787] <=  8'h00;      memory[32788] <=  8'h00;      memory[32789] <=  8'h00;      memory[32790] <=  8'h00;      memory[32791] <=  8'h00;      memory[32792] <=  8'h00;      memory[32793] <=  8'h00;      memory[32794] <=  8'h00;      memory[32795] <=  8'h00;      memory[32796] <=  8'h00;      memory[32797] <=  8'h00;      memory[32798] <=  8'h00;      memory[32799] <=  8'h00;      memory[32800] <=  8'h00;      memory[32801] <=  8'h00;      memory[32802] <=  8'h00;      memory[32803] <=  8'h00;      memory[32804] <=  8'h00;      memory[32805] <=  8'h00;      memory[32806] <=  8'h00;      memory[32807] <=  8'h00;      memory[32808] <=  8'h00;      memory[32809] <=  8'h00;      memory[32810] <=  8'h00;      memory[32811] <=  8'h00;      memory[32812] <=  8'h00;      memory[32813] <=  8'h00;      memory[32814] <=  8'h00;      memory[32815] <=  8'h00;      memory[32816] <=  8'h00;      memory[32817] <=  8'h00;      memory[32818] <=  8'h00;      memory[32819] <=  8'h00;      memory[32820] <=  8'h00;      memory[32821] <=  8'h00;      memory[32822] <=  8'h00;      memory[32823] <=  8'h00;      memory[32824] <=  8'h00;      memory[32825] <=  8'h00;      memory[32826] <=  8'h00;      memory[32827] <=  8'h00;      memory[32828] <=  8'h00;      memory[32829] <=  8'h00;      memory[32830] <=  8'h00;      memory[32831] <=  8'h00;      memory[32832] <=  8'h00;      memory[32833] <=  8'h00;      memory[32834] <=  8'h00;      memory[32835] <=  8'h00;      memory[32836] <=  8'h00;      memory[32837] <=  8'h00;      memory[32838] <=  8'h00;      memory[32839] <=  8'h00;      memory[32840] <=  8'h00;      memory[32841] <=  8'h00;      memory[32842] <=  8'h00;      memory[32843] <=  8'h00;      memory[32844] <=  8'h00;      memory[32845] <=  8'h00;      memory[32846] <=  8'h00;      memory[32847] <=  8'h00;      memory[32848] <=  8'h00;      memory[32849] <=  8'h00;      memory[32850] <=  8'h00;      memory[32851] <=  8'h00;      memory[32852] <=  8'h00;      memory[32853] <=  8'h00;      memory[32854] <=  8'h00;      memory[32855] <=  8'h00;      memory[32856] <=  8'h00;      memory[32857] <=  8'h00;      memory[32858] <=  8'h00;      memory[32859] <=  8'h00;      memory[32860] <=  8'h00;      memory[32861] <=  8'h00;      memory[32862] <=  8'h00;      memory[32863] <=  8'h00;      memory[32864] <=  8'h00;      memory[32865] <=  8'h00;      memory[32866] <=  8'h00;      memory[32867] <=  8'h00;      memory[32868] <=  8'h00;      memory[32869] <=  8'h00;      memory[32870] <=  8'h00;      memory[32871] <=  8'h00;      memory[32872] <=  8'h00;      memory[32873] <=  8'h00;      memory[32874] <=  8'h00;      memory[32875] <=  8'h00;      memory[32876] <=  8'h00;      memory[32877] <=  8'h00;      memory[32878] <=  8'h00;      memory[32879] <=  8'h00;      memory[32880] <=  8'h00;      memory[32881] <=  8'h00;      memory[32882] <=  8'h00;      memory[32883] <=  8'h00;      memory[32884] <=  8'h00;      memory[32885] <=  8'h00;      memory[32886] <=  8'h00;      memory[32887] <=  8'h00;      memory[32888] <=  8'h00;      memory[32889] <=  8'h00;      memory[32890] <=  8'h00;      memory[32891] <=  8'h00;      memory[32892] <=  8'h00;      memory[32893] <=  8'h00;      memory[32894] <=  8'h00;      memory[32895] <=  8'h00;      memory[32896] <=  8'h00;      memory[32897] <=  8'h00;      memory[32898] <=  8'h00;      memory[32899] <=  8'h00;      memory[32900] <=  8'h00;      memory[32901] <=  8'h00;      memory[32902] <=  8'h00;      memory[32903] <=  8'h00;      memory[32904] <=  8'h00;      memory[32905] <=  8'h00;      memory[32906] <=  8'h00;      memory[32907] <=  8'h00;      memory[32908] <=  8'h00;      memory[32909] <=  8'h00;      memory[32910] <=  8'h00;      memory[32911] <=  8'h00;      memory[32912] <=  8'h00;      memory[32913] <=  8'h00;      memory[32914] <=  8'h00;      memory[32915] <=  8'h00;      memory[32916] <=  8'h00;      memory[32917] <=  8'h00;      memory[32918] <=  8'h00;      memory[32919] <=  8'h00;      memory[32920] <=  8'h00;      memory[32921] <=  8'h00;      memory[32922] <=  8'h00;      memory[32923] <=  8'h00;      memory[32924] <=  8'h00;      memory[32925] <=  8'h00;      memory[32926] <=  8'h00;      memory[32927] <=  8'h00;      memory[32928] <=  8'h00;      memory[32929] <=  8'h00;      memory[32930] <=  8'h00;      memory[32931] <=  8'h00;      memory[32932] <=  8'h00;      memory[32933] <=  8'h00;      memory[32934] <=  8'h00;      memory[32935] <=  8'h00;      memory[32936] <=  8'h00;      memory[32937] <=  8'h00;      memory[32938] <=  8'h00;      memory[32939] <=  8'h00;      memory[32940] <=  8'h00;      memory[32941] <=  8'h00;      memory[32942] <=  8'h00;      memory[32943] <=  8'h00;      memory[32944] <=  8'h00;      memory[32945] <=  8'h00;      memory[32946] <=  8'h00;      memory[32947] <=  8'h00;      memory[32948] <=  8'h00;      memory[32949] <=  8'h00;      memory[32950] <=  8'h00;      memory[32951] <=  8'h00;      memory[32952] <=  8'h00;      memory[32953] <=  8'h00;      memory[32954] <=  8'h00;      memory[32955] <=  8'h00;      memory[32956] <=  8'h00;      memory[32957] <=  8'h00;      memory[32958] <=  8'h00;      memory[32959] <=  8'h00;      memory[32960] <=  8'h00;      memory[32961] <=  8'h00;      memory[32962] <=  8'h00;      memory[32963] <=  8'h00;      memory[32964] <=  8'h00;      memory[32965] <=  8'h00;      memory[32966] <=  8'h00;      memory[32967] <=  8'h00;      memory[32968] <=  8'h00;      memory[32969] <=  8'h00;      memory[32970] <=  8'h00;      memory[32971] <=  8'h00;      memory[32972] <=  8'h00;      memory[32973] <=  8'h00;      memory[32974] <=  8'h00;      memory[32975] <=  8'h00;      memory[32976] <=  8'h00;      memory[32977] <=  8'h00;      memory[32978] <=  8'h00;      memory[32979] <=  8'h00;      memory[32980] <=  8'h00;      memory[32981] <=  8'h00;      memory[32982] <=  8'h00;      memory[32983] <=  8'h00;      memory[32984] <=  8'h00;      memory[32985] <=  8'h00;      memory[32986] <=  8'h00;      memory[32987] <=  8'h00;      memory[32988] <=  8'h00;      memory[32989] <=  8'h00;      memory[32990] <=  8'h00;      memory[32991] <=  8'h00;      memory[32992] <=  8'h00;      memory[32993] <=  8'h00;      memory[32994] <=  8'h00;      memory[32995] <=  8'h00;      memory[32996] <=  8'h00;      memory[32997] <=  8'h00;      memory[32998] <=  8'h00;      memory[32999] <=  8'h00;      memory[33000] <=  8'h00;      memory[33001] <=  8'h00;      memory[33002] <=  8'h00;      memory[33003] <=  8'h00;      memory[33004] <=  8'h00;      memory[33005] <=  8'h00;      memory[33006] <=  8'h00;      memory[33007] <=  8'h00;      memory[33008] <=  8'h00;      memory[33009] <=  8'h00;      memory[33010] <=  8'h00;      memory[33011] <=  8'h00;      memory[33012] <=  8'h00;      memory[33013] <=  8'h00;      memory[33014] <=  8'h00;      memory[33015] <=  8'h00;      memory[33016] <=  8'h00;      memory[33017] <=  8'h00;      memory[33018] <=  8'h00;      memory[33019] <=  8'h00;      memory[33020] <=  8'h00;      memory[33021] <=  8'h00;      memory[33022] <=  8'h00;      memory[33023] <=  8'h00;      memory[33024] <=  8'h00;      memory[33025] <=  8'h00;      memory[33026] <=  8'h00;      memory[33027] <=  8'h00;      memory[33028] <=  8'h00;      memory[33029] <=  8'h00;      memory[33030] <=  8'h00;      memory[33031] <=  8'h00;      memory[33032] <=  8'h00;      memory[33033] <=  8'h00;      memory[33034] <=  8'h00;      memory[33035] <=  8'h00;      memory[33036] <=  8'h00;      memory[33037] <=  8'h00;      memory[33038] <=  8'h00;      memory[33039] <=  8'h00;      memory[33040] <=  8'h00;      memory[33041] <=  8'h00;      memory[33042] <=  8'h00;      memory[33043] <=  8'h00;      memory[33044] <=  8'h00;      memory[33045] <=  8'h00;      memory[33046] <=  8'h00;      memory[33047] <=  8'h00;      memory[33048] <=  8'h00;      memory[33049] <=  8'h00;      memory[33050] <=  8'h00;      memory[33051] <=  8'h00;      memory[33052] <=  8'h00;      memory[33053] <=  8'h00;      memory[33054] <=  8'h00;      memory[33055] <=  8'h00;      memory[33056] <=  8'h00;      memory[33057] <=  8'h00;      memory[33058] <=  8'h00;      memory[33059] <=  8'h00;      memory[33060] <=  8'h00;      memory[33061] <=  8'h00;      memory[33062] <=  8'h00;      memory[33063] <=  8'h00;      memory[33064] <=  8'h00;      memory[33065] <=  8'h00;      memory[33066] <=  8'h00;      memory[33067] <=  8'h00;      memory[33068] <=  8'h00;      memory[33069] <=  8'h00;      memory[33070] <=  8'h00;      memory[33071] <=  8'h00;      memory[33072] <=  8'h00;      memory[33073] <=  8'h00;      memory[33074] <=  8'h00;      memory[33075] <=  8'h00;      memory[33076] <=  8'h00;      memory[33077] <=  8'h00;      memory[33078] <=  8'h00;      memory[33079] <=  8'h00;      memory[33080] <=  8'h00;      memory[33081] <=  8'h00;      memory[33082] <=  8'h00;      memory[33083] <=  8'h00;      memory[33084] <=  8'h00;      memory[33085] <=  8'h00;      memory[33086] <=  8'h00;      memory[33087] <=  8'h00;      memory[33088] <=  8'h00;      memory[33089] <=  8'h00;      memory[33090] <=  8'h00;      memory[33091] <=  8'h00;      memory[33092] <=  8'h00;      memory[33093] <=  8'h00;      memory[33094] <=  8'h00;      memory[33095] <=  8'h00;      memory[33096] <=  8'h00;      memory[33097] <=  8'h00;      memory[33098] <=  8'h00;      memory[33099] <=  8'h00;      memory[33100] <=  8'h00;      memory[33101] <=  8'h00;      memory[33102] <=  8'h00;      memory[33103] <=  8'h00;      memory[33104] <=  8'h00;      memory[33105] <=  8'h00;      memory[33106] <=  8'h00;      memory[33107] <=  8'h00;      memory[33108] <=  8'h00;      memory[33109] <=  8'h00;      memory[33110] <=  8'h00;      memory[33111] <=  8'h00;      memory[33112] <=  8'h00;      memory[33113] <=  8'h00;      memory[33114] <=  8'h00;      memory[33115] <=  8'h00;      memory[33116] <=  8'h00;      memory[33117] <=  8'h00;      memory[33118] <=  8'h00;      memory[33119] <=  8'h00;      memory[33120] <=  8'h00;      memory[33121] <=  8'h00;      memory[33122] <=  8'h00;      memory[33123] <=  8'h00;      memory[33124] <=  8'h00;      memory[33125] <=  8'h00;      memory[33126] <=  8'h00;      memory[33127] <=  8'h00;      memory[33128] <=  8'h00;      memory[33129] <=  8'h00;      memory[33130] <=  8'h00;      memory[33131] <=  8'h00;      memory[33132] <=  8'h00;      memory[33133] <=  8'h00;      memory[33134] <=  8'h00;      memory[33135] <=  8'h00;      memory[33136] <=  8'h00;      memory[33137] <=  8'h00;      memory[33138] <=  8'h00;      memory[33139] <=  8'h00;      memory[33140] <=  8'h00;      memory[33141] <=  8'h00;      memory[33142] <=  8'h00;      memory[33143] <=  8'h00;      memory[33144] <=  8'h00;      memory[33145] <=  8'h00;      memory[33146] <=  8'h00;      memory[33147] <=  8'h00;      memory[33148] <=  8'h00;      memory[33149] <=  8'h00;      memory[33150] <=  8'h00;      memory[33151] <=  8'h00;      memory[33152] <=  8'h00;      memory[33153] <=  8'h00;      memory[33154] <=  8'h00;      memory[33155] <=  8'h00;      memory[33156] <=  8'h00;      memory[33157] <=  8'h00;      memory[33158] <=  8'h00;      memory[33159] <=  8'h00;      memory[33160] <=  8'h00;      memory[33161] <=  8'h00;      memory[33162] <=  8'h00;      memory[33163] <=  8'h00;      memory[33164] <=  8'h00;      memory[33165] <=  8'h00;      memory[33166] <=  8'h00;      memory[33167] <=  8'h00;      memory[33168] <=  8'h00;      memory[33169] <=  8'h00;      memory[33170] <=  8'h00;      memory[33171] <=  8'h00;      memory[33172] <=  8'h00;      memory[33173] <=  8'h00;      memory[33174] <=  8'h00;      memory[33175] <=  8'h00;      memory[33176] <=  8'h00;      memory[33177] <=  8'h00;      memory[33178] <=  8'h00;      memory[33179] <=  8'h00;      memory[33180] <=  8'h00;      memory[33181] <=  8'h00;      memory[33182] <=  8'h00;      memory[33183] <=  8'h00;      memory[33184] <=  8'h00;      memory[33185] <=  8'h00;      memory[33186] <=  8'h00;      memory[33187] <=  8'h00;      memory[33188] <=  8'h00;      memory[33189] <=  8'h00;      memory[33190] <=  8'h00;      memory[33191] <=  8'h00;      memory[33192] <=  8'h00;      memory[33193] <=  8'h00;      memory[33194] <=  8'h00;      memory[33195] <=  8'h00;      memory[33196] <=  8'h00;      memory[33197] <=  8'h00;      memory[33198] <=  8'h00;      memory[33199] <=  8'h00;      memory[33200] <=  8'h00;      memory[33201] <=  8'h00;      memory[33202] <=  8'h00;      memory[33203] <=  8'h00;      memory[33204] <=  8'h00;      memory[33205] <=  8'h00;      memory[33206] <=  8'h00;      memory[33207] <=  8'h00;      memory[33208] <=  8'h00;      memory[33209] <=  8'h00;      memory[33210] <=  8'h00;      memory[33211] <=  8'h00;      memory[33212] <=  8'h00;      memory[33213] <=  8'h00;      memory[33214] <=  8'h00;      memory[33215] <=  8'h00;      memory[33216] <=  8'h00;      memory[33217] <=  8'h00;      memory[33218] <=  8'h00;      memory[33219] <=  8'h00;      memory[33220] <=  8'h00;      memory[33221] <=  8'h00;      memory[33222] <=  8'h00;      memory[33223] <=  8'h00;      memory[33224] <=  8'h00;      memory[33225] <=  8'h00;      memory[33226] <=  8'h00;      memory[33227] <=  8'h00;      memory[33228] <=  8'h00;      memory[33229] <=  8'h00;      memory[33230] <=  8'h00;      memory[33231] <=  8'h00;      memory[33232] <=  8'h00;      memory[33233] <=  8'h00;      memory[33234] <=  8'h00;      memory[33235] <=  8'h00;      memory[33236] <=  8'h00;      memory[33237] <=  8'h00;      memory[33238] <=  8'h00;      memory[33239] <=  8'h00;      memory[33240] <=  8'h00;      memory[33241] <=  8'h00;      memory[33242] <=  8'h00;      memory[33243] <=  8'h00;      memory[33244] <=  8'h00;      memory[33245] <=  8'h00;      memory[33246] <=  8'h00;      memory[33247] <=  8'h00;      memory[33248] <=  8'h00;      memory[33249] <=  8'h00;      memory[33250] <=  8'h00;      memory[33251] <=  8'h00;      memory[33252] <=  8'h00;      memory[33253] <=  8'h00;      memory[33254] <=  8'h00;      memory[33255] <=  8'h00;      memory[33256] <=  8'h00;      memory[33257] <=  8'h00;      memory[33258] <=  8'h00;      memory[33259] <=  8'h00;      memory[33260] <=  8'h00;      memory[33261] <=  8'h00;      memory[33262] <=  8'h00;      memory[33263] <=  8'h00;      memory[33264] <=  8'h00;      memory[33265] <=  8'h00;      memory[33266] <=  8'h00;      memory[33267] <=  8'h00;      memory[33268] <=  8'h00;      memory[33269] <=  8'h00;      memory[33270] <=  8'h00;      memory[33271] <=  8'h00;      memory[33272] <=  8'h00;      memory[33273] <=  8'h00;      memory[33274] <=  8'h00;      memory[33275] <=  8'h00;      memory[33276] <=  8'h00;      memory[33277] <=  8'h00;      memory[33278] <=  8'h00;      memory[33279] <=  8'h00;      memory[33280] <=  8'h00;      memory[33281] <=  8'h00;      memory[33282] <=  8'h00;      memory[33283] <=  8'h00;      memory[33284] <=  8'h00;      memory[33285] <=  8'h00;      memory[33286] <=  8'h00;      memory[33287] <=  8'h00;      memory[33288] <=  8'h00;      memory[33289] <=  8'h00;      memory[33290] <=  8'h00;      memory[33291] <=  8'h00;      memory[33292] <=  8'h00;      memory[33293] <=  8'h00;      memory[33294] <=  8'h00;      memory[33295] <=  8'h00;      memory[33296] <=  8'h00;      memory[33297] <=  8'h00;      memory[33298] <=  8'h00;      memory[33299] <=  8'h00;      memory[33300] <=  8'h00;      memory[33301] <=  8'h00;      memory[33302] <=  8'h00;      memory[33303] <=  8'h00;      memory[33304] <=  8'h00;      memory[33305] <=  8'h00;      memory[33306] <=  8'h00;      memory[33307] <=  8'h00;      memory[33308] <=  8'h00;      memory[33309] <=  8'h00;      memory[33310] <=  8'h00;      memory[33311] <=  8'h00;      memory[33312] <=  8'h00;      memory[33313] <=  8'h00;      memory[33314] <=  8'h00;      memory[33315] <=  8'h00;      memory[33316] <=  8'h00;      memory[33317] <=  8'h00;      memory[33318] <=  8'h00;      memory[33319] <=  8'h00;      memory[33320] <=  8'h00;      memory[33321] <=  8'h00;      memory[33322] <=  8'h00;      memory[33323] <=  8'h00;      memory[33324] <=  8'h00;      memory[33325] <=  8'h00;      memory[33326] <=  8'h00;      memory[33327] <=  8'h00;      memory[33328] <=  8'h00;      memory[33329] <=  8'h00;      memory[33330] <=  8'h00;      memory[33331] <=  8'h00;      memory[33332] <=  8'h00;      memory[33333] <=  8'h00;      memory[33334] <=  8'h00;      memory[33335] <=  8'h00;      memory[33336] <=  8'h00;      memory[33337] <=  8'h00;      memory[33338] <=  8'h00;      memory[33339] <=  8'h00;      memory[33340] <=  8'h00;      memory[33341] <=  8'h00;      memory[33342] <=  8'h00;      memory[33343] <=  8'h00;      memory[33344] <=  8'h00;      memory[33345] <=  8'h00;      memory[33346] <=  8'h00;      memory[33347] <=  8'h00;      memory[33348] <=  8'h00;      memory[33349] <=  8'h00;      memory[33350] <=  8'h00;      memory[33351] <=  8'h00;      memory[33352] <=  8'h00;      memory[33353] <=  8'h00;      memory[33354] <=  8'h00;      memory[33355] <=  8'h00;      memory[33356] <=  8'h00;      memory[33357] <=  8'h00;      memory[33358] <=  8'h00;      memory[33359] <=  8'h00;      memory[33360] <=  8'h00;      memory[33361] <=  8'h00;      memory[33362] <=  8'h00;      memory[33363] <=  8'h00;      memory[33364] <=  8'h00;      memory[33365] <=  8'h00;      memory[33366] <=  8'h00;      memory[33367] <=  8'h00;      memory[33368] <=  8'h00;      memory[33369] <=  8'h00;      memory[33370] <=  8'h00;      memory[33371] <=  8'h00;      memory[33372] <=  8'h00;      memory[33373] <=  8'h00;      memory[33374] <=  8'h00;      memory[33375] <=  8'h00;      memory[33376] <=  8'h00;      memory[33377] <=  8'h00;      memory[33378] <=  8'h00;      memory[33379] <=  8'h00;      memory[33380] <=  8'h00;      memory[33381] <=  8'h00;      memory[33382] <=  8'h00;      memory[33383] <=  8'h00;      memory[33384] <=  8'h00;      memory[33385] <=  8'h00;      memory[33386] <=  8'h00;      memory[33387] <=  8'h00;      memory[33388] <=  8'h00;      memory[33389] <=  8'h00;      memory[33390] <=  8'h00;      memory[33391] <=  8'h00;      memory[33392] <=  8'h00;      memory[33393] <=  8'h00;      memory[33394] <=  8'h00;      memory[33395] <=  8'h00;      memory[33396] <=  8'h00;      memory[33397] <=  8'h00;      memory[33398] <=  8'h00;      memory[33399] <=  8'h00;      memory[33400] <=  8'h00;      memory[33401] <=  8'h00;      memory[33402] <=  8'h00;      memory[33403] <=  8'h00;      memory[33404] <=  8'h00;      memory[33405] <=  8'h00;      memory[33406] <=  8'h00;      memory[33407] <=  8'h00;      memory[33408] <=  8'h00;      memory[33409] <=  8'h00;      memory[33410] <=  8'h00;      memory[33411] <=  8'h00;      memory[33412] <=  8'h00;      memory[33413] <=  8'h00;      memory[33414] <=  8'h00;      memory[33415] <=  8'h00;      memory[33416] <=  8'h00;      memory[33417] <=  8'h00;      memory[33418] <=  8'h00;      memory[33419] <=  8'h00;      memory[33420] <=  8'h00;      memory[33421] <=  8'h00;      memory[33422] <=  8'h00;      memory[33423] <=  8'h00;      memory[33424] <=  8'h00;      memory[33425] <=  8'h00;      memory[33426] <=  8'h00;      memory[33427] <=  8'h00;      memory[33428] <=  8'h00;      memory[33429] <=  8'h00;      memory[33430] <=  8'h00;      memory[33431] <=  8'h00;      memory[33432] <=  8'h00;      memory[33433] <=  8'h00;      memory[33434] <=  8'h00;      memory[33435] <=  8'h00;      memory[33436] <=  8'h00;      memory[33437] <=  8'h00;      memory[33438] <=  8'h00;      memory[33439] <=  8'h00;      memory[33440] <=  8'h00;      memory[33441] <=  8'h00;      memory[33442] <=  8'h00;      memory[33443] <=  8'h00;      memory[33444] <=  8'h00;      memory[33445] <=  8'h00;      memory[33446] <=  8'h00;      memory[33447] <=  8'h00;      memory[33448] <=  8'h00;      memory[33449] <=  8'h00;      memory[33450] <=  8'h00;      memory[33451] <=  8'h00;      memory[33452] <=  8'h00;      memory[33453] <=  8'h00;      memory[33454] <=  8'h00;      memory[33455] <=  8'h00;      memory[33456] <=  8'h00;      memory[33457] <=  8'h00;      memory[33458] <=  8'h00;      memory[33459] <=  8'h00;      memory[33460] <=  8'h00;      memory[33461] <=  8'h00;      memory[33462] <=  8'h00;      memory[33463] <=  8'h00;      memory[33464] <=  8'h00;      memory[33465] <=  8'h00;      memory[33466] <=  8'h00;      memory[33467] <=  8'h00;      memory[33468] <=  8'h00;      memory[33469] <=  8'h00;      memory[33470] <=  8'h00;      memory[33471] <=  8'h00;      memory[33472] <=  8'h00;      memory[33473] <=  8'h00;      memory[33474] <=  8'h00;      memory[33475] <=  8'h00;      memory[33476] <=  8'h00;      memory[33477] <=  8'h00;      memory[33478] <=  8'h00;      memory[33479] <=  8'h00;      memory[33480] <=  8'h00;      memory[33481] <=  8'h00;      memory[33482] <=  8'h00;      memory[33483] <=  8'h00;      memory[33484] <=  8'h00;      memory[33485] <=  8'h00;      memory[33486] <=  8'h00;      memory[33487] <=  8'h00;      memory[33488] <=  8'h00;      memory[33489] <=  8'h00;      memory[33490] <=  8'h00;      memory[33491] <=  8'h00;      memory[33492] <=  8'h00;      memory[33493] <=  8'h00;      memory[33494] <=  8'h00;      memory[33495] <=  8'h00;      memory[33496] <=  8'h00;      memory[33497] <=  8'h00;      memory[33498] <=  8'h00;      memory[33499] <=  8'h00;      memory[33500] <=  8'h00;      memory[33501] <=  8'h00;      memory[33502] <=  8'h00;      memory[33503] <=  8'h00;      memory[33504] <=  8'h00;      memory[33505] <=  8'h00;      memory[33506] <=  8'h00;      memory[33507] <=  8'h00;      memory[33508] <=  8'h00;      memory[33509] <=  8'h00;      memory[33510] <=  8'h00;      memory[33511] <=  8'h00;      memory[33512] <=  8'h00;      memory[33513] <=  8'h00;      memory[33514] <=  8'h00;      memory[33515] <=  8'h00;      memory[33516] <=  8'h00;      memory[33517] <=  8'h00;      memory[33518] <=  8'h00;      memory[33519] <=  8'h00;      memory[33520] <=  8'h00;      memory[33521] <=  8'h00;      memory[33522] <=  8'h00;      memory[33523] <=  8'h00;      memory[33524] <=  8'h00;      memory[33525] <=  8'h00;      memory[33526] <=  8'h00;      memory[33527] <=  8'h00;      memory[33528] <=  8'h00;      memory[33529] <=  8'h00;      memory[33530] <=  8'h00;      memory[33531] <=  8'h00;      memory[33532] <=  8'h00;      memory[33533] <=  8'h00;      memory[33534] <=  8'h00;      memory[33535] <=  8'h00;      memory[33536] <=  8'h00;      memory[33537] <=  8'h00;      memory[33538] <=  8'h00;      memory[33539] <=  8'h00;      memory[33540] <=  8'h00;      memory[33541] <=  8'h00;      memory[33542] <=  8'h00;      memory[33543] <=  8'h00;      memory[33544] <=  8'h00;      memory[33545] <=  8'h00;      memory[33546] <=  8'h00;      memory[33547] <=  8'h00;      memory[33548] <=  8'h00;      memory[33549] <=  8'h00;      memory[33550] <=  8'h00;      memory[33551] <=  8'h00;      memory[33552] <=  8'h00;      memory[33553] <=  8'h00;      memory[33554] <=  8'h00;      memory[33555] <=  8'h00;      memory[33556] <=  8'h00;      memory[33557] <=  8'h00;      memory[33558] <=  8'h00;      memory[33559] <=  8'h00;      memory[33560] <=  8'h00;      memory[33561] <=  8'h00;      memory[33562] <=  8'h00;      memory[33563] <=  8'h00;      memory[33564] <=  8'h00;      memory[33565] <=  8'h00;      memory[33566] <=  8'h00;      memory[33567] <=  8'h00;      memory[33568] <=  8'h00;      memory[33569] <=  8'h00;      memory[33570] <=  8'h00;      memory[33571] <=  8'h00;      memory[33572] <=  8'h00;      memory[33573] <=  8'h00;      memory[33574] <=  8'h00;      memory[33575] <=  8'h00;      memory[33576] <=  8'h00;      memory[33577] <=  8'h00;      memory[33578] <=  8'h00;      memory[33579] <=  8'h00;      memory[33580] <=  8'h00;      memory[33581] <=  8'h00;      memory[33582] <=  8'h00;      memory[33583] <=  8'h00;      memory[33584] <=  8'h00;      memory[33585] <=  8'h00;      memory[33586] <=  8'h00;      memory[33587] <=  8'h00;      memory[33588] <=  8'h00;      memory[33589] <=  8'h00;      memory[33590] <=  8'h00;      memory[33591] <=  8'h00;      memory[33592] <=  8'h00;      memory[33593] <=  8'h00;      memory[33594] <=  8'h00;      memory[33595] <=  8'h00;      memory[33596] <=  8'h00;      memory[33597] <=  8'h00;      memory[33598] <=  8'h00;      memory[33599] <=  8'h00;      memory[33600] <=  8'h00;      memory[33601] <=  8'h00;      memory[33602] <=  8'h00;      memory[33603] <=  8'h00;      memory[33604] <=  8'h00;      memory[33605] <=  8'h00;      memory[33606] <=  8'h00;      memory[33607] <=  8'h00;      memory[33608] <=  8'h00;      memory[33609] <=  8'h00;      memory[33610] <=  8'h00;      memory[33611] <=  8'h00;      memory[33612] <=  8'h00;      memory[33613] <=  8'h00;      memory[33614] <=  8'h00;      memory[33615] <=  8'h00;      memory[33616] <=  8'h00;      memory[33617] <=  8'h00;      memory[33618] <=  8'h00;      memory[33619] <=  8'h00;      memory[33620] <=  8'h00;      memory[33621] <=  8'h00;      memory[33622] <=  8'h00;      memory[33623] <=  8'h00;      memory[33624] <=  8'h00;      memory[33625] <=  8'h00;      memory[33626] <=  8'h00;      memory[33627] <=  8'h00;      memory[33628] <=  8'h00;      memory[33629] <=  8'h00;      memory[33630] <=  8'h00;      memory[33631] <=  8'h00;      memory[33632] <=  8'h00;      memory[33633] <=  8'h00;      memory[33634] <=  8'h00;      memory[33635] <=  8'h00;      memory[33636] <=  8'h00;      memory[33637] <=  8'h00;      memory[33638] <=  8'h00;      memory[33639] <=  8'h00;      memory[33640] <=  8'h00;      memory[33641] <=  8'h00;      memory[33642] <=  8'h00;      memory[33643] <=  8'h00;      memory[33644] <=  8'h00;      memory[33645] <=  8'h00;      memory[33646] <=  8'h00;      memory[33647] <=  8'h00;      memory[33648] <=  8'h00;      memory[33649] <=  8'h00;      memory[33650] <=  8'h00;      memory[33651] <=  8'h00;      memory[33652] <=  8'h00;      memory[33653] <=  8'h00;      memory[33654] <=  8'h00;      memory[33655] <=  8'h00;      memory[33656] <=  8'h00;      memory[33657] <=  8'h00;      memory[33658] <=  8'h00;      memory[33659] <=  8'h00;      memory[33660] <=  8'h00;      memory[33661] <=  8'h00;      memory[33662] <=  8'h00;      memory[33663] <=  8'h00;      memory[33664] <=  8'h00;      memory[33665] <=  8'h00;      memory[33666] <=  8'h00;      memory[33667] <=  8'h00;      memory[33668] <=  8'h00;      memory[33669] <=  8'h00;      memory[33670] <=  8'h00;      memory[33671] <=  8'h00;      memory[33672] <=  8'h00;      memory[33673] <=  8'h00;      memory[33674] <=  8'h00;      memory[33675] <=  8'h00;      memory[33676] <=  8'h00;      memory[33677] <=  8'h00;      memory[33678] <=  8'h00;      memory[33679] <=  8'h00;      memory[33680] <=  8'h00;      memory[33681] <=  8'h00;      memory[33682] <=  8'h00;      memory[33683] <=  8'h00;      memory[33684] <=  8'h00;      memory[33685] <=  8'h00;      memory[33686] <=  8'h00;      memory[33687] <=  8'h00;      memory[33688] <=  8'h00;      memory[33689] <=  8'h00;      memory[33690] <=  8'h00;      memory[33691] <=  8'h00;      memory[33692] <=  8'h00;      memory[33693] <=  8'h00;      memory[33694] <=  8'h00;      memory[33695] <=  8'h00;      memory[33696] <=  8'h00;      memory[33697] <=  8'h00;      memory[33698] <=  8'h00;      memory[33699] <=  8'h00;      memory[33700] <=  8'h00;      memory[33701] <=  8'h00;      memory[33702] <=  8'h00;      memory[33703] <=  8'h00;      memory[33704] <=  8'h00;      memory[33705] <=  8'h00;      memory[33706] <=  8'h00;      memory[33707] <=  8'h00;      memory[33708] <=  8'h00;      memory[33709] <=  8'h00;      memory[33710] <=  8'h00;      memory[33711] <=  8'h00;      memory[33712] <=  8'h00;      memory[33713] <=  8'h00;      memory[33714] <=  8'h00;      memory[33715] <=  8'h00;      memory[33716] <=  8'h00;      memory[33717] <=  8'h00;      memory[33718] <=  8'h00;      memory[33719] <=  8'h00;      memory[33720] <=  8'h00;      memory[33721] <=  8'h00;      memory[33722] <=  8'h00;      memory[33723] <=  8'h00;      memory[33724] <=  8'h00;      memory[33725] <=  8'h00;      memory[33726] <=  8'h00;      memory[33727] <=  8'h00;      memory[33728] <=  8'h00;      memory[33729] <=  8'h00;      memory[33730] <=  8'h00;      memory[33731] <=  8'h00;      memory[33732] <=  8'h00;      memory[33733] <=  8'h00;      memory[33734] <=  8'h00;      memory[33735] <=  8'h00;      memory[33736] <=  8'h00;      memory[33737] <=  8'h00;      memory[33738] <=  8'h00;      memory[33739] <=  8'h00;      memory[33740] <=  8'h00;      memory[33741] <=  8'h00;      memory[33742] <=  8'h00;      memory[33743] <=  8'h00;      memory[33744] <=  8'h00;      memory[33745] <=  8'h00;      memory[33746] <=  8'h00;      memory[33747] <=  8'h00;      memory[33748] <=  8'h00;      memory[33749] <=  8'h00;      memory[33750] <=  8'h00;      memory[33751] <=  8'h00;      memory[33752] <=  8'h00;      memory[33753] <=  8'h00;      memory[33754] <=  8'h00;      memory[33755] <=  8'h00;      memory[33756] <=  8'h00;      memory[33757] <=  8'h00;      memory[33758] <=  8'h00;      memory[33759] <=  8'h00;      memory[33760] <=  8'h00;      memory[33761] <=  8'h00;      memory[33762] <=  8'h00;      memory[33763] <=  8'h00;      memory[33764] <=  8'h00;      memory[33765] <=  8'h00;      memory[33766] <=  8'h00;      memory[33767] <=  8'h00;      memory[33768] <=  8'h00;      memory[33769] <=  8'h00;      memory[33770] <=  8'h00;      memory[33771] <=  8'h00;      memory[33772] <=  8'h00;      memory[33773] <=  8'h00;      memory[33774] <=  8'h00;      memory[33775] <=  8'h00;      memory[33776] <=  8'h00;      memory[33777] <=  8'h00;      memory[33778] <=  8'h00;      memory[33779] <=  8'h00;      memory[33780] <=  8'h00;      memory[33781] <=  8'h00;      memory[33782] <=  8'h00;      memory[33783] <=  8'h00;      memory[33784] <=  8'h00;      memory[33785] <=  8'h00;      memory[33786] <=  8'h00;      memory[33787] <=  8'h00;      memory[33788] <=  8'h00;      memory[33789] <=  8'h00;      memory[33790] <=  8'h00;      memory[33791] <=  8'h00;      memory[33792] <=  8'h00;      memory[33793] <=  8'h00;      memory[33794] <=  8'h00;      memory[33795] <=  8'h00;      memory[33796] <=  8'h00;      memory[33797] <=  8'h00;      memory[33798] <=  8'h00;      memory[33799] <=  8'h00;      memory[33800] <=  8'h00;      memory[33801] <=  8'h00;      memory[33802] <=  8'h00;      memory[33803] <=  8'h00;      memory[33804] <=  8'h00;      memory[33805] <=  8'h00;      memory[33806] <=  8'h00;      memory[33807] <=  8'h00;      memory[33808] <=  8'h00;      memory[33809] <=  8'h00;      memory[33810] <=  8'h00;      memory[33811] <=  8'h00;      memory[33812] <=  8'h00;      memory[33813] <=  8'h00;      memory[33814] <=  8'h00;      memory[33815] <=  8'h00;      memory[33816] <=  8'h00;      memory[33817] <=  8'h00;      memory[33818] <=  8'h00;      memory[33819] <=  8'h00;      memory[33820] <=  8'h00;      memory[33821] <=  8'h00;      memory[33822] <=  8'h00;      memory[33823] <=  8'h00;      memory[33824] <=  8'h00;      memory[33825] <=  8'h00;      memory[33826] <=  8'h00;      memory[33827] <=  8'h00;      memory[33828] <=  8'h00;      memory[33829] <=  8'h00;      memory[33830] <=  8'h00;      memory[33831] <=  8'h00;      memory[33832] <=  8'h00;      memory[33833] <=  8'h00;      memory[33834] <=  8'h00;      memory[33835] <=  8'h00;      memory[33836] <=  8'h00;      memory[33837] <=  8'h00;      memory[33838] <=  8'h00;      memory[33839] <=  8'h00;      memory[33840] <=  8'h00;      memory[33841] <=  8'h00;      memory[33842] <=  8'h00;      memory[33843] <=  8'h00;      memory[33844] <=  8'h00;      memory[33845] <=  8'h00;      memory[33846] <=  8'h00;      memory[33847] <=  8'h00;      memory[33848] <=  8'h00;      memory[33849] <=  8'h00;      memory[33850] <=  8'h00;      memory[33851] <=  8'h00;      memory[33852] <=  8'h00;      memory[33853] <=  8'h00;      memory[33854] <=  8'h00;      memory[33855] <=  8'h00;      memory[33856] <=  8'h00;      memory[33857] <=  8'h00;      memory[33858] <=  8'h00;      memory[33859] <=  8'h00;      memory[33860] <=  8'h00;      memory[33861] <=  8'h00;      memory[33862] <=  8'h00;      memory[33863] <=  8'h00;      memory[33864] <=  8'h00;      memory[33865] <=  8'h00;      memory[33866] <=  8'h00;      memory[33867] <=  8'h00;      memory[33868] <=  8'h00;      memory[33869] <=  8'h00;      memory[33870] <=  8'h00;      memory[33871] <=  8'h00;      memory[33872] <=  8'h00;      memory[33873] <=  8'h00;      memory[33874] <=  8'h00;      memory[33875] <=  8'h00;      memory[33876] <=  8'h00;      memory[33877] <=  8'h00;      memory[33878] <=  8'h00;      memory[33879] <=  8'h00;      memory[33880] <=  8'h00;      memory[33881] <=  8'h00;      memory[33882] <=  8'h00;      memory[33883] <=  8'h00;      memory[33884] <=  8'h00;      memory[33885] <=  8'h00;      memory[33886] <=  8'h00;      memory[33887] <=  8'h00;      memory[33888] <=  8'h00;      memory[33889] <=  8'h00;      memory[33890] <=  8'h00;      memory[33891] <=  8'h00;      memory[33892] <=  8'h00;      memory[33893] <=  8'h00;      memory[33894] <=  8'h00;      memory[33895] <=  8'h00;      memory[33896] <=  8'h00;      memory[33897] <=  8'h00;      memory[33898] <=  8'h00;      memory[33899] <=  8'h00;      memory[33900] <=  8'h00;      memory[33901] <=  8'h00;      memory[33902] <=  8'h00;      memory[33903] <=  8'h00;      memory[33904] <=  8'h00;      memory[33905] <=  8'h00;      memory[33906] <=  8'h00;      memory[33907] <=  8'h00;      memory[33908] <=  8'h00;      memory[33909] <=  8'h00;      memory[33910] <=  8'h00;      memory[33911] <=  8'h00;      memory[33912] <=  8'h00;      memory[33913] <=  8'h00;      memory[33914] <=  8'h00;      memory[33915] <=  8'h00;      memory[33916] <=  8'h00;      memory[33917] <=  8'h00;      memory[33918] <=  8'h00;      memory[33919] <=  8'h00;      memory[33920] <=  8'h00;      memory[33921] <=  8'h00;      memory[33922] <=  8'h00;      memory[33923] <=  8'h00;      memory[33924] <=  8'h00;      memory[33925] <=  8'h00;      memory[33926] <=  8'h00;      memory[33927] <=  8'h00;      memory[33928] <=  8'h00;      memory[33929] <=  8'h00;      memory[33930] <=  8'h00;      memory[33931] <=  8'h00;      memory[33932] <=  8'h00;      memory[33933] <=  8'h00;      memory[33934] <=  8'h00;      memory[33935] <=  8'h00;      memory[33936] <=  8'h00;      memory[33937] <=  8'h00;      memory[33938] <=  8'h00;      memory[33939] <=  8'h00;      memory[33940] <=  8'h00;      memory[33941] <=  8'h00;      memory[33942] <=  8'h00;      memory[33943] <=  8'h00;      memory[33944] <=  8'h00;      memory[33945] <=  8'h00;      memory[33946] <=  8'h00;      memory[33947] <=  8'h00;      memory[33948] <=  8'h00;      memory[33949] <=  8'h00;      memory[33950] <=  8'h00;      memory[33951] <=  8'h00;      memory[33952] <=  8'h00;      memory[33953] <=  8'h00;      memory[33954] <=  8'h00;      memory[33955] <=  8'h00;      memory[33956] <=  8'h00;      memory[33957] <=  8'h00;      memory[33958] <=  8'h00;      memory[33959] <=  8'h00;      memory[33960] <=  8'h00;      memory[33961] <=  8'h00;      memory[33962] <=  8'h00;      memory[33963] <=  8'h00;      memory[33964] <=  8'h00;      memory[33965] <=  8'h00;      memory[33966] <=  8'h00;      memory[33967] <=  8'h00;      memory[33968] <=  8'h00;      memory[33969] <=  8'h00;      memory[33970] <=  8'h00;      memory[33971] <=  8'h00;      memory[33972] <=  8'h00;      memory[33973] <=  8'h00;      memory[33974] <=  8'h00;      memory[33975] <=  8'h00;      memory[33976] <=  8'h00;      memory[33977] <=  8'h00;      memory[33978] <=  8'h00;      memory[33979] <=  8'h00;      memory[33980] <=  8'h00;      memory[33981] <=  8'h00;      memory[33982] <=  8'h00;      memory[33983] <=  8'h00;      memory[33984] <=  8'h00;      memory[33985] <=  8'h00;      memory[33986] <=  8'h00;      memory[33987] <=  8'h00;      memory[33988] <=  8'h00;      memory[33989] <=  8'h00;      memory[33990] <=  8'h00;      memory[33991] <=  8'h00;      memory[33992] <=  8'h00;      memory[33993] <=  8'h00;      memory[33994] <=  8'h00;      memory[33995] <=  8'h00;      memory[33996] <=  8'h00;      memory[33997] <=  8'h00;      memory[33998] <=  8'h00;      memory[33999] <=  8'h00;      memory[34000] <=  8'h00;      memory[34001] <=  8'h00;      memory[34002] <=  8'h00;      memory[34003] <=  8'h00;      memory[34004] <=  8'h00;      memory[34005] <=  8'h00;      memory[34006] <=  8'h00;      memory[34007] <=  8'h00;      memory[34008] <=  8'h00;      memory[34009] <=  8'h00;      memory[34010] <=  8'h00;      memory[34011] <=  8'h00;      memory[34012] <=  8'h00;      memory[34013] <=  8'h00;      memory[34014] <=  8'h00;      memory[34015] <=  8'h00;      memory[34016] <=  8'h00;      memory[34017] <=  8'h00;      memory[34018] <=  8'h00;      memory[34019] <=  8'h00;      memory[34020] <=  8'h00;      memory[34021] <=  8'h00;      memory[34022] <=  8'h00;      memory[34023] <=  8'h00;      memory[34024] <=  8'h00;      memory[34025] <=  8'h00;      memory[34026] <=  8'h00;      memory[34027] <=  8'h00;      memory[34028] <=  8'h00;      memory[34029] <=  8'h00;      memory[34030] <=  8'h00;      memory[34031] <=  8'h00;      memory[34032] <=  8'h00;      memory[34033] <=  8'h00;      memory[34034] <=  8'h00;      memory[34035] <=  8'h00;      memory[34036] <=  8'h00;      memory[34037] <=  8'h00;      memory[34038] <=  8'h00;      memory[34039] <=  8'h00;      memory[34040] <=  8'h00;      memory[34041] <=  8'h00;      memory[34042] <=  8'h00;      memory[34043] <=  8'h00;      memory[34044] <=  8'h00;      memory[34045] <=  8'h00;      memory[34046] <=  8'h00;      memory[34047] <=  8'h00;      memory[34048] <=  8'h00;      memory[34049] <=  8'h00;      memory[34050] <=  8'h00;      memory[34051] <=  8'h00;      memory[34052] <=  8'h00;      memory[34053] <=  8'h00;      memory[34054] <=  8'h00;      memory[34055] <=  8'h00;      memory[34056] <=  8'h00;      memory[34057] <=  8'h00;      memory[34058] <=  8'h00;      memory[34059] <=  8'h00;      memory[34060] <=  8'h00;      memory[34061] <=  8'h00;      memory[34062] <=  8'h00;      memory[34063] <=  8'h00;      memory[34064] <=  8'h00;      memory[34065] <=  8'h00;      memory[34066] <=  8'h00;      memory[34067] <=  8'h00;      memory[34068] <=  8'h00;      memory[34069] <=  8'h00;      memory[34070] <=  8'h00;      memory[34071] <=  8'h00;      memory[34072] <=  8'h00;      memory[34073] <=  8'h00;      memory[34074] <=  8'h00;      memory[34075] <=  8'h00;      memory[34076] <=  8'h00;      memory[34077] <=  8'h00;      memory[34078] <=  8'h00;      memory[34079] <=  8'h00;      memory[34080] <=  8'h00;      memory[34081] <=  8'h00;      memory[34082] <=  8'h00;      memory[34083] <=  8'h00;      memory[34084] <=  8'h00;      memory[34085] <=  8'h00;      memory[34086] <=  8'h00;      memory[34087] <=  8'h00;      memory[34088] <=  8'h00;      memory[34089] <=  8'h00;      memory[34090] <=  8'h00;      memory[34091] <=  8'h00;      memory[34092] <=  8'h00;      memory[34093] <=  8'h00;      memory[34094] <=  8'h00;      memory[34095] <=  8'h00;      memory[34096] <=  8'h00;      memory[34097] <=  8'h00;      memory[34098] <=  8'h00;      memory[34099] <=  8'h00;      memory[34100] <=  8'h00;      memory[34101] <=  8'h00;      memory[34102] <=  8'h00;      memory[34103] <=  8'h00;      memory[34104] <=  8'h00;      memory[34105] <=  8'h00;      memory[34106] <=  8'h00;      memory[34107] <=  8'h00;      memory[34108] <=  8'h00;      memory[34109] <=  8'h00;      memory[34110] <=  8'h00;      memory[34111] <=  8'h00;      memory[34112] <=  8'h00;      memory[34113] <=  8'h00;      memory[34114] <=  8'h00;      memory[34115] <=  8'h00;      memory[34116] <=  8'h00;      memory[34117] <=  8'h00;      memory[34118] <=  8'h00;      memory[34119] <=  8'h00;      memory[34120] <=  8'h00;      memory[34121] <=  8'h00;      memory[34122] <=  8'h00;      memory[34123] <=  8'h00;      memory[34124] <=  8'h00;      memory[34125] <=  8'h00;      memory[34126] <=  8'h00;      memory[34127] <=  8'h00;      memory[34128] <=  8'h00;      memory[34129] <=  8'h00;      memory[34130] <=  8'h00;      memory[34131] <=  8'h00;      memory[34132] <=  8'h00;      memory[34133] <=  8'h00;      memory[34134] <=  8'h00;      memory[34135] <=  8'h00;      memory[34136] <=  8'h00;      memory[34137] <=  8'h00;      memory[34138] <=  8'h00;      memory[34139] <=  8'h00;      memory[34140] <=  8'h00;      memory[34141] <=  8'h00;      memory[34142] <=  8'h00;      memory[34143] <=  8'h00;      memory[34144] <=  8'h00;      memory[34145] <=  8'h00;      memory[34146] <=  8'h00;      memory[34147] <=  8'h00;      memory[34148] <=  8'h00;      memory[34149] <=  8'h00;      memory[34150] <=  8'h00;      memory[34151] <=  8'h00;      memory[34152] <=  8'h00;      memory[34153] <=  8'h00;      memory[34154] <=  8'h00;      memory[34155] <=  8'h00;      memory[34156] <=  8'h00;      memory[34157] <=  8'h00;      memory[34158] <=  8'h00;      memory[34159] <=  8'h00;      memory[34160] <=  8'h00;      memory[34161] <=  8'h00;      memory[34162] <=  8'h00;      memory[34163] <=  8'h00;      memory[34164] <=  8'h00;      memory[34165] <=  8'h00;      memory[34166] <=  8'h00;      memory[34167] <=  8'h00;      memory[34168] <=  8'h00;      memory[34169] <=  8'h00;      memory[34170] <=  8'h00;      memory[34171] <=  8'h00;      memory[34172] <=  8'h00;      memory[34173] <=  8'h00;      memory[34174] <=  8'h00;      memory[34175] <=  8'h00;      memory[34176] <=  8'h00;      memory[34177] <=  8'h00;      memory[34178] <=  8'h00;      memory[34179] <=  8'h00;      memory[34180] <=  8'h00;      memory[34181] <=  8'h00;      memory[34182] <=  8'h00;      memory[34183] <=  8'h00;      memory[34184] <=  8'h00;      memory[34185] <=  8'h00;      memory[34186] <=  8'h00;      memory[34187] <=  8'h00;      memory[34188] <=  8'h00;      memory[34189] <=  8'h00;      memory[34190] <=  8'h00;      memory[34191] <=  8'h00;      memory[34192] <=  8'h00;      memory[34193] <=  8'h00;      memory[34194] <=  8'h00;      memory[34195] <=  8'h00;      memory[34196] <=  8'h00;      memory[34197] <=  8'h00;      memory[34198] <=  8'h00;      memory[34199] <=  8'h00;      memory[34200] <=  8'h00;      memory[34201] <=  8'h00;      memory[34202] <=  8'h00;      memory[34203] <=  8'h00;      memory[34204] <=  8'h00;      memory[34205] <=  8'h00;      memory[34206] <=  8'h00;      memory[34207] <=  8'h00;      memory[34208] <=  8'h00;      memory[34209] <=  8'h00;      memory[34210] <=  8'h00;      memory[34211] <=  8'h00;      memory[34212] <=  8'h00;      memory[34213] <=  8'h00;      memory[34214] <=  8'h00;      memory[34215] <=  8'h00;      memory[34216] <=  8'h00;      memory[34217] <=  8'h00;      memory[34218] <=  8'h00;      memory[34219] <=  8'h00;      memory[34220] <=  8'h00;      memory[34221] <=  8'h00;      memory[34222] <=  8'h00;      memory[34223] <=  8'h00;      memory[34224] <=  8'h00;      memory[34225] <=  8'h00;      memory[34226] <=  8'h00;      memory[34227] <=  8'h00;      memory[34228] <=  8'h00;      memory[34229] <=  8'h00;      memory[34230] <=  8'h00;      memory[34231] <=  8'h00;      memory[34232] <=  8'h00;      memory[34233] <=  8'h00;      memory[34234] <=  8'h00;      memory[34235] <=  8'h00;      memory[34236] <=  8'h00;      memory[34237] <=  8'h00;      memory[34238] <=  8'h00;      memory[34239] <=  8'h00;      memory[34240] <=  8'h00;      memory[34241] <=  8'h00;      memory[34242] <=  8'h00;      memory[34243] <=  8'h00;      memory[34244] <=  8'h00;      memory[34245] <=  8'h00;      memory[34246] <=  8'h00;      memory[34247] <=  8'h00;      memory[34248] <=  8'h00;      memory[34249] <=  8'h00;      memory[34250] <=  8'h00;      memory[34251] <=  8'h00;      memory[34252] <=  8'h00;      memory[34253] <=  8'h00;      memory[34254] <=  8'h00;      memory[34255] <=  8'h00;      memory[34256] <=  8'h00;      memory[34257] <=  8'h00;      memory[34258] <=  8'h00;      memory[34259] <=  8'h00;      memory[34260] <=  8'h00;      memory[34261] <=  8'h00;      memory[34262] <=  8'h00;      memory[34263] <=  8'h00;      memory[34264] <=  8'h00;      memory[34265] <=  8'h00;      memory[34266] <=  8'h00;      memory[34267] <=  8'h00;      memory[34268] <=  8'h00;      memory[34269] <=  8'h00;      memory[34270] <=  8'h00;      memory[34271] <=  8'h00;      memory[34272] <=  8'h00;      memory[34273] <=  8'h00;      memory[34274] <=  8'h00;      memory[34275] <=  8'h00;      memory[34276] <=  8'h00;      memory[34277] <=  8'h00;      memory[34278] <=  8'h00;      memory[34279] <=  8'h00;      memory[34280] <=  8'h00;      memory[34281] <=  8'h00;      memory[34282] <=  8'h00;      memory[34283] <=  8'h00;      memory[34284] <=  8'h00;      memory[34285] <=  8'h00;      memory[34286] <=  8'h00;      memory[34287] <=  8'h00;      memory[34288] <=  8'h00;      memory[34289] <=  8'h00;      memory[34290] <=  8'h00;      memory[34291] <=  8'h00;      memory[34292] <=  8'h00;      memory[34293] <=  8'h00;      memory[34294] <=  8'h00;      memory[34295] <=  8'h00;      memory[34296] <=  8'h00;      memory[34297] <=  8'h00;      memory[34298] <=  8'h00;      memory[34299] <=  8'h00;      memory[34300] <=  8'h00;      memory[34301] <=  8'h00;      memory[34302] <=  8'h00;      memory[34303] <=  8'h00;      memory[34304] <=  8'h00;      memory[34305] <=  8'h00;      memory[34306] <=  8'h00;      memory[34307] <=  8'h00;      memory[34308] <=  8'h00;      memory[34309] <=  8'h00;      memory[34310] <=  8'h00;      memory[34311] <=  8'h00;      memory[34312] <=  8'h00;      memory[34313] <=  8'h00;      memory[34314] <=  8'h00;      memory[34315] <=  8'h00;      memory[34316] <=  8'h00;      memory[34317] <=  8'h00;      memory[34318] <=  8'h00;      memory[34319] <=  8'h00;      memory[34320] <=  8'h00;      memory[34321] <=  8'h00;      memory[34322] <=  8'h00;      memory[34323] <=  8'h00;      memory[34324] <=  8'h00;      memory[34325] <=  8'h00;      memory[34326] <=  8'h00;      memory[34327] <=  8'h00;      memory[34328] <=  8'h00;      memory[34329] <=  8'h00;      memory[34330] <=  8'h00;      memory[34331] <=  8'h00;      memory[34332] <=  8'h00;      memory[34333] <=  8'h00;      memory[34334] <=  8'h00;      memory[34335] <=  8'h00;      memory[34336] <=  8'h00;      memory[34337] <=  8'h00;      memory[34338] <=  8'h00;      memory[34339] <=  8'h00;      memory[34340] <=  8'h00;      memory[34341] <=  8'h00;      memory[34342] <=  8'h00;      memory[34343] <=  8'h00;      memory[34344] <=  8'h00;      memory[34345] <=  8'h00;      memory[34346] <=  8'h00;      memory[34347] <=  8'h00;      memory[34348] <=  8'h00;      memory[34349] <=  8'h00;      memory[34350] <=  8'h00;      memory[34351] <=  8'h00;      memory[34352] <=  8'h00;      memory[34353] <=  8'h00;      memory[34354] <=  8'h00;      memory[34355] <=  8'h00;      memory[34356] <=  8'h00;      memory[34357] <=  8'h00;      memory[34358] <=  8'h00;      memory[34359] <=  8'h00;      memory[34360] <=  8'h00;      memory[34361] <=  8'h00;      memory[34362] <=  8'h00;      memory[34363] <=  8'h00;      memory[34364] <=  8'h00;      memory[34365] <=  8'h00;      memory[34366] <=  8'h00;      memory[34367] <=  8'h00;      memory[34368] <=  8'h00;      memory[34369] <=  8'h00;      memory[34370] <=  8'h00;      memory[34371] <=  8'h00;      memory[34372] <=  8'h00;      memory[34373] <=  8'h00;      memory[34374] <=  8'h00;      memory[34375] <=  8'h00;      memory[34376] <=  8'h00;      memory[34377] <=  8'h00;      memory[34378] <=  8'h00;      memory[34379] <=  8'h00;      memory[34380] <=  8'h00;      memory[34381] <=  8'h00;      memory[34382] <=  8'h00;      memory[34383] <=  8'h00;      memory[34384] <=  8'h00;      memory[34385] <=  8'h00;      memory[34386] <=  8'h00;      memory[34387] <=  8'h00;      memory[34388] <=  8'h00;      memory[34389] <=  8'h00;      memory[34390] <=  8'h00;      memory[34391] <=  8'h00;      memory[34392] <=  8'h00;      memory[34393] <=  8'h00;      memory[34394] <=  8'h00;      memory[34395] <=  8'h00;      memory[34396] <=  8'h00;      memory[34397] <=  8'h00;      memory[34398] <=  8'h00;      memory[34399] <=  8'h00;      memory[34400] <=  8'h00;      memory[34401] <=  8'h00;      memory[34402] <=  8'h00;      memory[34403] <=  8'h00;      memory[34404] <=  8'h00;      memory[34405] <=  8'h00;      memory[34406] <=  8'h00;      memory[34407] <=  8'h00;      memory[34408] <=  8'h00;      memory[34409] <=  8'h00;      memory[34410] <=  8'h00;      memory[34411] <=  8'h00;      memory[34412] <=  8'h00;      memory[34413] <=  8'h00;      memory[34414] <=  8'h00;      memory[34415] <=  8'h00;      memory[34416] <=  8'h00;      memory[34417] <=  8'h00;      memory[34418] <=  8'h00;      memory[34419] <=  8'h00;      memory[34420] <=  8'h00;      memory[34421] <=  8'h00;      memory[34422] <=  8'h00;      memory[34423] <=  8'h00;      memory[34424] <=  8'h00;      memory[34425] <=  8'h00;      memory[34426] <=  8'h00;      memory[34427] <=  8'h00;      memory[34428] <=  8'h00;      memory[34429] <=  8'h00;      memory[34430] <=  8'h00;      memory[34431] <=  8'h00;      memory[34432] <=  8'h00;      memory[34433] <=  8'h00;      memory[34434] <=  8'h00;      memory[34435] <=  8'h00;      memory[34436] <=  8'h00;      memory[34437] <=  8'h00;      memory[34438] <=  8'h00;      memory[34439] <=  8'h00;      memory[34440] <=  8'h00;      memory[34441] <=  8'h00;      memory[34442] <=  8'h00;      memory[34443] <=  8'h00;      memory[34444] <=  8'h00;      memory[34445] <=  8'h00;      memory[34446] <=  8'h00;      memory[34447] <=  8'h00;      memory[34448] <=  8'h00;      memory[34449] <=  8'h00;      memory[34450] <=  8'h00;      memory[34451] <=  8'h00;      memory[34452] <=  8'h00;      memory[34453] <=  8'h00;      memory[34454] <=  8'h00;      memory[34455] <=  8'h00;      memory[34456] <=  8'h00;      memory[34457] <=  8'h00;      memory[34458] <=  8'h00;      memory[34459] <=  8'h00;      memory[34460] <=  8'h00;      memory[34461] <=  8'h00;      memory[34462] <=  8'h00;      memory[34463] <=  8'h00;      memory[34464] <=  8'h00;      memory[34465] <=  8'h00;      memory[34466] <=  8'h00;      memory[34467] <=  8'h00;      memory[34468] <=  8'h00;      memory[34469] <=  8'h00;      memory[34470] <=  8'h00;      memory[34471] <=  8'h00;      memory[34472] <=  8'h00;      memory[34473] <=  8'h00;      memory[34474] <=  8'h00;      memory[34475] <=  8'h00;      memory[34476] <=  8'h00;      memory[34477] <=  8'h00;      memory[34478] <=  8'h00;      memory[34479] <=  8'h00;      memory[34480] <=  8'h00;      memory[34481] <=  8'h00;      memory[34482] <=  8'h00;      memory[34483] <=  8'h00;      memory[34484] <=  8'h00;      memory[34485] <=  8'h00;      memory[34486] <=  8'h00;      memory[34487] <=  8'h00;      memory[34488] <=  8'h00;      memory[34489] <=  8'h00;      memory[34490] <=  8'h00;      memory[34491] <=  8'h00;      memory[34492] <=  8'h00;      memory[34493] <=  8'h00;      memory[34494] <=  8'h00;      memory[34495] <=  8'h00;      memory[34496] <=  8'h00;      memory[34497] <=  8'h00;      memory[34498] <=  8'h00;      memory[34499] <=  8'h00;      memory[34500] <=  8'h00;      memory[34501] <=  8'h00;      memory[34502] <=  8'h00;      memory[34503] <=  8'h00;      memory[34504] <=  8'h00;      memory[34505] <=  8'h00;      memory[34506] <=  8'h00;      memory[34507] <=  8'h00;      memory[34508] <=  8'h00;      memory[34509] <=  8'h00;      memory[34510] <=  8'h00;      memory[34511] <=  8'h00;      memory[34512] <=  8'h00;      memory[34513] <=  8'h00;      memory[34514] <=  8'h00;      memory[34515] <=  8'h00;      memory[34516] <=  8'h00;      memory[34517] <=  8'h00;      memory[34518] <=  8'h00;      memory[34519] <=  8'h00;      memory[34520] <=  8'h00;      memory[34521] <=  8'h00;      memory[34522] <=  8'h00;      memory[34523] <=  8'h00;      memory[34524] <=  8'h00;      memory[34525] <=  8'h00;      memory[34526] <=  8'h00;      memory[34527] <=  8'h00;      memory[34528] <=  8'h00;      memory[34529] <=  8'h00;      memory[34530] <=  8'h00;      memory[34531] <=  8'h00;      memory[34532] <=  8'h00;      memory[34533] <=  8'h00;      memory[34534] <=  8'h00;      memory[34535] <=  8'h00;      memory[34536] <=  8'h00;      memory[34537] <=  8'h00;      memory[34538] <=  8'h00;      memory[34539] <=  8'h00;      memory[34540] <=  8'h00;      memory[34541] <=  8'h00;      memory[34542] <=  8'h00;      memory[34543] <=  8'h00;      memory[34544] <=  8'h00;      memory[34545] <=  8'h00;      memory[34546] <=  8'h00;      memory[34547] <=  8'h00;      memory[34548] <=  8'h00;      memory[34549] <=  8'h00;      memory[34550] <=  8'h00;      memory[34551] <=  8'h00;      memory[34552] <=  8'h00;      memory[34553] <=  8'h00;      memory[34554] <=  8'h00;      memory[34555] <=  8'h00;      memory[34556] <=  8'h00;      memory[34557] <=  8'h00;      memory[34558] <=  8'h00;      memory[34559] <=  8'h00;      memory[34560] <=  8'h00;      memory[34561] <=  8'h00;      memory[34562] <=  8'h00;      memory[34563] <=  8'h00;      memory[34564] <=  8'h00;      memory[34565] <=  8'h00;      memory[34566] <=  8'h00;      memory[34567] <=  8'h00;      memory[34568] <=  8'h00;      memory[34569] <=  8'h00;      memory[34570] <=  8'h00;      memory[34571] <=  8'h00;      memory[34572] <=  8'h00;      memory[34573] <=  8'h00;      memory[34574] <=  8'h00;      memory[34575] <=  8'h00;      memory[34576] <=  8'h00;      memory[34577] <=  8'h00;      memory[34578] <=  8'h00;      memory[34579] <=  8'h00;      memory[34580] <=  8'h00;      memory[34581] <=  8'h00;      memory[34582] <=  8'h00;      memory[34583] <=  8'h00;      memory[34584] <=  8'h00;      memory[34585] <=  8'h00;      memory[34586] <=  8'h00;      memory[34587] <=  8'h00;      memory[34588] <=  8'h00;      memory[34589] <=  8'h00;      memory[34590] <=  8'h00;      memory[34591] <=  8'h00;      memory[34592] <=  8'h00;      memory[34593] <=  8'h00;      memory[34594] <=  8'h00;      memory[34595] <=  8'h00;      memory[34596] <=  8'h00;      memory[34597] <=  8'h00;      memory[34598] <=  8'h00;      memory[34599] <=  8'h00;      memory[34600] <=  8'h00;      memory[34601] <=  8'h00;      memory[34602] <=  8'h00;      memory[34603] <=  8'h00;      memory[34604] <=  8'h00;      memory[34605] <=  8'h00;      memory[34606] <=  8'h00;      memory[34607] <=  8'h00;      memory[34608] <=  8'h00;      memory[34609] <=  8'h00;      memory[34610] <=  8'h00;      memory[34611] <=  8'h00;      memory[34612] <=  8'h00;      memory[34613] <=  8'h00;      memory[34614] <=  8'h00;      memory[34615] <=  8'h00;      memory[34616] <=  8'h00;      memory[34617] <=  8'h00;      memory[34618] <=  8'h00;      memory[34619] <=  8'h00;      memory[34620] <=  8'h00;      memory[34621] <=  8'h00;      memory[34622] <=  8'h00;      memory[34623] <=  8'h00;      memory[34624] <=  8'h00;      memory[34625] <=  8'h00;      memory[34626] <=  8'h00;      memory[34627] <=  8'h00;      memory[34628] <=  8'h00;      memory[34629] <=  8'h00;      memory[34630] <=  8'h00;      memory[34631] <=  8'h00;      memory[34632] <=  8'h00;      memory[34633] <=  8'h00;      memory[34634] <=  8'h00;      memory[34635] <=  8'h00;      memory[34636] <=  8'h00;      memory[34637] <=  8'h00;      memory[34638] <=  8'h00;      memory[34639] <=  8'h00;      memory[34640] <=  8'h00;      memory[34641] <=  8'h00;      memory[34642] <=  8'h00;      memory[34643] <=  8'h00;      memory[34644] <=  8'h00;      memory[34645] <=  8'h00;      memory[34646] <=  8'h00;      memory[34647] <=  8'h00;      memory[34648] <=  8'h00;      memory[34649] <=  8'h00;      memory[34650] <=  8'h00;      memory[34651] <=  8'h00;      memory[34652] <=  8'h00;      memory[34653] <=  8'h00;      memory[34654] <=  8'h00;      memory[34655] <=  8'h00;      memory[34656] <=  8'h00;      memory[34657] <=  8'h00;      memory[34658] <=  8'h00;      memory[34659] <=  8'h00;      memory[34660] <=  8'h00;      memory[34661] <=  8'h00;      memory[34662] <=  8'h00;      memory[34663] <=  8'h00;      memory[34664] <=  8'h00;      memory[34665] <=  8'h00;      memory[34666] <=  8'h00;      memory[34667] <=  8'h00;      memory[34668] <=  8'h00;      memory[34669] <=  8'h00;      memory[34670] <=  8'h00;      memory[34671] <=  8'h00;      memory[34672] <=  8'h00;      memory[34673] <=  8'h00;      memory[34674] <=  8'h00;      memory[34675] <=  8'h00;      memory[34676] <=  8'h00;      memory[34677] <=  8'h00;      memory[34678] <=  8'h00;      memory[34679] <=  8'h00;      memory[34680] <=  8'h00;      memory[34681] <=  8'h00;      memory[34682] <=  8'h00;      memory[34683] <=  8'h00;      memory[34684] <=  8'h00;      memory[34685] <=  8'h00;      memory[34686] <=  8'h00;      memory[34687] <=  8'h00;      memory[34688] <=  8'h00;      memory[34689] <=  8'h00;      memory[34690] <=  8'h00;      memory[34691] <=  8'h00;      memory[34692] <=  8'h00;      memory[34693] <=  8'h00;      memory[34694] <=  8'h00;      memory[34695] <=  8'h00;      memory[34696] <=  8'h00;      memory[34697] <=  8'h00;      memory[34698] <=  8'h00;      memory[34699] <=  8'h00;      memory[34700] <=  8'h00;      memory[34701] <=  8'h00;      memory[34702] <=  8'h00;      memory[34703] <=  8'h00;      memory[34704] <=  8'h00;      memory[34705] <=  8'h00;      memory[34706] <=  8'h00;      memory[34707] <=  8'h00;      memory[34708] <=  8'h00;      memory[34709] <=  8'h00;      memory[34710] <=  8'h00;      memory[34711] <=  8'h00;      memory[34712] <=  8'h00;      memory[34713] <=  8'h00;      memory[34714] <=  8'h00;      memory[34715] <=  8'h00;      memory[34716] <=  8'h00;      memory[34717] <=  8'h00;      memory[34718] <=  8'h00;      memory[34719] <=  8'h00;      memory[34720] <=  8'h00;      memory[34721] <=  8'h00;      memory[34722] <=  8'h00;      memory[34723] <=  8'h00;      memory[34724] <=  8'h00;      memory[34725] <=  8'h00;      memory[34726] <=  8'h00;      memory[34727] <=  8'h00;      memory[34728] <=  8'h00;      memory[34729] <=  8'h00;      memory[34730] <=  8'h00;      memory[34731] <=  8'h00;      memory[34732] <=  8'h00;      memory[34733] <=  8'h00;      memory[34734] <=  8'h00;      memory[34735] <=  8'h00;      memory[34736] <=  8'h00;      memory[34737] <=  8'h00;      memory[34738] <=  8'h00;      memory[34739] <=  8'h00;      memory[34740] <=  8'h00;      memory[34741] <=  8'h00;      memory[34742] <=  8'h00;      memory[34743] <=  8'h00;      memory[34744] <=  8'h00;      memory[34745] <=  8'h00;      memory[34746] <=  8'h00;      memory[34747] <=  8'h00;      memory[34748] <=  8'h00;      memory[34749] <=  8'h00;      memory[34750] <=  8'h00;      memory[34751] <=  8'h00;      memory[34752] <=  8'h00;      memory[34753] <=  8'h00;      memory[34754] <=  8'h00;      memory[34755] <=  8'h00;      memory[34756] <=  8'h00;      memory[34757] <=  8'h00;      memory[34758] <=  8'h00;      memory[34759] <=  8'h00;      memory[34760] <=  8'h00;      memory[34761] <=  8'h00;      memory[34762] <=  8'h00;      memory[34763] <=  8'h00;      memory[34764] <=  8'h00;      memory[34765] <=  8'h00;      memory[34766] <=  8'h00;      memory[34767] <=  8'h00;      memory[34768] <=  8'h00;      memory[34769] <=  8'h00;      memory[34770] <=  8'h00;      memory[34771] <=  8'h00;      memory[34772] <=  8'h00;      memory[34773] <=  8'h00;      memory[34774] <=  8'h00;      memory[34775] <=  8'h00;      memory[34776] <=  8'h00;      memory[34777] <=  8'h00;      memory[34778] <=  8'h00;      memory[34779] <=  8'h00;      memory[34780] <=  8'h00;      memory[34781] <=  8'h00;      memory[34782] <=  8'h00;      memory[34783] <=  8'h00;      memory[34784] <=  8'h00;      memory[34785] <=  8'h00;      memory[34786] <=  8'h00;      memory[34787] <=  8'h00;      memory[34788] <=  8'h00;      memory[34789] <=  8'h00;      memory[34790] <=  8'h00;      memory[34791] <=  8'h00;      memory[34792] <=  8'h00;      memory[34793] <=  8'h00;      memory[34794] <=  8'h00;      memory[34795] <=  8'h00;      memory[34796] <=  8'h00;      memory[34797] <=  8'h00;      memory[34798] <=  8'h00;      memory[34799] <=  8'h00;      memory[34800] <=  8'h00;      memory[34801] <=  8'h00;      memory[34802] <=  8'h00;      memory[34803] <=  8'h00;      memory[34804] <=  8'h00;      memory[34805] <=  8'h00;      memory[34806] <=  8'h00;      memory[34807] <=  8'h00;      memory[34808] <=  8'h00;      memory[34809] <=  8'h00;      memory[34810] <=  8'h00;      memory[34811] <=  8'h00;      memory[34812] <=  8'h00;      memory[34813] <=  8'h00;      memory[34814] <=  8'h00;      memory[34815] <=  8'h00;      memory[34816] <=  8'h00;      memory[34817] <=  8'h00;      memory[34818] <=  8'h00;      memory[34819] <=  8'h00;      memory[34820] <=  8'h00;      memory[34821] <=  8'h00;      memory[34822] <=  8'h00;      memory[34823] <=  8'h00;      memory[34824] <=  8'h00;      memory[34825] <=  8'h00;      memory[34826] <=  8'h00;      memory[34827] <=  8'h00;      memory[34828] <=  8'h00;      memory[34829] <=  8'h00;      memory[34830] <=  8'h00;      memory[34831] <=  8'h00;      memory[34832] <=  8'h00;      memory[34833] <=  8'h00;      memory[34834] <=  8'h00;      memory[34835] <=  8'h00;      memory[34836] <=  8'h00;      memory[34837] <=  8'h00;      memory[34838] <=  8'h00;      memory[34839] <=  8'h00;      memory[34840] <=  8'h00;      memory[34841] <=  8'h00;      memory[34842] <=  8'h00;      memory[34843] <=  8'h00;      memory[34844] <=  8'h00;      memory[34845] <=  8'h00;      memory[34846] <=  8'h00;      memory[34847] <=  8'h00;      memory[34848] <=  8'h00;      memory[34849] <=  8'h00;      memory[34850] <=  8'h00;      memory[34851] <=  8'h00;      memory[34852] <=  8'h00;      memory[34853] <=  8'h00;      memory[34854] <=  8'h00;      memory[34855] <=  8'h00;      memory[34856] <=  8'h00;      memory[34857] <=  8'h00;      memory[34858] <=  8'h00;      memory[34859] <=  8'h00;      memory[34860] <=  8'h00;      memory[34861] <=  8'h00;      memory[34862] <=  8'h00;      memory[34863] <=  8'h00;      memory[34864] <=  8'h00;      memory[34865] <=  8'h00;      memory[34866] <=  8'h00;      memory[34867] <=  8'h00;      memory[34868] <=  8'h00;      memory[34869] <=  8'h00;      memory[34870] <=  8'h00;      memory[34871] <=  8'h00;      memory[34872] <=  8'h00;      memory[34873] <=  8'h00;      memory[34874] <=  8'h00;      memory[34875] <=  8'h00;      memory[34876] <=  8'h00;      memory[34877] <=  8'h00;      memory[34878] <=  8'h00;      memory[34879] <=  8'h00;      memory[34880] <=  8'h00;      memory[34881] <=  8'h00;      memory[34882] <=  8'h00;      memory[34883] <=  8'h00;      memory[34884] <=  8'h00;      memory[34885] <=  8'h00;      memory[34886] <=  8'h00;      memory[34887] <=  8'h00;      memory[34888] <=  8'h00;      memory[34889] <=  8'h00;      memory[34890] <=  8'h00;      memory[34891] <=  8'h00;      memory[34892] <=  8'h00;      memory[34893] <=  8'h00;      memory[34894] <=  8'h00;      memory[34895] <=  8'h00;      memory[34896] <=  8'h00;      memory[34897] <=  8'h00;      memory[34898] <=  8'h00;      memory[34899] <=  8'h00;      memory[34900] <=  8'h00;      memory[34901] <=  8'h00;      memory[34902] <=  8'h00;      memory[34903] <=  8'h00;      memory[34904] <=  8'h00;      memory[34905] <=  8'h00;      memory[34906] <=  8'h00;      memory[34907] <=  8'h00;      memory[34908] <=  8'h00;      memory[34909] <=  8'h00;      memory[34910] <=  8'h00;      memory[34911] <=  8'h00;      memory[34912] <=  8'h00;      memory[34913] <=  8'h00;      memory[34914] <=  8'h00;      memory[34915] <=  8'h00;      memory[34916] <=  8'h00;      memory[34917] <=  8'h00;      memory[34918] <=  8'h00;      memory[34919] <=  8'h00;      memory[34920] <=  8'h00;      memory[34921] <=  8'h00;      memory[34922] <=  8'h00;      memory[34923] <=  8'h00;      memory[34924] <=  8'h00;      memory[34925] <=  8'h00;      memory[34926] <=  8'h00;      memory[34927] <=  8'h00;      memory[34928] <=  8'h00;      memory[34929] <=  8'h00;      memory[34930] <=  8'h00;      memory[34931] <=  8'h00;      memory[34932] <=  8'h00;      memory[34933] <=  8'h00;      memory[34934] <=  8'h00;      memory[34935] <=  8'h00;      memory[34936] <=  8'h00;      memory[34937] <=  8'h00;      memory[34938] <=  8'h00;      memory[34939] <=  8'h00;      memory[34940] <=  8'h00;      memory[34941] <=  8'h00;      memory[34942] <=  8'h00;      memory[34943] <=  8'h00;      memory[34944] <=  8'h00;      memory[34945] <=  8'h00;      memory[34946] <=  8'h00;      memory[34947] <=  8'h00;      memory[34948] <=  8'h00;      memory[34949] <=  8'h00;      memory[34950] <=  8'h00;      memory[34951] <=  8'h00;      memory[34952] <=  8'h00;      memory[34953] <=  8'h00;      memory[34954] <=  8'h00;      memory[34955] <=  8'h00;      memory[34956] <=  8'h00;      memory[34957] <=  8'h00;      memory[34958] <=  8'h00;      memory[34959] <=  8'h00;      memory[34960] <=  8'h00;      memory[34961] <=  8'h00;      memory[34962] <=  8'h00;      memory[34963] <=  8'h00;      memory[34964] <=  8'h00;      memory[34965] <=  8'h00;      memory[34966] <=  8'h00;      memory[34967] <=  8'h00;      memory[34968] <=  8'h00;      memory[34969] <=  8'h00;      memory[34970] <=  8'h00;      memory[34971] <=  8'h00;      memory[34972] <=  8'h00;      memory[34973] <=  8'h00;      memory[34974] <=  8'h00;      memory[34975] <=  8'h00;      memory[34976] <=  8'h00;      memory[34977] <=  8'h00;      memory[34978] <=  8'h00;      memory[34979] <=  8'h00;      memory[34980] <=  8'h00;      memory[34981] <=  8'h00;      memory[34982] <=  8'h00;      memory[34983] <=  8'h00;      memory[34984] <=  8'h00;      memory[34985] <=  8'h00;      memory[34986] <=  8'h00;      memory[34987] <=  8'h00;      memory[34988] <=  8'h00;      memory[34989] <=  8'h00;      memory[34990] <=  8'h00;      memory[34991] <=  8'h00;      memory[34992] <=  8'h00;      memory[34993] <=  8'h00;      memory[34994] <=  8'h00;      memory[34995] <=  8'h00;      memory[34996] <=  8'h00;      memory[34997] <=  8'h00;      memory[34998] <=  8'h00;      memory[34999] <=  8'h00;      memory[35000] <=  8'h00;      memory[35001] <=  8'h00;      memory[35002] <=  8'h00;      memory[35003] <=  8'h00;      memory[35004] <=  8'h00;      memory[35005] <=  8'h00;      memory[35006] <=  8'h00;      memory[35007] <=  8'h00;      memory[35008] <=  8'h00;      memory[35009] <=  8'h00;      memory[35010] <=  8'h00;      memory[35011] <=  8'h00;      memory[35012] <=  8'h00;      memory[35013] <=  8'h00;      memory[35014] <=  8'h00;      memory[35015] <=  8'h00;      memory[35016] <=  8'h00;      memory[35017] <=  8'h00;      memory[35018] <=  8'h00;      memory[35019] <=  8'h00;      memory[35020] <=  8'h00;      memory[35021] <=  8'h00;      memory[35022] <=  8'h00;      memory[35023] <=  8'h00;      memory[35024] <=  8'h00;      memory[35025] <=  8'h00;      memory[35026] <=  8'h00;      memory[35027] <=  8'h00;      memory[35028] <=  8'h00;      memory[35029] <=  8'h00;      memory[35030] <=  8'h00;      memory[35031] <=  8'h00;      memory[35032] <=  8'h00;      memory[35033] <=  8'h00;      memory[35034] <=  8'h00;      memory[35035] <=  8'h00;      memory[35036] <=  8'h00;      memory[35037] <=  8'h00;      memory[35038] <=  8'h00;      memory[35039] <=  8'h00;      memory[35040] <=  8'h00;      memory[35041] <=  8'h00;      memory[35042] <=  8'h00;      memory[35043] <=  8'h00;      memory[35044] <=  8'h00;      memory[35045] <=  8'h00;      memory[35046] <=  8'h00;      memory[35047] <=  8'h00;      memory[35048] <=  8'h00;      memory[35049] <=  8'h00;      memory[35050] <=  8'h00;      memory[35051] <=  8'h00;      memory[35052] <=  8'h00;      memory[35053] <=  8'h00;      memory[35054] <=  8'h00;      memory[35055] <=  8'h00;      memory[35056] <=  8'h00;      memory[35057] <=  8'h00;      memory[35058] <=  8'h00;      memory[35059] <=  8'h00;      memory[35060] <=  8'h00;      memory[35061] <=  8'h00;      memory[35062] <=  8'h00;      memory[35063] <=  8'h00;      memory[35064] <=  8'h00;      memory[35065] <=  8'h00;      memory[35066] <=  8'h00;      memory[35067] <=  8'h00;      memory[35068] <=  8'h00;      memory[35069] <=  8'h00;      memory[35070] <=  8'h00;      memory[35071] <=  8'h00;      memory[35072] <=  8'h00;      memory[35073] <=  8'h00;      memory[35074] <=  8'h00;      memory[35075] <=  8'h00;      memory[35076] <=  8'h00;      memory[35077] <=  8'h00;      memory[35078] <=  8'h00;      memory[35079] <=  8'h00;      memory[35080] <=  8'h00;      memory[35081] <=  8'h00;      memory[35082] <=  8'h00;      memory[35083] <=  8'h00;      memory[35084] <=  8'h00;      memory[35085] <=  8'h00;      memory[35086] <=  8'h00;      memory[35087] <=  8'h00;      memory[35088] <=  8'h00;      memory[35089] <=  8'h00;      memory[35090] <=  8'h00;      memory[35091] <=  8'h00;      memory[35092] <=  8'h00;      memory[35093] <=  8'h00;      memory[35094] <=  8'h00;      memory[35095] <=  8'h00;      memory[35096] <=  8'h00;      memory[35097] <=  8'h00;      memory[35098] <=  8'h00;      memory[35099] <=  8'h00;      memory[35100] <=  8'h00;      memory[35101] <=  8'h00;      memory[35102] <=  8'h00;      memory[35103] <=  8'h00;      memory[35104] <=  8'h00;      memory[35105] <=  8'h00;      memory[35106] <=  8'h00;      memory[35107] <=  8'h00;      memory[35108] <=  8'h00;      memory[35109] <=  8'h00;      memory[35110] <=  8'h00;      memory[35111] <=  8'h00;      memory[35112] <=  8'h00;      memory[35113] <=  8'h00;      memory[35114] <=  8'h00;      memory[35115] <=  8'h00;      memory[35116] <=  8'h00;      memory[35117] <=  8'h00;      memory[35118] <=  8'h00;      memory[35119] <=  8'h00;      memory[35120] <=  8'h00;      memory[35121] <=  8'h00;      memory[35122] <=  8'h00;      memory[35123] <=  8'h00;      memory[35124] <=  8'h00;      memory[35125] <=  8'h00;      memory[35126] <=  8'h00;      memory[35127] <=  8'h00;      memory[35128] <=  8'h00;      memory[35129] <=  8'h00;      memory[35130] <=  8'h00;      memory[35131] <=  8'h00;      memory[35132] <=  8'h00;      memory[35133] <=  8'h00;      memory[35134] <=  8'h00;      memory[35135] <=  8'h00;      memory[35136] <=  8'h00;      memory[35137] <=  8'h00;      memory[35138] <=  8'h00;      memory[35139] <=  8'h00;      memory[35140] <=  8'h00;      memory[35141] <=  8'h00;      memory[35142] <=  8'h00;      memory[35143] <=  8'h00;      memory[35144] <=  8'h00;      memory[35145] <=  8'h00;      memory[35146] <=  8'h00;      memory[35147] <=  8'h00;      memory[35148] <=  8'h00;      memory[35149] <=  8'h00;      memory[35150] <=  8'h00;      memory[35151] <=  8'h00;      memory[35152] <=  8'h00;      memory[35153] <=  8'h00;      memory[35154] <=  8'h00;      memory[35155] <=  8'h00;      memory[35156] <=  8'h00;      memory[35157] <=  8'h00;      memory[35158] <=  8'h00;      memory[35159] <=  8'h00;      memory[35160] <=  8'h00;      memory[35161] <=  8'h00;      memory[35162] <=  8'h00;      memory[35163] <=  8'h00;      memory[35164] <=  8'h00;      memory[35165] <=  8'h00;      memory[35166] <=  8'h00;      memory[35167] <=  8'h00;      memory[35168] <=  8'h00;      memory[35169] <=  8'h00;      memory[35170] <=  8'h00;      memory[35171] <=  8'h00;      memory[35172] <=  8'h00;      memory[35173] <=  8'h00;      memory[35174] <=  8'h00;      memory[35175] <=  8'h00;      memory[35176] <=  8'h00;      memory[35177] <=  8'h00;      memory[35178] <=  8'h00;      memory[35179] <=  8'h00;      memory[35180] <=  8'h00;      memory[35181] <=  8'h00;      memory[35182] <=  8'h00;      memory[35183] <=  8'h00;      memory[35184] <=  8'h00;      memory[35185] <=  8'h00;      memory[35186] <=  8'h00;      memory[35187] <=  8'h00;      memory[35188] <=  8'h00;      memory[35189] <=  8'h00;      memory[35190] <=  8'h00;      memory[35191] <=  8'h00;      memory[35192] <=  8'h00;      memory[35193] <=  8'h00;      memory[35194] <=  8'h00;      memory[35195] <=  8'h00;      memory[35196] <=  8'h00;      memory[35197] <=  8'h00;      memory[35198] <=  8'h00;      memory[35199] <=  8'h00;      memory[35200] <=  8'h00;      memory[35201] <=  8'h00;      memory[35202] <=  8'h00;      memory[35203] <=  8'h00;      memory[35204] <=  8'h00;      memory[35205] <=  8'h00;      memory[35206] <=  8'h00;      memory[35207] <=  8'h00;      memory[35208] <=  8'h00;      memory[35209] <=  8'h00;      memory[35210] <=  8'h00;      memory[35211] <=  8'h00;      memory[35212] <=  8'h00;      memory[35213] <=  8'h00;      memory[35214] <=  8'h00;      memory[35215] <=  8'h00;      memory[35216] <=  8'h00;      memory[35217] <=  8'h00;      memory[35218] <=  8'h00;      memory[35219] <=  8'h00;      memory[35220] <=  8'h00;      memory[35221] <=  8'h00;      memory[35222] <=  8'h00;      memory[35223] <=  8'h00;      memory[35224] <=  8'h00;      memory[35225] <=  8'h00;      memory[35226] <=  8'h00;      memory[35227] <=  8'h00;      memory[35228] <=  8'h00;      memory[35229] <=  8'h00;      memory[35230] <=  8'h00;      memory[35231] <=  8'h00;      memory[35232] <=  8'h00;      memory[35233] <=  8'h00;      memory[35234] <=  8'h00;      memory[35235] <=  8'h00;      memory[35236] <=  8'h00;      memory[35237] <=  8'h00;      memory[35238] <=  8'h00;      memory[35239] <=  8'h00;      memory[35240] <=  8'h00;      memory[35241] <=  8'h00;      memory[35242] <=  8'h00;      memory[35243] <=  8'h00;      memory[35244] <=  8'h00;      memory[35245] <=  8'h00;      memory[35246] <=  8'h00;      memory[35247] <=  8'h00;      memory[35248] <=  8'h00;      memory[35249] <=  8'h00;      memory[35250] <=  8'h00;      memory[35251] <=  8'h00;      memory[35252] <=  8'h00;      memory[35253] <=  8'h00;      memory[35254] <=  8'h00;      memory[35255] <=  8'h00;      memory[35256] <=  8'h00;      memory[35257] <=  8'h00;      memory[35258] <=  8'h00;      memory[35259] <=  8'h00;      memory[35260] <=  8'h00;      memory[35261] <=  8'h00;      memory[35262] <=  8'h00;      memory[35263] <=  8'h00;      memory[35264] <=  8'h00;      memory[35265] <=  8'h00;      memory[35266] <=  8'h00;      memory[35267] <=  8'h00;      memory[35268] <=  8'h00;      memory[35269] <=  8'h00;      memory[35270] <=  8'h00;      memory[35271] <=  8'h00;      memory[35272] <=  8'h00;      memory[35273] <=  8'h00;      memory[35274] <=  8'h00;      memory[35275] <=  8'h00;      memory[35276] <=  8'h00;      memory[35277] <=  8'h00;      memory[35278] <=  8'h00;      memory[35279] <=  8'h00;      memory[35280] <=  8'h00;      memory[35281] <=  8'h00;      memory[35282] <=  8'h00;      memory[35283] <=  8'h00;      memory[35284] <=  8'h00;      memory[35285] <=  8'h00;      memory[35286] <=  8'h00;      memory[35287] <=  8'h00;      memory[35288] <=  8'h00;      memory[35289] <=  8'h00;      memory[35290] <=  8'h00;      memory[35291] <=  8'h00;      memory[35292] <=  8'h00;      memory[35293] <=  8'h00;      memory[35294] <=  8'h00;      memory[35295] <=  8'h00;      memory[35296] <=  8'h00;      memory[35297] <=  8'h00;      memory[35298] <=  8'h00;      memory[35299] <=  8'h00;      memory[35300] <=  8'h00;      memory[35301] <=  8'h00;      memory[35302] <=  8'h00;      memory[35303] <=  8'h00;      memory[35304] <=  8'h00;      memory[35305] <=  8'h00;      memory[35306] <=  8'h00;      memory[35307] <=  8'h00;      memory[35308] <=  8'h00;      memory[35309] <=  8'h00;      memory[35310] <=  8'h00;      memory[35311] <=  8'h00;      memory[35312] <=  8'h00;      memory[35313] <=  8'h00;      memory[35314] <=  8'h00;      memory[35315] <=  8'h00;      memory[35316] <=  8'h00;      memory[35317] <=  8'h00;      memory[35318] <=  8'h00;      memory[35319] <=  8'h00;      memory[35320] <=  8'h00;      memory[35321] <=  8'h00;      memory[35322] <=  8'h00;      memory[35323] <=  8'h00;      memory[35324] <=  8'h00;      memory[35325] <=  8'h00;      memory[35326] <=  8'h00;      memory[35327] <=  8'h00;      memory[35328] <=  8'h00;      memory[35329] <=  8'h00;      memory[35330] <=  8'h00;      memory[35331] <=  8'h00;      memory[35332] <=  8'h00;      memory[35333] <=  8'h00;      memory[35334] <=  8'h00;      memory[35335] <=  8'h00;      memory[35336] <=  8'h00;      memory[35337] <=  8'h00;      memory[35338] <=  8'h00;      memory[35339] <=  8'h00;      memory[35340] <=  8'h00;      memory[35341] <=  8'h00;      memory[35342] <=  8'h00;      memory[35343] <=  8'h00;      memory[35344] <=  8'h00;      memory[35345] <=  8'h00;      memory[35346] <=  8'h00;      memory[35347] <=  8'h00;      memory[35348] <=  8'h00;      memory[35349] <=  8'h00;      memory[35350] <=  8'h00;      memory[35351] <=  8'h00;      memory[35352] <=  8'h00;      memory[35353] <=  8'h00;      memory[35354] <=  8'h00;      memory[35355] <=  8'h00;      memory[35356] <=  8'h00;      memory[35357] <=  8'h00;      memory[35358] <=  8'h00;      memory[35359] <=  8'h00;      memory[35360] <=  8'h00;      memory[35361] <=  8'h00;      memory[35362] <=  8'h00;      memory[35363] <=  8'h00;      memory[35364] <=  8'h00;      memory[35365] <=  8'h00;      memory[35366] <=  8'h00;      memory[35367] <=  8'h00;      memory[35368] <=  8'h00;      memory[35369] <=  8'h00;      memory[35370] <=  8'h00;      memory[35371] <=  8'h00;      memory[35372] <=  8'h00;      memory[35373] <=  8'h00;      memory[35374] <=  8'h00;      memory[35375] <=  8'h00;      memory[35376] <=  8'h00;      memory[35377] <=  8'h00;      memory[35378] <=  8'h00;      memory[35379] <=  8'h00;      memory[35380] <=  8'h00;      memory[35381] <=  8'h00;      memory[35382] <=  8'h00;      memory[35383] <=  8'h00;      memory[35384] <=  8'h00;      memory[35385] <=  8'h00;      memory[35386] <=  8'h00;      memory[35387] <=  8'h00;      memory[35388] <=  8'h00;      memory[35389] <=  8'h00;      memory[35390] <=  8'h00;      memory[35391] <=  8'h00;      memory[35392] <=  8'h00;      memory[35393] <=  8'h00;      memory[35394] <=  8'h00;      memory[35395] <=  8'h00;      memory[35396] <=  8'h00;      memory[35397] <=  8'h00;      memory[35398] <=  8'h00;      memory[35399] <=  8'h00;      memory[35400] <=  8'h00;      memory[35401] <=  8'h00;      memory[35402] <=  8'h00;      memory[35403] <=  8'h00;      memory[35404] <=  8'h00;      memory[35405] <=  8'h00;      memory[35406] <=  8'h00;      memory[35407] <=  8'h00;      memory[35408] <=  8'h00;      memory[35409] <=  8'h00;      memory[35410] <=  8'h00;      memory[35411] <=  8'h00;      memory[35412] <=  8'h00;      memory[35413] <=  8'h00;      memory[35414] <=  8'h00;      memory[35415] <=  8'h00;      memory[35416] <=  8'h00;      memory[35417] <=  8'h00;      memory[35418] <=  8'h00;      memory[35419] <=  8'h00;      memory[35420] <=  8'h00;      memory[35421] <=  8'h00;      memory[35422] <=  8'h00;      memory[35423] <=  8'h00;      memory[35424] <=  8'h00;      memory[35425] <=  8'h00;      memory[35426] <=  8'h00;      memory[35427] <=  8'h00;      memory[35428] <=  8'h00;      memory[35429] <=  8'h00;      memory[35430] <=  8'h00;      memory[35431] <=  8'h00;      memory[35432] <=  8'h00;      memory[35433] <=  8'h00;      memory[35434] <=  8'h00;      memory[35435] <=  8'h00;      memory[35436] <=  8'h00;      memory[35437] <=  8'h00;      memory[35438] <=  8'h00;      memory[35439] <=  8'h00;      memory[35440] <=  8'h00;      memory[35441] <=  8'h00;      memory[35442] <=  8'h00;      memory[35443] <=  8'h00;      memory[35444] <=  8'h00;      memory[35445] <=  8'h00;      memory[35446] <=  8'h00;      memory[35447] <=  8'h00;      memory[35448] <=  8'h00;      memory[35449] <=  8'h00;      memory[35450] <=  8'h00;      memory[35451] <=  8'h00;      memory[35452] <=  8'h00;      memory[35453] <=  8'h00;      memory[35454] <=  8'h00;      memory[35455] <=  8'h00;      memory[35456] <=  8'h00;      memory[35457] <=  8'h00;      memory[35458] <=  8'h00;      memory[35459] <=  8'h00;      memory[35460] <=  8'h00;      memory[35461] <=  8'h00;      memory[35462] <=  8'h00;      memory[35463] <=  8'h00;      memory[35464] <=  8'h00;      memory[35465] <=  8'h00;      memory[35466] <=  8'h00;      memory[35467] <=  8'h00;      memory[35468] <=  8'h00;      memory[35469] <=  8'h00;      memory[35470] <=  8'h00;      memory[35471] <=  8'h00;      memory[35472] <=  8'h00;      memory[35473] <=  8'h00;      memory[35474] <=  8'h00;      memory[35475] <=  8'h00;      memory[35476] <=  8'h00;      memory[35477] <=  8'h00;      memory[35478] <=  8'h00;      memory[35479] <=  8'h00;      memory[35480] <=  8'h00;      memory[35481] <=  8'h00;      memory[35482] <=  8'h00;      memory[35483] <=  8'h00;      memory[35484] <=  8'h00;      memory[35485] <=  8'h00;      memory[35486] <=  8'h00;      memory[35487] <=  8'h00;      memory[35488] <=  8'h00;      memory[35489] <=  8'h00;      memory[35490] <=  8'h00;      memory[35491] <=  8'h00;      memory[35492] <=  8'h00;      memory[35493] <=  8'h00;      memory[35494] <=  8'h00;      memory[35495] <=  8'h00;      memory[35496] <=  8'h00;      memory[35497] <=  8'h00;      memory[35498] <=  8'h00;      memory[35499] <=  8'h00;      memory[35500] <=  8'h00;      memory[35501] <=  8'h00;      memory[35502] <=  8'h00;      memory[35503] <=  8'h00;      memory[35504] <=  8'h00;      memory[35505] <=  8'h00;      memory[35506] <=  8'h00;      memory[35507] <=  8'h00;      memory[35508] <=  8'h00;      memory[35509] <=  8'h00;      memory[35510] <=  8'h00;      memory[35511] <=  8'h00;      memory[35512] <=  8'h00;      memory[35513] <=  8'h00;      memory[35514] <=  8'h00;      memory[35515] <=  8'h00;      memory[35516] <=  8'h00;      memory[35517] <=  8'h00;      memory[35518] <=  8'h00;      memory[35519] <=  8'h00;      memory[35520] <=  8'h00;      memory[35521] <=  8'h00;      memory[35522] <=  8'h00;      memory[35523] <=  8'h00;      memory[35524] <=  8'h00;      memory[35525] <=  8'h00;      memory[35526] <=  8'h00;      memory[35527] <=  8'h00;      memory[35528] <=  8'h00;      memory[35529] <=  8'h00;      memory[35530] <=  8'h00;      memory[35531] <=  8'h00;      memory[35532] <=  8'h00;      memory[35533] <=  8'h00;      memory[35534] <=  8'h00;      memory[35535] <=  8'h00;      memory[35536] <=  8'h00;      memory[35537] <=  8'h00;      memory[35538] <=  8'h00;      memory[35539] <=  8'h00;      memory[35540] <=  8'h00;      memory[35541] <=  8'h00;      memory[35542] <=  8'h00;      memory[35543] <=  8'h00;      memory[35544] <=  8'h00;      memory[35545] <=  8'h00;      memory[35546] <=  8'h00;      memory[35547] <=  8'h00;      memory[35548] <=  8'h00;      memory[35549] <=  8'h00;      memory[35550] <=  8'h00;      memory[35551] <=  8'h00;      memory[35552] <=  8'h00;      memory[35553] <=  8'h00;      memory[35554] <=  8'h00;      memory[35555] <=  8'h00;      memory[35556] <=  8'h00;      memory[35557] <=  8'h00;      memory[35558] <=  8'h00;      memory[35559] <=  8'h00;      memory[35560] <=  8'h00;      memory[35561] <=  8'h00;      memory[35562] <=  8'h00;      memory[35563] <=  8'h00;      memory[35564] <=  8'h00;      memory[35565] <=  8'h00;      memory[35566] <=  8'h00;      memory[35567] <=  8'h00;      memory[35568] <=  8'h00;      memory[35569] <=  8'h00;      memory[35570] <=  8'h00;      memory[35571] <=  8'h00;      memory[35572] <=  8'h00;      memory[35573] <=  8'h00;      memory[35574] <=  8'h00;      memory[35575] <=  8'h00;      memory[35576] <=  8'h00;      memory[35577] <=  8'h00;      memory[35578] <=  8'h00;      memory[35579] <=  8'h00;      memory[35580] <=  8'h00;      memory[35581] <=  8'h00;      memory[35582] <=  8'h00;      memory[35583] <=  8'h00;      memory[35584] <=  8'h00;      memory[35585] <=  8'h00;      memory[35586] <=  8'h00;      memory[35587] <=  8'h00;      memory[35588] <=  8'h00;      memory[35589] <=  8'h00;      memory[35590] <=  8'h00;      memory[35591] <=  8'h00;      memory[35592] <=  8'h00;      memory[35593] <=  8'h00;      memory[35594] <=  8'h00;      memory[35595] <=  8'h00;      memory[35596] <=  8'h00;      memory[35597] <=  8'h00;      memory[35598] <=  8'h00;      memory[35599] <=  8'h00;      memory[35600] <=  8'h00;      memory[35601] <=  8'h00;      memory[35602] <=  8'h00;      memory[35603] <=  8'h00;      memory[35604] <=  8'h00;      memory[35605] <=  8'h00;      memory[35606] <=  8'h00;      memory[35607] <=  8'h00;      memory[35608] <=  8'h00;      memory[35609] <=  8'h00;      memory[35610] <=  8'h00;      memory[35611] <=  8'h00;      memory[35612] <=  8'h00;      memory[35613] <=  8'h00;      memory[35614] <=  8'h00;      memory[35615] <=  8'h00;      memory[35616] <=  8'h00;      memory[35617] <=  8'h00;      memory[35618] <=  8'h00;      memory[35619] <=  8'h00;      memory[35620] <=  8'h00;      memory[35621] <=  8'h00;      memory[35622] <=  8'h00;      memory[35623] <=  8'h00;      memory[35624] <=  8'h00;      memory[35625] <=  8'h00;      memory[35626] <=  8'h00;      memory[35627] <=  8'h00;      memory[35628] <=  8'h00;      memory[35629] <=  8'h00;      memory[35630] <=  8'h00;      memory[35631] <=  8'h00;      memory[35632] <=  8'h00;      memory[35633] <=  8'h00;      memory[35634] <=  8'h00;      memory[35635] <=  8'h00;      memory[35636] <=  8'h00;      memory[35637] <=  8'h00;      memory[35638] <=  8'h00;      memory[35639] <=  8'h00;      memory[35640] <=  8'h00;      memory[35641] <=  8'h00;      memory[35642] <=  8'h00;      memory[35643] <=  8'h00;      memory[35644] <=  8'h00;      memory[35645] <=  8'h00;      memory[35646] <=  8'h00;      memory[35647] <=  8'h00;      memory[35648] <=  8'h00;      memory[35649] <=  8'h00;      memory[35650] <=  8'h00;      memory[35651] <=  8'h00;      memory[35652] <=  8'h00;      memory[35653] <=  8'h00;      memory[35654] <=  8'h00;      memory[35655] <=  8'h00;      memory[35656] <=  8'h00;      memory[35657] <=  8'h00;      memory[35658] <=  8'h00;      memory[35659] <=  8'h00;      memory[35660] <=  8'h00;      memory[35661] <=  8'h00;      memory[35662] <=  8'h00;      memory[35663] <=  8'h00;      memory[35664] <=  8'h00;      memory[35665] <=  8'h00;      memory[35666] <=  8'h00;      memory[35667] <=  8'h00;      memory[35668] <=  8'h00;      memory[35669] <=  8'h00;      memory[35670] <=  8'h00;      memory[35671] <=  8'h00;      memory[35672] <=  8'h00;      memory[35673] <=  8'h00;      memory[35674] <=  8'h00;      memory[35675] <=  8'h00;      memory[35676] <=  8'h00;      memory[35677] <=  8'h00;      memory[35678] <=  8'h00;      memory[35679] <=  8'h00;      memory[35680] <=  8'h00;      memory[35681] <=  8'h00;      memory[35682] <=  8'h00;      memory[35683] <=  8'h00;      memory[35684] <=  8'h00;      memory[35685] <=  8'h00;      memory[35686] <=  8'h00;      memory[35687] <=  8'h00;      memory[35688] <=  8'h00;      memory[35689] <=  8'h00;      memory[35690] <=  8'h00;      memory[35691] <=  8'h00;      memory[35692] <=  8'h00;      memory[35693] <=  8'h00;      memory[35694] <=  8'h00;      memory[35695] <=  8'h00;      memory[35696] <=  8'h00;      memory[35697] <=  8'h00;      memory[35698] <=  8'h00;      memory[35699] <=  8'h00;      memory[35700] <=  8'h00;      memory[35701] <=  8'h00;      memory[35702] <=  8'h00;      memory[35703] <=  8'h00;      memory[35704] <=  8'h00;      memory[35705] <=  8'h00;      memory[35706] <=  8'h00;      memory[35707] <=  8'h00;      memory[35708] <=  8'h00;      memory[35709] <=  8'h00;      memory[35710] <=  8'h00;      memory[35711] <=  8'h00;      memory[35712] <=  8'h00;      memory[35713] <=  8'h00;      memory[35714] <=  8'h00;      memory[35715] <=  8'h00;      memory[35716] <=  8'h00;      memory[35717] <=  8'h00;      memory[35718] <=  8'h00;      memory[35719] <=  8'h00;      memory[35720] <=  8'h00;      memory[35721] <=  8'h00;      memory[35722] <=  8'h00;      memory[35723] <=  8'h00;      memory[35724] <=  8'h00;      memory[35725] <=  8'h00;      memory[35726] <=  8'h00;      memory[35727] <=  8'h00;      memory[35728] <=  8'h00;      memory[35729] <=  8'h00;      memory[35730] <=  8'h00;      memory[35731] <=  8'h00;      memory[35732] <=  8'h00;      memory[35733] <=  8'h00;      memory[35734] <=  8'h00;      memory[35735] <=  8'h00;      memory[35736] <=  8'h00;      memory[35737] <=  8'h00;      memory[35738] <=  8'h00;      memory[35739] <=  8'h00;      memory[35740] <=  8'h00;      memory[35741] <=  8'h00;      memory[35742] <=  8'h00;      memory[35743] <=  8'h00;      memory[35744] <=  8'h00;      memory[35745] <=  8'h00;      memory[35746] <=  8'h00;      memory[35747] <=  8'h00;      memory[35748] <=  8'h00;      memory[35749] <=  8'h00;      memory[35750] <=  8'h00;      memory[35751] <=  8'h00;      memory[35752] <=  8'h00;      memory[35753] <=  8'h00;      memory[35754] <=  8'h00;      memory[35755] <=  8'h00;      memory[35756] <=  8'h00;      memory[35757] <=  8'h00;      memory[35758] <=  8'h00;      memory[35759] <=  8'h00;      memory[35760] <=  8'h00;      memory[35761] <=  8'h00;      memory[35762] <=  8'h00;      memory[35763] <=  8'h00;      memory[35764] <=  8'h00;      memory[35765] <=  8'h00;      memory[35766] <=  8'h00;      memory[35767] <=  8'h00;      memory[35768] <=  8'h00;      memory[35769] <=  8'h00;      memory[35770] <=  8'h00;      memory[35771] <=  8'h00;      memory[35772] <=  8'h00;      memory[35773] <=  8'h00;      memory[35774] <=  8'h00;      memory[35775] <=  8'h00;      memory[35776] <=  8'h00;      memory[35777] <=  8'h00;      memory[35778] <=  8'h00;      memory[35779] <=  8'h00;      memory[35780] <=  8'h00;      memory[35781] <=  8'h00;      memory[35782] <=  8'h00;      memory[35783] <=  8'h00;      memory[35784] <=  8'h00;      memory[35785] <=  8'h00;      memory[35786] <=  8'h00;      memory[35787] <=  8'h00;      memory[35788] <=  8'h00;      memory[35789] <=  8'h00;      memory[35790] <=  8'h00;      memory[35791] <=  8'h00;      memory[35792] <=  8'h00;      memory[35793] <=  8'h00;      memory[35794] <=  8'h00;      memory[35795] <=  8'h00;      memory[35796] <=  8'h00;      memory[35797] <=  8'h00;      memory[35798] <=  8'h00;      memory[35799] <=  8'h00;      memory[35800] <=  8'h00;      memory[35801] <=  8'h00;      memory[35802] <=  8'h00;      memory[35803] <=  8'h00;      memory[35804] <=  8'h00;      memory[35805] <=  8'h00;      memory[35806] <=  8'h00;      memory[35807] <=  8'h00;      memory[35808] <=  8'h00;      memory[35809] <=  8'h00;      memory[35810] <=  8'h00;      memory[35811] <=  8'h00;      memory[35812] <=  8'h00;      memory[35813] <=  8'h00;      memory[35814] <=  8'h00;      memory[35815] <=  8'h00;      memory[35816] <=  8'h00;      memory[35817] <=  8'h00;      memory[35818] <=  8'h00;      memory[35819] <=  8'h00;      memory[35820] <=  8'h00;      memory[35821] <=  8'h00;      memory[35822] <=  8'h00;      memory[35823] <=  8'h00;      memory[35824] <=  8'h00;      memory[35825] <=  8'h00;      memory[35826] <=  8'h00;      memory[35827] <=  8'h00;      memory[35828] <=  8'h00;      memory[35829] <=  8'h00;      memory[35830] <=  8'h00;      memory[35831] <=  8'h00;      memory[35832] <=  8'h00;      memory[35833] <=  8'h00;      memory[35834] <=  8'h00;      memory[35835] <=  8'h00;      memory[35836] <=  8'h00;      memory[35837] <=  8'h00;      memory[35838] <=  8'h00;      memory[35839] <=  8'h00;      memory[35840] <=  8'h00;      memory[35841] <=  8'h00;      memory[35842] <=  8'h00;      memory[35843] <=  8'h00;      memory[35844] <=  8'h00;      memory[35845] <=  8'h00;      memory[35846] <=  8'h00;      memory[35847] <=  8'h00;      memory[35848] <=  8'h00;      memory[35849] <=  8'h00;      memory[35850] <=  8'h00;      memory[35851] <=  8'h00;      memory[35852] <=  8'h00;      memory[35853] <=  8'h00;      memory[35854] <=  8'h00;      memory[35855] <=  8'h00;      memory[35856] <=  8'h00;      memory[35857] <=  8'h00;      memory[35858] <=  8'h00;      memory[35859] <=  8'h00;      memory[35860] <=  8'h00;      memory[35861] <=  8'h00;      memory[35862] <=  8'h00;      memory[35863] <=  8'h00;      memory[35864] <=  8'h00;      memory[35865] <=  8'h00;      memory[35866] <=  8'h00;      memory[35867] <=  8'h00;      memory[35868] <=  8'h00;      memory[35869] <=  8'h00;      memory[35870] <=  8'h00;      memory[35871] <=  8'h00;      memory[35872] <=  8'h00;      memory[35873] <=  8'h00;      memory[35874] <=  8'h00;      memory[35875] <=  8'h00;      memory[35876] <=  8'h00;      memory[35877] <=  8'h00;      memory[35878] <=  8'h00;      memory[35879] <=  8'h00;      memory[35880] <=  8'h00;      memory[35881] <=  8'h00;      memory[35882] <=  8'h00;      memory[35883] <=  8'h00;      memory[35884] <=  8'h00;      memory[35885] <=  8'h00;      memory[35886] <=  8'h00;      memory[35887] <=  8'h00;      memory[35888] <=  8'h00;      memory[35889] <=  8'h00;      memory[35890] <=  8'h00;      memory[35891] <=  8'h00;      memory[35892] <=  8'h00;      memory[35893] <=  8'h00;      memory[35894] <=  8'h00;      memory[35895] <=  8'h00;      memory[35896] <=  8'h00;      memory[35897] <=  8'h00;      memory[35898] <=  8'h00;      memory[35899] <=  8'h00;      memory[35900] <=  8'h00;      memory[35901] <=  8'h00;      memory[35902] <=  8'h00;      memory[35903] <=  8'h00;      memory[35904] <=  8'h00;      memory[35905] <=  8'h00;      memory[35906] <=  8'h00;      memory[35907] <=  8'h00;      memory[35908] <=  8'h00;      memory[35909] <=  8'h00;      memory[35910] <=  8'h00;      memory[35911] <=  8'h00;      memory[35912] <=  8'h00;      memory[35913] <=  8'h00;      memory[35914] <=  8'h00;      memory[35915] <=  8'h00;      memory[35916] <=  8'h00;      memory[35917] <=  8'h00;      memory[35918] <=  8'h00;      memory[35919] <=  8'h00;      memory[35920] <=  8'h00;      memory[35921] <=  8'h00;      memory[35922] <=  8'h00;      memory[35923] <=  8'h00;      memory[35924] <=  8'h00;      memory[35925] <=  8'h00;      memory[35926] <=  8'h00;      memory[35927] <=  8'h00;      memory[35928] <=  8'h00;      memory[35929] <=  8'h00;      memory[35930] <=  8'h00;      memory[35931] <=  8'h00;      memory[35932] <=  8'h00;      memory[35933] <=  8'h00;      memory[35934] <=  8'h00;      memory[35935] <=  8'h00;      memory[35936] <=  8'h00;      memory[35937] <=  8'h00;      memory[35938] <=  8'h00;      memory[35939] <=  8'h00;      memory[35940] <=  8'h00;      memory[35941] <=  8'h00;      memory[35942] <=  8'h00;      memory[35943] <=  8'h00;      memory[35944] <=  8'h00;      memory[35945] <=  8'h00;      memory[35946] <=  8'h00;      memory[35947] <=  8'h00;      memory[35948] <=  8'h00;      memory[35949] <=  8'h00;      memory[35950] <=  8'h00;      memory[35951] <=  8'h00;      memory[35952] <=  8'h00;      memory[35953] <=  8'h00;      memory[35954] <=  8'h00;      memory[35955] <=  8'h00;      memory[35956] <=  8'h00;      memory[35957] <=  8'h00;      memory[35958] <=  8'h00;      memory[35959] <=  8'h00;      memory[35960] <=  8'h00;      memory[35961] <=  8'h00;      memory[35962] <=  8'h00;      memory[35963] <=  8'h00;      memory[35964] <=  8'h00;      memory[35965] <=  8'h00;      memory[35966] <=  8'h00;      memory[35967] <=  8'h00;      memory[35968] <=  8'h00;      memory[35969] <=  8'h00;      memory[35970] <=  8'h00;      memory[35971] <=  8'h00;      memory[35972] <=  8'h00;      memory[35973] <=  8'h00;      memory[35974] <=  8'h00;      memory[35975] <=  8'h00;      memory[35976] <=  8'h00;      memory[35977] <=  8'h00;      memory[35978] <=  8'h00;      memory[35979] <=  8'h00;      memory[35980] <=  8'h00;      memory[35981] <=  8'h00;      memory[35982] <=  8'h00;      memory[35983] <=  8'h00;      memory[35984] <=  8'h00;      memory[35985] <=  8'h00;      memory[35986] <=  8'h00;      memory[35987] <=  8'h00;      memory[35988] <=  8'h00;      memory[35989] <=  8'h00;      memory[35990] <=  8'h00;      memory[35991] <=  8'h00;      memory[35992] <=  8'h00;      memory[35993] <=  8'h00;      memory[35994] <=  8'h00;      memory[35995] <=  8'h00;      memory[35996] <=  8'h00;      memory[35997] <=  8'h00;      memory[35998] <=  8'h00;      memory[35999] <=  8'h00;      memory[36000] <=  8'h00;      memory[36001] <=  8'h00;      memory[36002] <=  8'h00;      memory[36003] <=  8'h00;      memory[36004] <=  8'h00;      memory[36005] <=  8'h00;      memory[36006] <=  8'h00;      memory[36007] <=  8'h00;      memory[36008] <=  8'h00;      memory[36009] <=  8'h00;      memory[36010] <=  8'h00;      memory[36011] <=  8'h00;      memory[36012] <=  8'h00;      memory[36013] <=  8'h00;      memory[36014] <=  8'h00;      memory[36015] <=  8'h00;      memory[36016] <=  8'h00;      memory[36017] <=  8'h00;      memory[36018] <=  8'h00;      memory[36019] <=  8'h00;      memory[36020] <=  8'h00;      memory[36021] <=  8'h00;      memory[36022] <=  8'h00;      memory[36023] <=  8'h00;      memory[36024] <=  8'h00;      memory[36025] <=  8'h00;      memory[36026] <=  8'h00;      memory[36027] <=  8'h00;      memory[36028] <=  8'h00;      memory[36029] <=  8'h00;      memory[36030] <=  8'h00;      memory[36031] <=  8'h00;      memory[36032] <=  8'h00;      memory[36033] <=  8'h00;      memory[36034] <=  8'h00;      memory[36035] <=  8'h00;      memory[36036] <=  8'h00;      memory[36037] <=  8'h00;      memory[36038] <=  8'h00;      memory[36039] <=  8'h00;      memory[36040] <=  8'h00;      memory[36041] <=  8'h00;      memory[36042] <=  8'h00;      memory[36043] <=  8'h00;      memory[36044] <=  8'h00;      memory[36045] <=  8'h00;      memory[36046] <=  8'h00;      memory[36047] <=  8'h00;      memory[36048] <=  8'h00;      memory[36049] <=  8'h00;      memory[36050] <=  8'h00;      memory[36051] <=  8'h00;      memory[36052] <=  8'h00;      memory[36053] <=  8'h00;      memory[36054] <=  8'h00;      memory[36055] <=  8'h00;      memory[36056] <=  8'h00;      memory[36057] <=  8'h00;      memory[36058] <=  8'h00;      memory[36059] <=  8'h00;      memory[36060] <=  8'h00;      memory[36061] <=  8'h00;      memory[36062] <=  8'h00;      memory[36063] <=  8'h00;      memory[36064] <=  8'h00;      memory[36065] <=  8'h00;      memory[36066] <=  8'h00;      memory[36067] <=  8'h00;      memory[36068] <=  8'h00;      memory[36069] <=  8'h00;      memory[36070] <=  8'h00;      memory[36071] <=  8'h00;      memory[36072] <=  8'h00;      memory[36073] <=  8'h00;      memory[36074] <=  8'h00;      memory[36075] <=  8'h00;      memory[36076] <=  8'h00;      memory[36077] <=  8'h00;      memory[36078] <=  8'h00;      memory[36079] <=  8'h00;      memory[36080] <=  8'h00;      memory[36081] <=  8'h00;      memory[36082] <=  8'h00;      memory[36083] <=  8'h00;      memory[36084] <=  8'h00;      memory[36085] <=  8'h00;      memory[36086] <=  8'h00;      memory[36087] <=  8'h00;      memory[36088] <=  8'h00;      memory[36089] <=  8'h00;      memory[36090] <=  8'h00;      memory[36091] <=  8'h00;      memory[36092] <=  8'h00;      memory[36093] <=  8'h00;      memory[36094] <=  8'h00;      memory[36095] <=  8'h00;      memory[36096] <=  8'h00;      memory[36097] <=  8'h00;      memory[36098] <=  8'h00;      memory[36099] <=  8'h00;      memory[36100] <=  8'h00;      memory[36101] <=  8'h00;      memory[36102] <=  8'h00;      memory[36103] <=  8'h00;      memory[36104] <=  8'h00;      memory[36105] <=  8'h00;      memory[36106] <=  8'h00;      memory[36107] <=  8'h00;      memory[36108] <=  8'h00;      memory[36109] <=  8'h00;      memory[36110] <=  8'h00;      memory[36111] <=  8'h00;      memory[36112] <=  8'h00;      memory[36113] <=  8'h00;      memory[36114] <=  8'h00;      memory[36115] <=  8'h00;      memory[36116] <=  8'h00;      memory[36117] <=  8'h00;      memory[36118] <=  8'h00;      memory[36119] <=  8'h00;      memory[36120] <=  8'h00;      memory[36121] <=  8'h00;      memory[36122] <=  8'h00;      memory[36123] <=  8'h00;      memory[36124] <=  8'h00;      memory[36125] <=  8'h00;      memory[36126] <=  8'h00;      memory[36127] <=  8'h00;      memory[36128] <=  8'h00;      memory[36129] <=  8'h00;      memory[36130] <=  8'h00;      memory[36131] <=  8'h00;      memory[36132] <=  8'h00;      memory[36133] <=  8'h00;      memory[36134] <=  8'h00;      memory[36135] <=  8'h00;      memory[36136] <=  8'h00;      memory[36137] <=  8'h00;      memory[36138] <=  8'h00;      memory[36139] <=  8'h00;      memory[36140] <=  8'h00;      memory[36141] <=  8'h00;      memory[36142] <=  8'h00;      memory[36143] <=  8'h00;      memory[36144] <=  8'h00;      memory[36145] <=  8'h00;      memory[36146] <=  8'h00;      memory[36147] <=  8'h00;      memory[36148] <=  8'h00;      memory[36149] <=  8'h00;      memory[36150] <=  8'h00;      memory[36151] <=  8'h00;      memory[36152] <=  8'h00;      memory[36153] <=  8'h00;      memory[36154] <=  8'h00;      memory[36155] <=  8'h00;      memory[36156] <=  8'h00;      memory[36157] <=  8'h00;      memory[36158] <=  8'h00;      memory[36159] <=  8'h00;      memory[36160] <=  8'h00;      memory[36161] <=  8'h00;      memory[36162] <=  8'h00;      memory[36163] <=  8'h00;      memory[36164] <=  8'h00;      memory[36165] <=  8'h00;      memory[36166] <=  8'h00;      memory[36167] <=  8'h00;      memory[36168] <=  8'h00;      memory[36169] <=  8'h00;      memory[36170] <=  8'h00;      memory[36171] <=  8'h00;      memory[36172] <=  8'h00;      memory[36173] <=  8'h00;      memory[36174] <=  8'h00;      memory[36175] <=  8'h00;      memory[36176] <=  8'h00;      memory[36177] <=  8'h00;      memory[36178] <=  8'h00;      memory[36179] <=  8'h00;      memory[36180] <=  8'h00;      memory[36181] <=  8'h00;      memory[36182] <=  8'h00;      memory[36183] <=  8'h00;      memory[36184] <=  8'h00;      memory[36185] <=  8'h00;      memory[36186] <=  8'h00;      memory[36187] <=  8'h00;      memory[36188] <=  8'h00;      memory[36189] <=  8'h00;      memory[36190] <=  8'h00;      memory[36191] <=  8'h00;      memory[36192] <=  8'h00;      memory[36193] <=  8'h00;      memory[36194] <=  8'h00;      memory[36195] <=  8'h00;      memory[36196] <=  8'h00;      memory[36197] <=  8'h00;      memory[36198] <=  8'h00;      memory[36199] <=  8'h00;      memory[36200] <=  8'h00;      memory[36201] <=  8'h00;      memory[36202] <=  8'h00;      memory[36203] <=  8'h00;      memory[36204] <=  8'h00;      memory[36205] <=  8'h00;      memory[36206] <=  8'h00;      memory[36207] <=  8'h00;      memory[36208] <=  8'h00;      memory[36209] <=  8'h00;      memory[36210] <=  8'h00;      memory[36211] <=  8'h00;      memory[36212] <=  8'h00;      memory[36213] <=  8'h00;      memory[36214] <=  8'h00;      memory[36215] <=  8'h00;      memory[36216] <=  8'h00;      memory[36217] <=  8'h00;      memory[36218] <=  8'h00;      memory[36219] <=  8'h00;      memory[36220] <=  8'h00;      memory[36221] <=  8'h00;      memory[36222] <=  8'h00;      memory[36223] <=  8'h00;      memory[36224] <=  8'h00;      memory[36225] <=  8'h00;      memory[36226] <=  8'h00;      memory[36227] <=  8'h00;      memory[36228] <=  8'h00;      memory[36229] <=  8'h00;      memory[36230] <=  8'h00;      memory[36231] <=  8'h00;      memory[36232] <=  8'h00;      memory[36233] <=  8'h00;      memory[36234] <=  8'h00;      memory[36235] <=  8'h00;      memory[36236] <=  8'h00;      memory[36237] <=  8'h00;      memory[36238] <=  8'h00;      memory[36239] <=  8'h00;      memory[36240] <=  8'h00;      memory[36241] <=  8'h00;      memory[36242] <=  8'h00;      memory[36243] <=  8'h00;      memory[36244] <=  8'h00;      memory[36245] <=  8'h00;      memory[36246] <=  8'h00;      memory[36247] <=  8'h00;      memory[36248] <=  8'h00;      memory[36249] <=  8'h00;      memory[36250] <=  8'h00;      memory[36251] <=  8'h00;      memory[36252] <=  8'h00;      memory[36253] <=  8'h00;      memory[36254] <=  8'h00;      memory[36255] <=  8'h00;      memory[36256] <=  8'h00;      memory[36257] <=  8'h00;      memory[36258] <=  8'h00;      memory[36259] <=  8'h00;      memory[36260] <=  8'h00;      memory[36261] <=  8'h00;      memory[36262] <=  8'h00;      memory[36263] <=  8'h00;      memory[36264] <=  8'h00;      memory[36265] <=  8'h00;      memory[36266] <=  8'h00;      memory[36267] <=  8'h00;      memory[36268] <=  8'h00;      memory[36269] <=  8'h00;      memory[36270] <=  8'h00;      memory[36271] <=  8'h00;      memory[36272] <=  8'h00;      memory[36273] <=  8'h00;      memory[36274] <=  8'h00;      memory[36275] <=  8'h00;      memory[36276] <=  8'h00;      memory[36277] <=  8'h00;      memory[36278] <=  8'h00;      memory[36279] <=  8'h00;      memory[36280] <=  8'h00;      memory[36281] <=  8'h00;      memory[36282] <=  8'h00;      memory[36283] <=  8'h00;      memory[36284] <=  8'h00;      memory[36285] <=  8'h00;      memory[36286] <=  8'h00;      memory[36287] <=  8'h00;      memory[36288] <=  8'h00;      memory[36289] <=  8'h00;      memory[36290] <=  8'h00;      memory[36291] <=  8'h00;      memory[36292] <=  8'h00;      memory[36293] <=  8'h00;      memory[36294] <=  8'h00;      memory[36295] <=  8'h00;      memory[36296] <=  8'h00;      memory[36297] <=  8'h00;      memory[36298] <=  8'h00;      memory[36299] <=  8'h00;      memory[36300] <=  8'h00;      memory[36301] <=  8'h00;      memory[36302] <=  8'h00;      memory[36303] <=  8'h00;      memory[36304] <=  8'h00;      memory[36305] <=  8'h00;      memory[36306] <=  8'h00;      memory[36307] <=  8'h00;      memory[36308] <=  8'h00;      memory[36309] <=  8'h00;      memory[36310] <=  8'h00;      memory[36311] <=  8'h00;      memory[36312] <=  8'h00;      memory[36313] <=  8'h00;      memory[36314] <=  8'h00;      memory[36315] <=  8'h00;      memory[36316] <=  8'h00;      memory[36317] <=  8'h00;      memory[36318] <=  8'h00;      memory[36319] <=  8'h00;      memory[36320] <=  8'h00;      memory[36321] <=  8'h00;      memory[36322] <=  8'h00;      memory[36323] <=  8'h00;      memory[36324] <=  8'h00;      memory[36325] <=  8'h00;      memory[36326] <=  8'h00;      memory[36327] <=  8'h00;      memory[36328] <=  8'h00;      memory[36329] <=  8'h00;      memory[36330] <=  8'h00;      memory[36331] <=  8'h00;      memory[36332] <=  8'h00;      memory[36333] <=  8'h00;      memory[36334] <=  8'h00;      memory[36335] <=  8'h00;      memory[36336] <=  8'h00;      memory[36337] <=  8'h00;      memory[36338] <=  8'h00;      memory[36339] <=  8'h00;      memory[36340] <=  8'h00;      memory[36341] <=  8'h00;      memory[36342] <=  8'h00;      memory[36343] <=  8'h00;      memory[36344] <=  8'h00;      memory[36345] <=  8'h00;      memory[36346] <=  8'h00;      memory[36347] <=  8'h00;      memory[36348] <=  8'h00;      memory[36349] <=  8'h00;      memory[36350] <=  8'h00;      memory[36351] <=  8'h00;      memory[36352] <=  8'h00;      memory[36353] <=  8'h00;      memory[36354] <=  8'h00;      memory[36355] <=  8'h00;      memory[36356] <=  8'h00;      memory[36357] <=  8'h00;      memory[36358] <=  8'h00;      memory[36359] <=  8'h00;      memory[36360] <=  8'h00;      memory[36361] <=  8'h00;      memory[36362] <=  8'h00;      memory[36363] <=  8'h00;      memory[36364] <=  8'h00;      memory[36365] <=  8'h00;      memory[36366] <=  8'h00;      memory[36367] <=  8'h00;      memory[36368] <=  8'h00;      memory[36369] <=  8'h00;      memory[36370] <=  8'h00;      memory[36371] <=  8'h00;      memory[36372] <=  8'h00;      memory[36373] <=  8'h00;      memory[36374] <=  8'h00;      memory[36375] <=  8'h00;      memory[36376] <=  8'h00;      memory[36377] <=  8'h00;      memory[36378] <=  8'h00;      memory[36379] <=  8'h00;      memory[36380] <=  8'h00;      memory[36381] <=  8'h00;      memory[36382] <=  8'h00;      memory[36383] <=  8'h00;      memory[36384] <=  8'h00;      memory[36385] <=  8'h00;      memory[36386] <=  8'h00;      memory[36387] <=  8'h00;      memory[36388] <=  8'h00;      memory[36389] <=  8'h00;      memory[36390] <=  8'h00;      memory[36391] <=  8'h00;      memory[36392] <=  8'h00;      memory[36393] <=  8'h00;      memory[36394] <=  8'h00;      memory[36395] <=  8'h00;      memory[36396] <=  8'h00;      memory[36397] <=  8'h00;      memory[36398] <=  8'h00;      memory[36399] <=  8'h00;      memory[36400] <=  8'h00;      memory[36401] <=  8'h00;      memory[36402] <=  8'h00;      memory[36403] <=  8'h00;      memory[36404] <=  8'h00;      memory[36405] <=  8'h00;      memory[36406] <=  8'h00;      memory[36407] <=  8'h00;      memory[36408] <=  8'h00;      memory[36409] <=  8'h00;      memory[36410] <=  8'h00;      memory[36411] <=  8'h00;      memory[36412] <=  8'h00;      memory[36413] <=  8'h00;      memory[36414] <=  8'h00;      memory[36415] <=  8'h00;      memory[36416] <=  8'h00;      memory[36417] <=  8'h00;      memory[36418] <=  8'h00;      memory[36419] <=  8'h00;      memory[36420] <=  8'h00;      memory[36421] <=  8'h00;      memory[36422] <=  8'h00;      memory[36423] <=  8'h00;      memory[36424] <=  8'h00;      memory[36425] <=  8'h00;      memory[36426] <=  8'h00;      memory[36427] <=  8'h00;      memory[36428] <=  8'h00;      memory[36429] <=  8'h00;      memory[36430] <=  8'h00;      memory[36431] <=  8'h00;      memory[36432] <=  8'h00;      memory[36433] <=  8'h00;      memory[36434] <=  8'h00;      memory[36435] <=  8'h00;      memory[36436] <=  8'h00;      memory[36437] <=  8'h00;      memory[36438] <=  8'h00;      memory[36439] <=  8'h00;      memory[36440] <=  8'h00;      memory[36441] <=  8'h00;      memory[36442] <=  8'h00;      memory[36443] <=  8'h00;      memory[36444] <=  8'h00;      memory[36445] <=  8'h00;      memory[36446] <=  8'h00;      memory[36447] <=  8'h00;      memory[36448] <=  8'h00;      memory[36449] <=  8'h00;      memory[36450] <=  8'h00;      memory[36451] <=  8'h00;      memory[36452] <=  8'h00;      memory[36453] <=  8'h00;      memory[36454] <=  8'h00;      memory[36455] <=  8'h00;      memory[36456] <=  8'h00;      memory[36457] <=  8'h00;      memory[36458] <=  8'h00;      memory[36459] <=  8'h00;      memory[36460] <=  8'h00;      memory[36461] <=  8'h00;      memory[36462] <=  8'h00;      memory[36463] <=  8'h00;      memory[36464] <=  8'h00;      memory[36465] <=  8'h00;      memory[36466] <=  8'h00;      memory[36467] <=  8'h00;      memory[36468] <=  8'h00;      memory[36469] <=  8'h00;      memory[36470] <=  8'h00;      memory[36471] <=  8'h00;      memory[36472] <=  8'h00;      memory[36473] <=  8'h00;      memory[36474] <=  8'h00;      memory[36475] <=  8'h00;      memory[36476] <=  8'h00;      memory[36477] <=  8'h00;      memory[36478] <=  8'h00;      memory[36479] <=  8'h00;      memory[36480] <=  8'h00;      memory[36481] <=  8'h00;      memory[36482] <=  8'h00;      memory[36483] <=  8'h00;      memory[36484] <=  8'h00;      memory[36485] <=  8'h00;      memory[36486] <=  8'h00;      memory[36487] <=  8'h00;      memory[36488] <=  8'h00;      memory[36489] <=  8'h00;      memory[36490] <=  8'h00;      memory[36491] <=  8'h00;      memory[36492] <=  8'h00;      memory[36493] <=  8'h00;      memory[36494] <=  8'h00;      memory[36495] <=  8'h00;      memory[36496] <=  8'h00;      memory[36497] <=  8'h00;      memory[36498] <=  8'h00;      memory[36499] <=  8'h00;      memory[36500] <=  8'h00;      memory[36501] <=  8'h00;      memory[36502] <=  8'h00;      memory[36503] <=  8'h00;      memory[36504] <=  8'h00;      memory[36505] <=  8'h00;      memory[36506] <=  8'h00;      memory[36507] <=  8'h00;      memory[36508] <=  8'h00;      memory[36509] <=  8'h00;      memory[36510] <=  8'h00;      memory[36511] <=  8'h00;      memory[36512] <=  8'h00;      memory[36513] <=  8'h00;      memory[36514] <=  8'h00;      memory[36515] <=  8'h00;      memory[36516] <=  8'h00;      memory[36517] <=  8'h00;      memory[36518] <=  8'h00;      memory[36519] <=  8'h00;      memory[36520] <=  8'h00;      memory[36521] <=  8'h00;      memory[36522] <=  8'h00;      memory[36523] <=  8'h00;      memory[36524] <=  8'h00;      memory[36525] <=  8'h00;      memory[36526] <=  8'h00;      memory[36527] <=  8'h00;      memory[36528] <=  8'h00;      memory[36529] <=  8'h00;      memory[36530] <=  8'h00;      memory[36531] <=  8'h00;      memory[36532] <=  8'h00;      memory[36533] <=  8'h00;      memory[36534] <=  8'h00;      memory[36535] <=  8'h00;      memory[36536] <=  8'h00;      memory[36537] <=  8'h00;      memory[36538] <=  8'h00;      memory[36539] <=  8'h00;      memory[36540] <=  8'h00;      memory[36541] <=  8'h00;      memory[36542] <=  8'h00;      memory[36543] <=  8'h00;      memory[36544] <=  8'h00;      memory[36545] <=  8'h00;      memory[36546] <=  8'h00;      memory[36547] <=  8'h00;      memory[36548] <=  8'h00;      memory[36549] <=  8'h00;      memory[36550] <=  8'h00;      memory[36551] <=  8'h00;      memory[36552] <=  8'h00;      memory[36553] <=  8'h00;      memory[36554] <=  8'h00;      memory[36555] <=  8'h00;      memory[36556] <=  8'h00;      memory[36557] <=  8'h00;      memory[36558] <=  8'h00;      memory[36559] <=  8'h00;      memory[36560] <=  8'h00;      memory[36561] <=  8'h00;      memory[36562] <=  8'h00;      memory[36563] <=  8'h00;      memory[36564] <=  8'h00;      memory[36565] <=  8'h00;      memory[36566] <=  8'h00;      memory[36567] <=  8'h00;      memory[36568] <=  8'h00;      memory[36569] <=  8'h00;      memory[36570] <=  8'h00;      memory[36571] <=  8'h00;      memory[36572] <=  8'h00;      memory[36573] <=  8'h00;      memory[36574] <=  8'h00;      memory[36575] <=  8'h00;      memory[36576] <=  8'h00;      memory[36577] <=  8'h00;      memory[36578] <=  8'h00;      memory[36579] <=  8'h00;      memory[36580] <=  8'h00;      memory[36581] <=  8'h00;      memory[36582] <=  8'h00;      memory[36583] <=  8'h00;      memory[36584] <=  8'h00;      memory[36585] <=  8'h00;      memory[36586] <=  8'h00;      memory[36587] <=  8'h00;      memory[36588] <=  8'h00;      memory[36589] <=  8'h00;      memory[36590] <=  8'h00;      memory[36591] <=  8'h00;      memory[36592] <=  8'h00;      memory[36593] <=  8'h00;      memory[36594] <=  8'h00;      memory[36595] <=  8'h00;      memory[36596] <=  8'h00;      memory[36597] <=  8'h00;      memory[36598] <=  8'h00;      memory[36599] <=  8'h00;      memory[36600] <=  8'h00;      memory[36601] <=  8'h00;      memory[36602] <=  8'h00;      memory[36603] <=  8'h00;      memory[36604] <=  8'h00;      memory[36605] <=  8'h00;      memory[36606] <=  8'h00;      memory[36607] <=  8'h00;      memory[36608] <=  8'h00;      memory[36609] <=  8'h00;      memory[36610] <=  8'h00;      memory[36611] <=  8'h00;      memory[36612] <=  8'h00;      memory[36613] <=  8'h00;      memory[36614] <=  8'h00;      memory[36615] <=  8'h00;      memory[36616] <=  8'h00;      memory[36617] <=  8'h00;      memory[36618] <=  8'h00;      memory[36619] <=  8'h00;      memory[36620] <=  8'h00;      memory[36621] <=  8'h00;      memory[36622] <=  8'h00;      memory[36623] <=  8'h00;      memory[36624] <=  8'h00;      memory[36625] <=  8'h00;      memory[36626] <=  8'h00;      memory[36627] <=  8'h00;      memory[36628] <=  8'h00;      memory[36629] <=  8'h00;      memory[36630] <=  8'h00;      memory[36631] <=  8'h00;      memory[36632] <=  8'h00;      memory[36633] <=  8'h00;      memory[36634] <=  8'h00;      memory[36635] <=  8'h00;      memory[36636] <=  8'h00;      memory[36637] <=  8'h00;      memory[36638] <=  8'h00;      memory[36639] <=  8'h00;      memory[36640] <=  8'h00;      memory[36641] <=  8'h00;      memory[36642] <=  8'h00;      memory[36643] <=  8'h00;      memory[36644] <=  8'h00;      memory[36645] <=  8'h00;      memory[36646] <=  8'h00;      memory[36647] <=  8'h00;      memory[36648] <=  8'h00;      memory[36649] <=  8'h00;      memory[36650] <=  8'h00;      memory[36651] <=  8'h00;      memory[36652] <=  8'h00;      memory[36653] <=  8'h00;      memory[36654] <=  8'h00;      memory[36655] <=  8'h00;      memory[36656] <=  8'h00;      memory[36657] <=  8'h00;      memory[36658] <=  8'h00;      memory[36659] <=  8'h00;      memory[36660] <=  8'h00;      memory[36661] <=  8'h00;      memory[36662] <=  8'h00;      memory[36663] <=  8'h00;      memory[36664] <=  8'h00;      memory[36665] <=  8'h00;      memory[36666] <=  8'h00;      memory[36667] <=  8'h00;      memory[36668] <=  8'h00;      memory[36669] <=  8'h00;      memory[36670] <=  8'h00;      memory[36671] <=  8'h00;      memory[36672] <=  8'h00;      memory[36673] <=  8'h00;      memory[36674] <=  8'h00;      memory[36675] <=  8'h00;      memory[36676] <=  8'h00;      memory[36677] <=  8'h00;      memory[36678] <=  8'h00;      memory[36679] <=  8'h00;      memory[36680] <=  8'h00;      memory[36681] <=  8'h00;      memory[36682] <=  8'h00;      memory[36683] <=  8'h00;      memory[36684] <=  8'h00;      memory[36685] <=  8'h00;      memory[36686] <=  8'h00;      memory[36687] <=  8'h00;      memory[36688] <=  8'h00;      memory[36689] <=  8'h00;      memory[36690] <=  8'h00;      memory[36691] <=  8'h00;      memory[36692] <=  8'h00;      memory[36693] <=  8'h00;      memory[36694] <=  8'h00;      memory[36695] <=  8'h00;      memory[36696] <=  8'h00;      memory[36697] <=  8'h00;      memory[36698] <=  8'h00;      memory[36699] <=  8'h00;      memory[36700] <=  8'h00;      memory[36701] <=  8'h00;      memory[36702] <=  8'h00;      memory[36703] <=  8'h00;      memory[36704] <=  8'h00;      memory[36705] <=  8'h00;      memory[36706] <=  8'h00;      memory[36707] <=  8'h00;      memory[36708] <=  8'h00;      memory[36709] <=  8'h00;      memory[36710] <=  8'h00;      memory[36711] <=  8'h00;      memory[36712] <=  8'h00;      memory[36713] <=  8'h00;      memory[36714] <=  8'h00;      memory[36715] <=  8'h00;      memory[36716] <=  8'h00;      memory[36717] <=  8'h00;      memory[36718] <=  8'h00;      memory[36719] <=  8'h00;      memory[36720] <=  8'h00;      memory[36721] <=  8'h00;      memory[36722] <=  8'h00;      memory[36723] <=  8'h00;      memory[36724] <=  8'h00;      memory[36725] <=  8'h00;      memory[36726] <=  8'h00;      memory[36727] <=  8'h00;      memory[36728] <=  8'h00;      memory[36729] <=  8'h00;      memory[36730] <=  8'h00;      memory[36731] <=  8'h00;      memory[36732] <=  8'h00;      memory[36733] <=  8'h00;      memory[36734] <=  8'h00;      memory[36735] <=  8'h00;      memory[36736] <=  8'h00;      memory[36737] <=  8'h00;      memory[36738] <=  8'h00;      memory[36739] <=  8'h00;      memory[36740] <=  8'h00;      memory[36741] <=  8'h00;      memory[36742] <=  8'h00;      memory[36743] <=  8'h00;      memory[36744] <=  8'h00;      memory[36745] <=  8'h00;      memory[36746] <=  8'h00;      memory[36747] <=  8'h00;      memory[36748] <=  8'h00;      memory[36749] <=  8'h00;      memory[36750] <=  8'h00;      memory[36751] <=  8'h00;      memory[36752] <=  8'h00;      memory[36753] <=  8'h00;      memory[36754] <=  8'h00;      memory[36755] <=  8'h00;      memory[36756] <=  8'h00;      memory[36757] <=  8'h00;      memory[36758] <=  8'h00;      memory[36759] <=  8'h00;      memory[36760] <=  8'h00;      memory[36761] <=  8'h00;      memory[36762] <=  8'h00;      memory[36763] <=  8'h00;      memory[36764] <=  8'h00;      memory[36765] <=  8'h00;      memory[36766] <=  8'h00;      memory[36767] <=  8'h00;      memory[36768] <=  8'h00;      memory[36769] <=  8'h00;      memory[36770] <=  8'h00;      memory[36771] <=  8'h00;      memory[36772] <=  8'h00;      memory[36773] <=  8'h00;      memory[36774] <=  8'h00;      memory[36775] <=  8'h00;      memory[36776] <=  8'h00;      memory[36777] <=  8'h00;      memory[36778] <=  8'h00;      memory[36779] <=  8'h00;      memory[36780] <=  8'h00;      memory[36781] <=  8'h00;      memory[36782] <=  8'h00;      memory[36783] <=  8'h00;      memory[36784] <=  8'h00;      memory[36785] <=  8'h00;      memory[36786] <=  8'h00;      memory[36787] <=  8'h00;      memory[36788] <=  8'h00;      memory[36789] <=  8'h00;      memory[36790] <=  8'h00;      memory[36791] <=  8'h00;      memory[36792] <=  8'h00;      memory[36793] <=  8'h00;      memory[36794] <=  8'h00;      memory[36795] <=  8'h00;      memory[36796] <=  8'h00;      memory[36797] <=  8'h00;      memory[36798] <=  8'h00;      memory[36799] <=  8'h00;      memory[36800] <=  8'h00;      memory[36801] <=  8'h00;      memory[36802] <=  8'h00;      memory[36803] <=  8'h00;      memory[36804] <=  8'h00;      memory[36805] <=  8'h00;      memory[36806] <=  8'h00;      memory[36807] <=  8'h00;      memory[36808] <=  8'h00;      memory[36809] <=  8'h00;      memory[36810] <=  8'h00;      memory[36811] <=  8'h00;      memory[36812] <=  8'h00;      memory[36813] <=  8'h00;      memory[36814] <=  8'h00;      memory[36815] <=  8'h00;      memory[36816] <=  8'h00;      memory[36817] <=  8'h00;      memory[36818] <=  8'h00;      memory[36819] <=  8'h00;      memory[36820] <=  8'h00;      memory[36821] <=  8'h00;      memory[36822] <=  8'h00;      memory[36823] <=  8'h00;      memory[36824] <=  8'h00;      memory[36825] <=  8'h00;      memory[36826] <=  8'h00;      memory[36827] <=  8'h00;      memory[36828] <=  8'h00;      memory[36829] <=  8'h00;      memory[36830] <=  8'h00;      memory[36831] <=  8'h00;      memory[36832] <=  8'h00;      memory[36833] <=  8'h00;      memory[36834] <=  8'h00;      memory[36835] <=  8'h00;      memory[36836] <=  8'h00;      memory[36837] <=  8'h00;      memory[36838] <=  8'h00;      memory[36839] <=  8'h00;      memory[36840] <=  8'h00;      memory[36841] <=  8'h00;      memory[36842] <=  8'h00;      memory[36843] <=  8'h00;      memory[36844] <=  8'h00;      memory[36845] <=  8'h00;      memory[36846] <=  8'h00;      memory[36847] <=  8'h00;      memory[36848] <=  8'h00;      memory[36849] <=  8'h00;      memory[36850] <=  8'h00;      memory[36851] <=  8'h00;      memory[36852] <=  8'h00;      memory[36853] <=  8'h00;      memory[36854] <=  8'h00;      memory[36855] <=  8'h00;      memory[36856] <=  8'h00;      memory[36857] <=  8'h00;      memory[36858] <=  8'h00;      memory[36859] <=  8'h00;      memory[36860] <=  8'h00;      memory[36861] <=  8'h00;      memory[36862] <=  8'h00;      memory[36863] <=  8'h00;      memory[36864] <=  8'h00;      memory[36865] <=  8'h00;      memory[36866] <=  8'h00;      memory[36867] <=  8'h00;      memory[36868] <=  8'h00;      memory[36869] <=  8'h00;      memory[36870] <=  8'h00;      memory[36871] <=  8'h00;      memory[36872] <=  8'h00;      memory[36873] <=  8'h00;      memory[36874] <=  8'h00;      memory[36875] <=  8'h00;      memory[36876] <=  8'h00;      memory[36877] <=  8'h00;      memory[36878] <=  8'h00;      memory[36879] <=  8'h00;      memory[36880] <=  8'h00;      memory[36881] <=  8'h00;      memory[36882] <=  8'h00;      memory[36883] <=  8'h00;      memory[36884] <=  8'h00;      memory[36885] <=  8'h00;      memory[36886] <=  8'h00;      memory[36887] <=  8'h00;      memory[36888] <=  8'h00;      memory[36889] <=  8'h00;      memory[36890] <=  8'h00;      memory[36891] <=  8'h00;      memory[36892] <=  8'h00;      memory[36893] <=  8'h00;      memory[36894] <=  8'h00;      memory[36895] <=  8'h00;      memory[36896] <=  8'h00;      memory[36897] <=  8'h00;      memory[36898] <=  8'h00;      memory[36899] <=  8'h00;      memory[36900] <=  8'h00;      memory[36901] <=  8'h00;      memory[36902] <=  8'h00;      memory[36903] <=  8'h00;      memory[36904] <=  8'h00;      memory[36905] <=  8'h00;      memory[36906] <=  8'h00;      memory[36907] <=  8'h00;      memory[36908] <=  8'h00;      memory[36909] <=  8'h00;      memory[36910] <=  8'h00;      memory[36911] <=  8'h00;      memory[36912] <=  8'h00;      memory[36913] <=  8'h00;      memory[36914] <=  8'h00;      memory[36915] <=  8'h00;      memory[36916] <=  8'h00;      memory[36917] <=  8'h00;      memory[36918] <=  8'h00;      memory[36919] <=  8'h00;      memory[36920] <=  8'h00;      memory[36921] <=  8'h00;      memory[36922] <=  8'h00;      memory[36923] <=  8'h00;      memory[36924] <=  8'h00;      memory[36925] <=  8'h00;      memory[36926] <=  8'h00;      memory[36927] <=  8'h00;      memory[36928] <=  8'h00;      memory[36929] <=  8'h00;      memory[36930] <=  8'h00;      memory[36931] <=  8'h00;      memory[36932] <=  8'h00;      memory[36933] <=  8'h00;      memory[36934] <=  8'h00;      memory[36935] <=  8'h00;      memory[36936] <=  8'h00;      memory[36937] <=  8'h00;      memory[36938] <=  8'h00;      memory[36939] <=  8'h00;      memory[36940] <=  8'h00;      memory[36941] <=  8'h00;      memory[36942] <=  8'h00;      memory[36943] <=  8'h00;      memory[36944] <=  8'h00;      memory[36945] <=  8'h00;      memory[36946] <=  8'h00;      memory[36947] <=  8'h00;      memory[36948] <=  8'h00;      memory[36949] <=  8'h00;      memory[36950] <=  8'h00;      memory[36951] <=  8'h00;      memory[36952] <=  8'h00;      memory[36953] <=  8'h00;      memory[36954] <=  8'h00;      memory[36955] <=  8'h00;      memory[36956] <=  8'h00;      memory[36957] <=  8'h00;      memory[36958] <=  8'h00;      memory[36959] <=  8'h00;      memory[36960] <=  8'h00;      memory[36961] <=  8'h00;      memory[36962] <=  8'h00;      memory[36963] <=  8'h00;      memory[36964] <=  8'h00;      memory[36965] <=  8'h00;      memory[36966] <=  8'h00;      memory[36967] <=  8'h00;      memory[36968] <=  8'h00;      memory[36969] <=  8'h00;      memory[36970] <=  8'h00;      memory[36971] <=  8'h00;      memory[36972] <=  8'h00;      memory[36973] <=  8'h00;      memory[36974] <=  8'h00;      memory[36975] <=  8'h00;      memory[36976] <=  8'h00;      memory[36977] <=  8'h00;      memory[36978] <=  8'h00;      memory[36979] <=  8'h00;      memory[36980] <=  8'h00;      memory[36981] <=  8'h00;      memory[36982] <=  8'h00;      memory[36983] <=  8'h00;      memory[36984] <=  8'h00;      memory[36985] <=  8'h00;      memory[36986] <=  8'h00;      memory[36987] <=  8'h00;      memory[36988] <=  8'h00;      memory[36989] <=  8'h00;      memory[36990] <=  8'h00;      memory[36991] <=  8'h00;      memory[36992] <=  8'h00;      memory[36993] <=  8'h00;      memory[36994] <=  8'h00;      memory[36995] <=  8'h00;      memory[36996] <=  8'h00;      memory[36997] <=  8'h00;      memory[36998] <=  8'h00;      memory[36999] <=  8'h00;      memory[37000] <=  8'h00;      memory[37001] <=  8'h00;      memory[37002] <=  8'h00;      memory[37003] <=  8'h00;      memory[37004] <=  8'h00;      memory[37005] <=  8'h00;      memory[37006] <=  8'h00;      memory[37007] <=  8'h00;      memory[37008] <=  8'h00;      memory[37009] <=  8'h00;      memory[37010] <=  8'h00;      memory[37011] <=  8'h00;      memory[37012] <=  8'h00;      memory[37013] <=  8'h00;      memory[37014] <=  8'h00;      memory[37015] <=  8'h00;      memory[37016] <=  8'h00;      memory[37017] <=  8'h00;      memory[37018] <=  8'h00;      memory[37019] <=  8'h00;      memory[37020] <=  8'h00;      memory[37021] <=  8'h00;      memory[37022] <=  8'h00;      memory[37023] <=  8'h00;      memory[37024] <=  8'h00;      memory[37025] <=  8'h00;      memory[37026] <=  8'h00;      memory[37027] <=  8'h00;      memory[37028] <=  8'h00;      memory[37029] <=  8'h00;      memory[37030] <=  8'h00;      memory[37031] <=  8'h00;      memory[37032] <=  8'h00;      memory[37033] <=  8'h00;      memory[37034] <=  8'h00;      memory[37035] <=  8'h00;      memory[37036] <=  8'h00;      memory[37037] <=  8'h00;      memory[37038] <=  8'h00;      memory[37039] <=  8'h00;      memory[37040] <=  8'h00;      memory[37041] <=  8'h00;      memory[37042] <=  8'h00;      memory[37043] <=  8'h00;      memory[37044] <=  8'h00;      memory[37045] <=  8'h00;      memory[37046] <=  8'h00;      memory[37047] <=  8'h00;      memory[37048] <=  8'h00;      memory[37049] <=  8'h00;      memory[37050] <=  8'h00;      memory[37051] <=  8'h00;      memory[37052] <=  8'h00;      memory[37053] <=  8'h00;      memory[37054] <=  8'h00;      memory[37055] <=  8'h00;      memory[37056] <=  8'h00;      memory[37057] <=  8'h00;      memory[37058] <=  8'h00;      memory[37059] <=  8'h00;      memory[37060] <=  8'h00;      memory[37061] <=  8'h00;      memory[37062] <=  8'h00;      memory[37063] <=  8'h00;      memory[37064] <=  8'h00;      memory[37065] <=  8'h00;      memory[37066] <=  8'h00;      memory[37067] <=  8'h00;      memory[37068] <=  8'h00;      memory[37069] <=  8'h00;      memory[37070] <=  8'h00;      memory[37071] <=  8'h00;      memory[37072] <=  8'h00;      memory[37073] <=  8'h00;      memory[37074] <=  8'h00;      memory[37075] <=  8'h00;      memory[37076] <=  8'h00;      memory[37077] <=  8'h00;      memory[37078] <=  8'h00;      memory[37079] <=  8'h00;      memory[37080] <=  8'h00;      memory[37081] <=  8'h00;      memory[37082] <=  8'h00;      memory[37083] <=  8'h00;      memory[37084] <=  8'h00;      memory[37085] <=  8'h00;      memory[37086] <=  8'h00;      memory[37087] <=  8'h00;      memory[37088] <=  8'h00;      memory[37089] <=  8'h00;      memory[37090] <=  8'h00;      memory[37091] <=  8'h00;      memory[37092] <=  8'h00;      memory[37093] <=  8'h00;      memory[37094] <=  8'h00;      memory[37095] <=  8'h00;      memory[37096] <=  8'h00;      memory[37097] <=  8'h00;      memory[37098] <=  8'h00;      memory[37099] <=  8'h00;      memory[37100] <=  8'h00;      memory[37101] <=  8'h00;      memory[37102] <=  8'h00;      memory[37103] <=  8'h00;      memory[37104] <=  8'h00;      memory[37105] <=  8'h00;      memory[37106] <=  8'h00;      memory[37107] <=  8'h00;      memory[37108] <=  8'h00;      memory[37109] <=  8'h00;      memory[37110] <=  8'h00;      memory[37111] <=  8'h00;      memory[37112] <=  8'h00;      memory[37113] <=  8'h00;      memory[37114] <=  8'h00;      memory[37115] <=  8'h00;      memory[37116] <=  8'h00;      memory[37117] <=  8'h00;      memory[37118] <=  8'h00;      memory[37119] <=  8'h00;      memory[37120] <=  8'h00;      memory[37121] <=  8'h00;      memory[37122] <=  8'h00;      memory[37123] <=  8'h00;      memory[37124] <=  8'h00;      memory[37125] <=  8'h00;      memory[37126] <=  8'h00;      memory[37127] <=  8'h00;      memory[37128] <=  8'h00;      memory[37129] <=  8'h00;      memory[37130] <=  8'h00;      memory[37131] <=  8'h00;      memory[37132] <=  8'h00;      memory[37133] <=  8'h00;      memory[37134] <=  8'h00;      memory[37135] <=  8'h00;      memory[37136] <=  8'h00;      memory[37137] <=  8'h00;      memory[37138] <=  8'h00;      memory[37139] <=  8'h00;      memory[37140] <=  8'h00;      memory[37141] <=  8'h00;      memory[37142] <=  8'h00;      memory[37143] <=  8'h00;      memory[37144] <=  8'h00;      memory[37145] <=  8'h00;      memory[37146] <=  8'h00;      memory[37147] <=  8'h00;      memory[37148] <=  8'h00;      memory[37149] <=  8'h00;      memory[37150] <=  8'h00;      memory[37151] <=  8'h00;      memory[37152] <=  8'h00;      memory[37153] <=  8'h00;      memory[37154] <=  8'h00;      memory[37155] <=  8'h00;      memory[37156] <=  8'h00;      memory[37157] <=  8'h00;      memory[37158] <=  8'h00;      memory[37159] <=  8'h00;      memory[37160] <=  8'h00;      memory[37161] <=  8'h00;      memory[37162] <=  8'h00;      memory[37163] <=  8'h00;      memory[37164] <=  8'h00;      memory[37165] <=  8'h00;      memory[37166] <=  8'h00;      memory[37167] <=  8'h00;      memory[37168] <=  8'h00;      memory[37169] <=  8'h00;      memory[37170] <=  8'h00;      memory[37171] <=  8'h00;      memory[37172] <=  8'h00;      memory[37173] <=  8'h00;      memory[37174] <=  8'h00;      memory[37175] <=  8'h00;      memory[37176] <=  8'h00;      memory[37177] <=  8'h00;      memory[37178] <=  8'h00;      memory[37179] <=  8'h00;      memory[37180] <=  8'h00;      memory[37181] <=  8'h00;      memory[37182] <=  8'h00;      memory[37183] <=  8'h00;      memory[37184] <=  8'h00;      memory[37185] <=  8'h00;      memory[37186] <=  8'h00;      memory[37187] <=  8'h00;      memory[37188] <=  8'h00;      memory[37189] <=  8'h00;      memory[37190] <=  8'h00;      memory[37191] <=  8'h00;      memory[37192] <=  8'h00;      memory[37193] <=  8'h00;      memory[37194] <=  8'h00;      memory[37195] <=  8'h00;      memory[37196] <=  8'h00;      memory[37197] <=  8'h00;      memory[37198] <=  8'h00;      memory[37199] <=  8'h00;      memory[37200] <=  8'h00;      memory[37201] <=  8'h00;      memory[37202] <=  8'h00;      memory[37203] <=  8'h00;      memory[37204] <=  8'h00;      memory[37205] <=  8'h00;      memory[37206] <=  8'h00;      memory[37207] <=  8'h00;      memory[37208] <=  8'h00;      memory[37209] <=  8'h00;      memory[37210] <=  8'h00;      memory[37211] <=  8'h00;      memory[37212] <=  8'h00;      memory[37213] <=  8'h00;      memory[37214] <=  8'h00;      memory[37215] <=  8'h00;      memory[37216] <=  8'h00;      memory[37217] <=  8'h00;      memory[37218] <=  8'h00;      memory[37219] <=  8'h00;      memory[37220] <=  8'h00;      memory[37221] <=  8'h00;      memory[37222] <=  8'h00;      memory[37223] <=  8'h00;      memory[37224] <=  8'h00;      memory[37225] <=  8'h00;      memory[37226] <=  8'h00;      memory[37227] <=  8'h00;      memory[37228] <=  8'h00;      memory[37229] <=  8'h00;      memory[37230] <=  8'h00;      memory[37231] <=  8'h00;      memory[37232] <=  8'h00;      memory[37233] <=  8'h00;      memory[37234] <=  8'h00;      memory[37235] <=  8'h00;      memory[37236] <=  8'h00;      memory[37237] <=  8'h00;      memory[37238] <=  8'h00;      memory[37239] <=  8'h00;      memory[37240] <=  8'h00;      memory[37241] <=  8'h00;      memory[37242] <=  8'h00;      memory[37243] <=  8'h00;      memory[37244] <=  8'h00;      memory[37245] <=  8'h00;      memory[37246] <=  8'h00;      memory[37247] <=  8'h00;      memory[37248] <=  8'h00;      memory[37249] <=  8'h00;      memory[37250] <=  8'h00;      memory[37251] <=  8'h00;      memory[37252] <=  8'h00;      memory[37253] <=  8'h00;      memory[37254] <=  8'h00;      memory[37255] <=  8'h00;      memory[37256] <=  8'h00;      memory[37257] <=  8'h00;      memory[37258] <=  8'h00;      memory[37259] <=  8'h00;      memory[37260] <=  8'h00;      memory[37261] <=  8'h00;      memory[37262] <=  8'h00;      memory[37263] <=  8'h00;      memory[37264] <=  8'h00;      memory[37265] <=  8'h00;      memory[37266] <=  8'h00;      memory[37267] <=  8'h00;      memory[37268] <=  8'h00;      memory[37269] <=  8'h00;      memory[37270] <=  8'h00;      memory[37271] <=  8'h00;      memory[37272] <=  8'h00;      memory[37273] <=  8'h00;      memory[37274] <=  8'h00;      memory[37275] <=  8'h00;      memory[37276] <=  8'h00;      memory[37277] <=  8'h00;      memory[37278] <=  8'h00;      memory[37279] <=  8'h00;      memory[37280] <=  8'h00;      memory[37281] <=  8'h00;      memory[37282] <=  8'h00;      memory[37283] <=  8'h00;      memory[37284] <=  8'h00;      memory[37285] <=  8'h00;      memory[37286] <=  8'h00;      memory[37287] <=  8'h00;      memory[37288] <=  8'h00;      memory[37289] <=  8'h00;      memory[37290] <=  8'h00;      memory[37291] <=  8'h00;      memory[37292] <=  8'h00;      memory[37293] <=  8'h00;      memory[37294] <=  8'h00;      memory[37295] <=  8'h00;      memory[37296] <=  8'h00;      memory[37297] <=  8'h00;      memory[37298] <=  8'h00;      memory[37299] <=  8'h00;      memory[37300] <=  8'h00;      memory[37301] <=  8'h00;      memory[37302] <=  8'h00;      memory[37303] <=  8'h00;      memory[37304] <=  8'h00;      memory[37305] <=  8'h00;      memory[37306] <=  8'h00;      memory[37307] <=  8'h00;      memory[37308] <=  8'h00;      memory[37309] <=  8'h00;      memory[37310] <=  8'h00;      memory[37311] <=  8'h00;      memory[37312] <=  8'h00;      memory[37313] <=  8'h00;      memory[37314] <=  8'h00;      memory[37315] <=  8'h00;      memory[37316] <=  8'h00;      memory[37317] <=  8'h00;      memory[37318] <=  8'h00;      memory[37319] <=  8'h00;      memory[37320] <=  8'h00;      memory[37321] <=  8'h00;      memory[37322] <=  8'h00;      memory[37323] <=  8'h00;      memory[37324] <=  8'h00;      memory[37325] <=  8'h00;      memory[37326] <=  8'h00;      memory[37327] <=  8'h00;      memory[37328] <=  8'h00;      memory[37329] <=  8'h00;      memory[37330] <=  8'h00;      memory[37331] <=  8'h00;      memory[37332] <=  8'h00;      memory[37333] <=  8'h00;      memory[37334] <=  8'h00;      memory[37335] <=  8'h00;      memory[37336] <=  8'h00;      memory[37337] <=  8'h00;      memory[37338] <=  8'h00;      memory[37339] <=  8'h00;      memory[37340] <=  8'h00;      memory[37341] <=  8'h00;      memory[37342] <=  8'h00;      memory[37343] <=  8'h00;      memory[37344] <=  8'h00;      memory[37345] <=  8'h00;      memory[37346] <=  8'h00;      memory[37347] <=  8'h00;      memory[37348] <=  8'h00;      memory[37349] <=  8'h00;      memory[37350] <=  8'h00;      memory[37351] <=  8'h00;      memory[37352] <=  8'h00;      memory[37353] <=  8'h00;      memory[37354] <=  8'h00;      memory[37355] <=  8'h00;      memory[37356] <=  8'h00;      memory[37357] <=  8'h00;      memory[37358] <=  8'h00;      memory[37359] <=  8'h00;      memory[37360] <=  8'h00;      memory[37361] <=  8'h00;      memory[37362] <=  8'h00;      memory[37363] <=  8'h00;      memory[37364] <=  8'h00;      memory[37365] <=  8'h00;      memory[37366] <=  8'h00;      memory[37367] <=  8'h00;      memory[37368] <=  8'h00;      memory[37369] <=  8'h00;      memory[37370] <=  8'h00;      memory[37371] <=  8'h00;      memory[37372] <=  8'h00;      memory[37373] <=  8'h00;      memory[37374] <=  8'h00;      memory[37375] <=  8'h00;      memory[37376] <=  8'h00;      memory[37377] <=  8'h00;      memory[37378] <=  8'h00;      memory[37379] <=  8'h00;      memory[37380] <=  8'h00;      memory[37381] <=  8'h00;      memory[37382] <=  8'h00;      memory[37383] <=  8'h00;      memory[37384] <=  8'h00;      memory[37385] <=  8'h00;      memory[37386] <=  8'h00;      memory[37387] <=  8'h00;      memory[37388] <=  8'h00;      memory[37389] <=  8'h00;      memory[37390] <=  8'h00;      memory[37391] <=  8'h00;      memory[37392] <=  8'h00;      memory[37393] <=  8'h00;      memory[37394] <=  8'h00;      memory[37395] <=  8'h00;      memory[37396] <=  8'h00;      memory[37397] <=  8'h00;      memory[37398] <=  8'h00;      memory[37399] <=  8'h00;      memory[37400] <=  8'h00;      memory[37401] <=  8'h00;      memory[37402] <=  8'h00;      memory[37403] <=  8'h00;      memory[37404] <=  8'h00;      memory[37405] <=  8'h00;      memory[37406] <=  8'h00;      memory[37407] <=  8'h00;      memory[37408] <=  8'h00;      memory[37409] <=  8'h00;      memory[37410] <=  8'h00;      memory[37411] <=  8'h00;      memory[37412] <=  8'h00;      memory[37413] <=  8'h00;      memory[37414] <=  8'h00;      memory[37415] <=  8'h00;      memory[37416] <=  8'h00;      memory[37417] <=  8'h00;      memory[37418] <=  8'h00;      memory[37419] <=  8'h00;      memory[37420] <=  8'h00;      memory[37421] <=  8'h00;      memory[37422] <=  8'h00;      memory[37423] <=  8'h00;      memory[37424] <=  8'h00;      memory[37425] <=  8'h00;      memory[37426] <=  8'h00;      memory[37427] <=  8'h00;      memory[37428] <=  8'h00;      memory[37429] <=  8'h00;      memory[37430] <=  8'h00;      memory[37431] <=  8'h00;      memory[37432] <=  8'h00;      memory[37433] <=  8'h00;      memory[37434] <=  8'h00;      memory[37435] <=  8'h00;      memory[37436] <=  8'h00;      memory[37437] <=  8'h00;      memory[37438] <=  8'h00;      memory[37439] <=  8'h00;      memory[37440] <=  8'h00;      memory[37441] <=  8'h00;      memory[37442] <=  8'h00;      memory[37443] <=  8'h00;      memory[37444] <=  8'h00;      memory[37445] <=  8'h00;      memory[37446] <=  8'h00;      memory[37447] <=  8'h00;      memory[37448] <=  8'h00;      memory[37449] <=  8'h00;      memory[37450] <=  8'h00;      memory[37451] <=  8'h00;      memory[37452] <=  8'h00;      memory[37453] <=  8'h00;      memory[37454] <=  8'h00;      memory[37455] <=  8'h00;      memory[37456] <=  8'h00;      memory[37457] <=  8'h00;      memory[37458] <=  8'h00;      memory[37459] <=  8'h00;      memory[37460] <=  8'h00;      memory[37461] <=  8'h00;      memory[37462] <=  8'h00;      memory[37463] <=  8'h00;      memory[37464] <=  8'h00;      memory[37465] <=  8'h00;      memory[37466] <=  8'h00;      memory[37467] <=  8'h00;      memory[37468] <=  8'h00;      memory[37469] <=  8'h00;      memory[37470] <=  8'h00;      memory[37471] <=  8'h00;      memory[37472] <=  8'h00;      memory[37473] <=  8'h00;      memory[37474] <=  8'h00;      memory[37475] <=  8'h00;      memory[37476] <=  8'h00;      memory[37477] <=  8'h00;      memory[37478] <=  8'h00;      memory[37479] <=  8'h00;      memory[37480] <=  8'h00;      memory[37481] <=  8'h00;      memory[37482] <=  8'h00;      memory[37483] <=  8'h00;      memory[37484] <=  8'h00;      memory[37485] <=  8'h00;      memory[37486] <=  8'h00;      memory[37487] <=  8'h00;      memory[37488] <=  8'h00;      memory[37489] <=  8'h00;      memory[37490] <=  8'h00;      memory[37491] <=  8'h00;      memory[37492] <=  8'h00;      memory[37493] <=  8'h00;      memory[37494] <=  8'h00;      memory[37495] <=  8'h00;      memory[37496] <=  8'h00;      memory[37497] <=  8'h00;      memory[37498] <=  8'h00;      memory[37499] <=  8'h00;      memory[37500] <=  8'h00;      memory[37501] <=  8'h00;      memory[37502] <=  8'h00;      memory[37503] <=  8'h00;      memory[37504] <=  8'h00;      memory[37505] <=  8'h00;      memory[37506] <=  8'h00;      memory[37507] <=  8'h00;      memory[37508] <=  8'h00;      memory[37509] <=  8'h00;      memory[37510] <=  8'h00;      memory[37511] <=  8'h00;      memory[37512] <=  8'h00;      memory[37513] <=  8'h00;      memory[37514] <=  8'h00;      memory[37515] <=  8'h00;      memory[37516] <=  8'h00;      memory[37517] <=  8'h00;      memory[37518] <=  8'h00;      memory[37519] <=  8'h00;      memory[37520] <=  8'h00;      memory[37521] <=  8'h00;      memory[37522] <=  8'h00;      memory[37523] <=  8'h00;      memory[37524] <=  8'h00;      memory[37525] <=  8'h00;      memory[37526] <=  8'h00;      memory[37527] <=  8'h00;      memory[37528] <=  8'h00;      memory[37529] <=  8'h00;      memory[37530] <=  8'h00;      memory[37531] <=  8'h00;      memory[37532] <=  8'h00;      memory[37533] <=  8'h00;      memory[37534] <=  8'h00;      memory[37535] <=  8'h00;      memory[37536] <=  8'h00;      memory[37537] <=  8'h00;      memory[37538] <=  8'h00;      memory[37539] <=  8'h00;      memory[37540] <=  8'h00;      memory[37541] <=  8'h00;      memory[37542] <=  8'h00;      memory[37543] <=  8'h00;      memory[37544] <=  8'h00;      memory[37545] <=  8'h00;      memory[37546] <=  8'h00;      memory[37547] <=  8'h00;      memory[37548] <=  8'h00;      memory[37549] <=  8'h00;      memory[37550] <=  8'h00;      memory[37551] <=  8'h00;      memory[37552] <=  8'h00;      memory[37553] <=  8'h00;      memory[37554] <=  8'h00;      memory[37555] <=  8'h00;      memory[37556] <=  8'h00;      memory[37557] <=  8'h00;      memory[37558] <=  8'h00;      memory[37559] <=  8'h00;      memory[37560] <=  8'h00;      memory[37561] <=  8'h00;      memory[37562] <=  8'h00;      memory[37563] <=  8'h00;      memory[37564] <=  8'h00;      memory[37565] <=  8'h00;      memory[37566] <=  8'h00;      memory[37567] <=  8'h00;      memory[37568] <=  8'h00;      memory[37569] <=  8'h00;      memory[37570] <=  8'h00;      memory[37571] <=  8'h00;      memory[37572] <=  8'h00;      memory[37573] <=  8'h00;      memory[37574] <=  8'h00;      memory[37575] <=  8'h00;      memory[37576] <=  8'h00;      memory[37577] <=  8'h00;      memory[37578] <=  8'h00;      memory[37579] <=  8'h00;      memory[37580] <=  8'h00;      memory[37581] <=  8'h00;      memory[37582] <=  8'h00;      memory[37583] <=  8'h00;      memory[37584] <=  8'h00;      memory[37585] <=  8'h00;      memory[37586] <=  8'h00;      memory[37587] <=  8'h00;      memory[37588] <=  8'h00;      memory[37589] <=  8'h00;      memory[37590] <=  8'h00;      memory[37591] <=  8'h00;      memory[37592] <=  8'h00;      memory[37593] <=  8'h00;      memory[37594] <=  8'h00;      memory[37595] <=  8'h00;      memory[37596] <=  8'h00;      memory[37597] <=  8'h00;      memory[37598] <=  8'h00;      memory[37599] <=  8'h00;      memory[37600] <=  8'h00;      memory[37601] <=  8'h00;      memory[37602] <=  8'h00;      memory[37603] <=  8'h00;      memory[37604] <=  8'h00;      memory[37605] <=  8'h00;      memory[37606] <=  8'h00;      memory[37607] <=  8'h00;      memory[37608] <=  8'h00;      memory[37609] <=  8'h00;      memory[37610] <=  8'h00;      memory[37611] <=  8'h00;      memory[37612] <=  8'h00;      memory[37613] <=  8'h00;      memory[37614] <=  8'h00;      memory[37615] <=  8'h00;      memory[37616] <=  8'h00;      memory[37617] <=  8'h00;      memory[37618] <=  8'h00;      memory[37619] <=  8'h00;      memory[37620] <=  8'h00;      memory[37621] <=  8'h00;      memory[37622] <=  8'h00;      memory[37623] <=  8'h00;      memory[37624] <=  8'h00;      memory[37625] <=  8'h00;      memory[37626] <=  8'h00;      memory[37627] <=  8'h00;      memory[37628] <=  8'h00;      memory[37629] <=  8'h00;      memory[37630] <=  8'h00;      memory[37631] <=  8'h00;      memory[37632] <=  8'h00;      memory[37633] <=  8'h00;      memory[37634] <=  8'h00;      memory[37635] <=  8'h00;      memory[37636] <=  8'h00;      memory[37637] <=  8'h00;      memory[37638] <=  8'h00;      memory[37639] <=  8'h00;      memory[37640] <=  8'h00;      memory[37641] <=  8'h00;      memory[37642] <=  8'h00;      memory[37643] <=  8'h00;      memory[37644] <=  8'h00;      memory[37645] <=  8'h00;      memory[37646] <=  8'h00;      memory[37647] <=  8'h00;      memory[37648] <=  8'h00;      memory[37649] <=  8'h00;      memory[37650] <=  8'h00;      memory[37651] <=  8'h00;      memory[37652] <=  8'h00;      memory[37653] <=  8'h00;      memory[37654] <=  8'h00;      memory[37655] <=  8'h00;      memory[37656] <=  8'h00;      memory[37657] <=  8'h00;      memory[37658] <=  8'h00;      memory[37659] <=  8'h00;      memory[37660] <=  8'h00;      memory[37661] <=  8'h00;      memory[37662] <=  8'h00;      memory[37663] <=  8'h00;      memory[37664] <=  8'h00;      memory[37665] <=  8'h00;      memory[37666] <=  8'h00;      memory[37667] <=  8'h00;      memory[37668] <=  8'h00;      memory[37669] <=  8'h00;      memory[37670] <=  8'h00;      memory[37671] <=  8'h00;      memory[37672] <=  8'h00;      memory[37673] <=  8'h00;      memory[37674] <=  8'h00;      memory[37675] <=  8'h00;      memory[37676] <=  8'h00;      memory[37677] <=  8'h00;      memory[37678] <=  8'h00;      memory[37679] <=  8'h00;      memory[37680] <=  8'h00;      memory[37681] <=  8'h00;      memory[37682] <=  8'h00;      memory[37683] <=  8'h00;      memory[37684] <=  8'h00;      memory[37685] <=  8'h00;      memory[37686] <=  8'h00;      memory[37687] <=  8'h00;      memory[37688] <=  8'h00;      memory[37689] <=  8'h00;      memory[37690] <=  8'h00;      memory[37691] <=  8'h00;      memory[37692] <=  8'h00;      memory[37693] <=  8'h00;      memory[37694] <=  8'h00;      memory[37695] <=  8'h00;      memory[37696] <=  8'h00;      memory[37697] <=  8'h00;      memory[37698] <=  8'h00;      memory[37699] <=  8'h00;      memory[37700] <=  8'h00;      memory[37701] <=  8'h00;      memory[37702] <=  8'h00;      memory[37703] <=  8'h00;      memory[37704] <=  8'h00;      memory[37705] <=  8'h00;      memory[37706] <=  8'h00;      memory[37707] <=  8'h00;      memory[37708] <=  8'h00;      memory[37709] <=  8'h00;      memory[37710] <=  8'h00;      memory[37711] <=  8'h00;      memory[37712] <=  8'h00;      memory[37713] <=  8'h00;      memory[37714] <=  8'h00;      memory[37715] <=  8'h00;      memory[37716] <=  8'h00;      memory[37717] <=  8'h00;      memory[37718] <=  8'h00;      memory[37719] <=  8'h00;      memory[37720] <=  8'h00;      memory[37721] <=  8'h00;      memory[37722] <=  8'h00;      memory[37723] <=  8'h00;      memory[37724] <=  8'h00;      memory[37725] <=  8'h00;      memory[37726] <=  8'h00;      memory[37727] <=  8'h00;      memory[37728] <=  8'h00;      memory[37729] <=  8'h00;      memory[37730] <=  8'h00;      memory[37731] <=  8'h00;      memory[37732] <=  8'h00;      memory[37733] <=  8'h00;      memory[37734] <=  8'h00;      memory[37735] <=  8'h00;      memory[37736] <=  8'h00;      memory[37737] <=  8'h00;      memory[37738] <=  8'h00;      memory[37739] <=  8'h00;      memory[37740] <=  8'h00;      memory[37741] <=  8'h00;      memory[37742] <=  8'h00;      memory[37743] <=  8'h00;      memory[37744] <=  8'h00;      memory[37745] <=  8'h00;      memory[37746] <=  8'h00;      memory[37747] <=  8'h00;      memory[37748] <=  8'h00;      memory[37749] <=  8'h00;      memory[37750] <=  8'h00;      memory[37751] <=  8'h00;      memory[37752] <=  8'h00;      memory[37753] <=  8'h00;      memory[37754] <=  8'h00;      memory[37755] <=  8'h00;      memory[37756] <=  8'h00;      memory[37757] <=  8'h00;      memory[37758] <=  8'h00;      memory[37759] <=  8'h00;      memory[37760] <=  8'h00;      memory[37761] <=  8'h00;      memory[37762] <=  8'h00;      memory[37763] <=  8'h00;      memory[37764] <=  8'h00;      memory[37765] <=  8'h00;      memory[37766] <=  8'h00;      memory[37767] <=  8'h00;      memory[37768] <=  8'h00;      memory[37769] <=  8'h00;      memory[37770] <=  8'h00;      memory[37771] <=  8'h00;      memory[37772] <=  8'h00;      memory[37773] <=  8'h00;      memory[37774] <=  8'h00;      memory[37775] <=  8'h00;      memory[37776] <=  8'h00;      memory[37777] <=  8'h00;      memory[37778] <=  8'h00;      memory[37779] <=  8'h00;      memory[37780] <=  8'h00;      memory[37781] <=  8'h00;      memory[37782] <=  8'h00;      memory[37783] <=  8'h00;      memory[37784] <=  8'h00;      memory[37785] <=  8'h00;      memory[37786] <=  8'h00;      memory[37787] <=  8'h00;      memory[37788] <=  8'h00;      memory[37789] <=  8'h00;      memory[37790] <=  8'h00;      memory[37791] <=  8'h00;      memory[37792] <=  8'h00;      memory[37793] <=  8'h00;      memory[37794] <=  8'h00;      memory[37795] <=  8'h00;      memory[37796] <=  8'h00;      memory[37797] <=  8'h00;      memory[37798] <=  8'h00;      memory[37799] <=  8'h00;      memory[37800] <=  8'h00;      memory[37801] <=  8'h00;      memory[37802] <=  8'h00;      memory[37803] <=  8'h00;      memory[37804] <=  8'h00;      memory[37805] <=  8'h00;      memory[37806] <=  8'h00;      memory[37807] <=  8'h00;      memory[37808] <=  8'h00;      memory[37809] <=  8'h00;      memory[37810] <=  8'h00;      memory[37811] <=  8'h00;      memory[37812] <=  8'h00;      memory[37813] <=  8'h00;      memory[37814] <=  8'h00;      memory[37815] <=  8'h00;      memory[37816] <=  8'h00;      memory[37817] <=  8'h00;      memory[37818] <=  8'h00;      memory[37819] <=  8'h00;      memory[37820] <=  8'h00;      memory[37821] <=  8'h00;      memory[37822] <=  8'h00;      memory[37823] <=  8'h00;      memory[37824] <=  8'h00;      memory[37825] <=  8'h00;      memory[37826] <=  8'h00;      memory[37827] <=  8'h00;      memory[37828] <=  8'h00;      memory[37829] <=  8'h00;      memory[37830] <=  8'h00;      memory[37831] <=  8'h00;      memory[37832] <=  8'h00;      memory[37833] <=  8'h00;      memory[37834] <=  8'h00;      memory[37835] <=  8'h00;      memory[37836] <=  8'h00;      memory[37837] <=  8'h00;      memory[37838] <=  8'h00;      memory[37839] <=  8'h00;      memory[37840] <=  8'h00;      memory[37841] <=  8'h00;      memory[37842] <=  8'h00;      memory[37843] <=  8'h00;      memory[37844] <=  8'h00;      memory[37845] <=  8'h00;      memory[37846] <=  8'h00;      memory[37847] <=  8'h00;      memory[37848] <=  8'h00;      memory[37849] <=  8'h00;      memory[37850] <=  8'h00;      memory[37851] <=  8'h00;      memory[37852] <=  8'h00;      memory[37853] <=  8'h00;      memory[37854] <=  8'h00;      memory[37855] <=  8'h00;      memory[37856] <=  8'h00;      memory[37857] <=  8'h00;      memory[37858] <=  8'h00;      memory[37859] <=  8'h00;      memory[37860] <=  8'h00;      memory[37861] <=  8'h00;      memory[37862] <=  8'h00;      memory[37863] <=  8'h00;      memory[37864] <=  8'h00;      memory[37865] <=  8'h00;      memory[37866] <=  8'h00;      memory[37867] <=  8'h00;      memory[37868] <=  8'h00;      memory[37869] <=  8'h00;      memory[37870] <=  8'h00;      memory[37871] <=  8'h00;      memory[37872] <=  8'h00;      memory[37873] <=  8'h00;      memory[37874] <=  8'h00;      memory[37875] <=  8'h00;      memory[37876] <=  8'h00;      memory[37877] <=  8'h00;      memory[37878] <=  8'h00;      memory[37879] <=  8'h00;      memory[37880] <=  8'h00;      memory[37881] <=  8'h00;      memory[37882] <=  8'h00;      memory[37883] <=  8'h00;      memory[37884] <=  8'h00;      memory[37885] <=  8'h00;      memory[37886] <=  8'h00;      memory[37887] <=  8'h00;      memory[37888] <=  8'h00;      memory[37889] <=  8'h00;      memory[37890] <=  8'h00;      memory[37891] <=  8'h00;      memory[37892] <=  8'h00;      memory[37893] <=  8'h00;      memory[37894] <=  8'h00;      memory[37895] <=  8'h00;      memory[37896] <=  8'h00;      memory[37897] <=  8'h00;      memory[37898] <=  8'h00;      memory[37899] <=  8'h00;      memory[37900] <=  8'h00;      memory[37901] <=  8'h00;      memory[37902] <=  8'h00;      memory[37903] <=  8'h00;      memory[37904] <=  8'h00;      memory[37905] <=  8'h00;      memory[37906] <=  8'h00;      memory[37907] <=  8'h00;      memory[37908] <=  8'h00;      memory[37909] <=  8'h00;      memory[37910] <=  8'h00;      memory[37911] <=  8'h00;      memory[37912] <=  8'h00;      memory[37913] <=  8'h00;      memory[37914] <=  8'h00;      memory[37915] <=  8'h00;      memory[37916] <=  8'h00;      memory[37917] <=  8'h00;      memory[37918] <=  8'h00;      memory[37919] <=  8'h00;      memory[37920] <=  8'h00;      memory[37921] <=  8'h00;      memory[37922] <=  8'h00;      memory[37923] <=  8'h00;      memory[37924] <=  8'h00;      memory[37925] <=  8'h00;      memory[37926] <=  8'h00;      memory[37927] <=  8'h00;      memory[37928] <=  8'h00;      memory[37929] <=  8'h00;      memory[37930] <=  8'h00;      memory[37931] <=  8'h00;      memory[37932] <=  8'h00;      memory[37933] <=  8'h00;      memory[37934] <=  8'h00;      memory[37935] <=  8'h00;      memory[37936] <=  8'h00;      memory[37937] <=  8'h00;      memory[37938] <=  8'h00;      memory[37939] <=  8'h00;      memory[37940] <=  8'h00;      memory[37941] <=  8'h00;      memory[37942] <=  8'h00;      memory[37943] <=  8'h00;      memory[37944] <=  8'h00;      memory[37945] <=  8'h00;      memory[37946] <=  8'h00;      memory[37947] <=  8'h00;      memory[37948] <=  8'h00;      memory[37949] <=  8'h00;      memory[37950] <=  8'h00;      memory[37951] <=  8'h00;      memory[37952] <=  8'h00;      memory[37953] <=  8'h00;      memory[37954] <=  8'h00;      memory[37955] <=  8'h00;      memory[37956] <=  8'h00;      memory[37957] <=  8'h00;      memory[37958] <=  8'h00;      memory[37959] <=  8'h00;      memory[37960] <=  8'h00;      memory[37961] <=  8'h00;      memory[37962] <=  8'h00;      memory[37963] <=  8'h00;      memory[37964] <=  8'h00;      memory[37965] <=  8'h00;      memory[37966] <=  8'h00;      memory[37967] <=  8'h00;      memory[37968] <=  8'h00;      memory[37969] <=  8'h00;      memory[37970] <=  8'h00;      memory[37971] <=  8'h00;      memory[37972] <=  8'h00;      memory[37973] <=  8'h00;      memory[37974] <=  8'h00;      memory[37975] <=  8'h00;      memory[37976] <=  8'h00;      memory[37977] <=  8'h00;      memory[37978] <=  8'h00;      memory[37979] <=  8'h00;      memory[37980] <=  8'h00;      memory[37981] <=  8'h00;      memory[37982] <=  8'h00;      memory[37983] <=  8'h00;      memory[37984] <=  8'h00;      memory[37985] <=  8'h00;      memory[37986] <=  8'h00;      memory[37987] <=  8'h00;      memory[37988] <=  8'h00;      memory[37989] <=  8'h00;      memory[37990] <=  8'h00;      memory[37991] <=  8'h00;      memory[37992] <=  8'h00;      memory[37993] <=  8'h00;      memory[37994] <=  8'h00;      memory[37995] <=  8'h00;      memory[37996] <=  8'h00;      memory[37997] <=  8'h00;      memory[37998] <=  8'h00;      memory[37999] <=  8'h00;      memory[38000] <=  8'h00;      memory[38001] <=  8'h00;      memory[38002] <=  8'h00;      memory[38003] <=  8'h00;      memory[38004] <=  8'h00;      memory[38005] <=  8'h00;      memory[38006] <=  8'h00;      memory[38007] <=  8'h00;      memory[38008] <=  8'h00;      memory[38009] <=  8'h00;      memory[38010] <=  8'h00;      memory[38011] <=  8'h00;      memory[38012] <=  8'h00;      memory[38013] <=  8'h00;      memory[38014] <=  8'h00;      memory[38015] <=  8'h00;      memory[38016] <=  8'h00;      memory[38017] <=  8'h00;      memory[38018] <=  8'h00;      memory[38019] <=  8'h00;      memory[38020] <=  8'h00;      memory[38021] <=  8'h00;      memory[38022] <=  8'h00;      memory[38023] <=  8'h00;      memory[38024] <=  8'h00;      memory[38025] <=  8'h00;      memory[38026] <=  8'h00;      memory[38027] <=  8'h00;      memory[38028] <=  8'h00;      memory[38029] <=  8'h00;      memory[38030] <=  8'h00;      memory[38031] <=  8'h00;      memory[38032] <=  8'h00;      memory[38033] <=  8'h00;      memory[38034] <=  8'h00;      memory[38035] <=  8'h00;      memory[38036] <=  8'h00;      memory[38037] <=  8'h00;      memory[38038] <=  8'h00;      memory[38039] <=  8'h00;      memory[38040] <=  8'h00;      memory[38041] <=  8'h00;      memory[38042] <=  8'h00;      memory[38043] <=  8'h00;      memory[38044] <=  8'h00;      memory[38045] <=  8'h00;      memory[38046] <=  8'h00;      memory[38047] <=  8'h00;      memory[38048] <=  8'h00;      memory[38049] <=  8'h00;      memory[38050] <=  8'h00;      memory[38051] <=  8'h00;      memory[38052] <=  8'h00;      memory[38053] <=  8'h00;      memory[38054] <=  8'h00;      memory[38055] <=  8'h00;      memory[38056] <=  8'h00;      memory[38057] <=  8'h00;      memory[38058] <=  8'h00;      memory[38059] <=  8'h00;      memory[38060] <=  8'h00;      memory[38061] <=  8'h00;      memory[38062] <=  8'h00;      memory[38063] <=  8'h00;      memory[38064] <=  8'h00;      memory[38065] <=  8'h00;      memory[38066] <=  8'h00;      memory[38067] <=  8'h00;      memory[38068] <=  8'h00;      memory[38069] <=  8'h00;      memory[38070] <=  8'h00;      memory[38071] <=  8'h00;      memory[38072] <=  8'h00;      memory[38073] <=  8'h00;      memory[38074] <=  8'h00;      memory[38075] <=  8'h00;      memory[38076] <=  8'h00;      memory[38077] <=  8'h00;      memory[38078] <=  8'h00;      memory[38079] <=  8'h00;      memory[38080] <=  8'h00;      memory[38081] <=  8'h00;      memory[38082] <=  8'h00;      memory[38083] <=  8'h00;      memory[38084] <=  8'h00;      memory[38085] <=  8'h00;      memory[38086] <=  8'h00;      memory[38087] <=  8'h00;      memory[38088] <=  8'h00;      memory[38089] <=  8'h00;      memory[38090] <=  8'h00;      memory[38091] <=  8'h00;      memory[38092] <=  8'h00;      memory[38093] <=  8'h00;      memory[38094] <=  8'h00;      memory[38095] <=  8'h00;      memory[38096] <=  8'h00;      memory[38097] <=  8'h00;      memory[38098] <=  8'h00;      memory[38099] <=  8'h00;      memory[38100] <=  8'h00;      memory[38101] <=  8'h00;      memory[38102] <=  8'h00;      memory[38103] <=  8'h00;      memory[38104] <=  8'h00;      memory[38105] <=  8'h00;      memory[38106] <=  8'h00;      memory[38107] <=  8'h00;      memory[38108] <=  8'h00;      memory[38109] <=  8'h00;      memory[38110] <=  8'h00;      memory[38111] <=  8'h00;      memory[38112] <=  8'h00;      memory[38113] <=  8'h00;      memory[38114] <=  8'h00;      memory[38115] <=  8'h00;      memory[38116] <=  8'h00;      memory[38117] <=  8'h00;      memory[38118] <=  8'h00;      memory[38119] <=  8'h00;      memory[38120] <=  8'h00;      memory[38121] <=  8'h00;      memory[38122] <=  8'h00;      memory[38123] <=  8'h00;      memory[38124] <=  8'h00;      memory[38125] <=  8'h00;      memory[38126] <=  8'h00;      memory[38127] <=  8'h00;      memory[38128] <=  8'h00;      memory[38129] <=  8'h00;      memory[38130] <=  8'h00;      memory[38131] <=  8'h00;      memory[38132] <=  8'h00;      memory[38133] <=  8'h00;      memory[38134] <=  8'h00;      memory[38135] <=  8'h00;      memory[38136] <=  8'h00;      memory[38137] <=  8'h00;      memory[38138] <=  8'h00;      memory[38139] <=  8'h00;      memory[38140] <=  8'h00;      memory[38141] <=  8'h00;      memory[38142] <=  8'h00;      memory[38143] <=  8'h00;      memory[38144] <=  8'h00;      memory[38145] <=  8'h00;      memory[38146] <=  8'h00;      memory[38147] <=  8'h00;      memory[38148] <=  8'h00;      memory[38149] <=  8'h00;      memory[38150] <=  8'h00;      memory[38151] <=  8'h00;      memory[38152] <=  8'h00;      memory[38153] <=  8'h00;      memory[38154] <=  8'h00;      memory[38155] <=  8'h00;      memory[38156] <=  8'h00;      memory[38157] <=  8'h00;      memory[38158] <=  8'h00;      memory[38159] <=  8'h00;      memory[38160] <=  8'h00;      memory[38161] <=  8'h00;      memory[38162] <=  8'h00;      memory[38163] <=  8'h00;      memory[38164] <=  8'h00;      memory[38165] <=  8'h00;      memory[38166] <=  8'h00;      memory[38167] <=  8'h00;      memory[38168] <=  8'h00;      memory[38169] <=  8'h00;      memory[38170] <=  8'h00;      memory[38171] <=  8'h00;      memory[38172] <=  8'h00;      memory[38173] <=  8'h00;      memory[38174] <=  8'h00;      memory[38175] <=  8'h00;      memory[38176] <=  8'h00;      memory[38177] <=  8'h00;      memory[38178] <=  8'h00;      memory[38179] <=  8'h00;      memory[38180] <=  8'h00;      memory[38181] <=  8'h00;      memory[38182] <=  8'h00;      memory[38183] <=  8'h00;      memory[38184] <=  8'h00;      memory[38185] <=  8'h00;      memory[38186] <=  8'h00;      memory[38187] <=  8'h00;      memory[38188] <=  8'h00;      memory[38189] <=  8'h00;      memory[38190] <=  8'h00;      memory[38191] <=  8'h00;      memory[38192] <=  8'h00;      memory[38193] <=  8'h00;      memory[38194] <=  8'h00;      memory[38195] <=  8'h00;      memory[38196] <=  8'h00;      memory[38197] <=  8'h00;      memory[38198] <=  8'h00;      memory[38199] <=  8'h00;      memory[38200] <=  8'h00;      memory[38201] <=  8'h00;      memory[38202] <=  8'h00;      memory[38203] <=  8'h00;      memory[38204] <=  8'h00;      memory[38205] <=  8'h00;      memory[38206] <=  8'h00;      memory[38207] <=  8'h00;      memory[38208] <=  8'h00;      memory[38209] <=  8'h00;      memory[38210] <=  8'h00;      memory[38211] <=  8'h00;      memory[38212] <=  8'h00;      memory[38213] <=  8'h00;      memory[38214] <=  8'h00;      memory[38215] <=  8'h00;      memory[38216] <=  8'h00;      memory[38217] <=  8'h00;      memory[38218] <=  8'h00;      memory[38219] <=  8'h00;      memory[38220] <=  8'h00;      memory[38221] <=  8'h00;      memory[38222] <=  8'h00;      memory[38223] <=  8'h00;      memory[38224] <=  8'h00;      memory[38225] <=  8'h00;      memory[38226] <=  8'h00;      memory[38227] <=  8'h00;      memory[38228] <=  8'h00;      memory[38229] <=  8'h00;      memory[38230] <=  8'h00;      memory[38231] <=  8'h00;      memory[38232] <=  8'h00;      memory[38233] <=  8'h00;      memory[38234] <=  8'h00;      memory[38235] <=  8'h00;      memory[38236] <=  8'h00;      memory[38237] <=  8'h00;      memory[38238] <=  8'h00;      memory[38239] <=  8'h00;      memory[38240] <=  8'h00;      memory[38241] <=  8'h00;      memory[38242] <=  8'h00;      memory[38243] <=  8'h00;      memory[38244] <=  8'h00;      memory[38245] <=  8'h00;      memory[38246] <=  8'h00;      memory[38247] <=  8'h00;      memory[38248] <=  8'h00;      memory[38249] <=  8'h00;      memory[38250] <=  8'h00;      memory[38251] <=  8'h00;      memory[38252] <=  8'h00;      memory[38253] <=  8'h00;      memory[38254] <=  8'h00;      memory[38255] <=  8'h00;      memory[38256] <=  8'h00;      memory[38257] <=  8'h00;      memory[38258] <=  8'h00;      memory[38259] <=  8'h00;      memory[38260] <=  8'h00;      memory[38261] <=  8'h00;      memory[38262] <=  8'h00;      memory[38263] <=  8'h00;      memory[38264] <=  8'h00;      memory[38265] <=  8'h00;      memory[38266] <=  8'h00;      memory[38267] <=  8'h00;      memory[38268] <=  8'h00;      memory[38269] <=  8'h00;      memory[38270] <=  8'h00;      memory[38271] <=  8'h00;      memory[38272] <=  8'h00;      memory[38273] <=  8'h00;      memory[38274] <=  8'h00;      memory[38275] <=  8'h00;      memory[38276] <=  8'h00;      memory[38277] <=  8'h00;      memory[38278] <=  8'h00;      memory[38279] <=  8'h00;      memory[38280] <=  8'h00;      memory[38281] <=  8'h00;      memory[38282] <=  8'h00;      memory[38283] <=  8'h00;      memory[38284] <=  8'h00;      memory[38285] <=  8'h00;      memory[38286] <=  8'h00;      memory[38287] <=  8'h00;      memory[38288] <=  8'h00;      memory[38289] <=  8'h00;      memory[38290] <=  8'h00;      memory[38291] <=  8'h00;      memory[38292] <=  8'h00;      memory[38293] <=  8'h00;      memory[38294] <=  8'h00;      memory[38295] <=  8'h00;      memory[38296] <=  8'h00;      memory[38297] <=  8'h00;      memory[38298] <=  8'h00;      memory[38299] <=  8'h00;      memory[38300] <=  8'h00;      memory[38301] <=  8'h00;      memory[38302] <=  8'h00;      memory[38303] <=  8'h00;      memory[38304] <=  8'h00;      memory[38305] <=  8'h00;      memory[38306] <=  8'h00;      memory[38307] <=  8'h00;      memory[38308] <=  8'h00;      memory[38309] <=  8'h00;      memory[38310] <=  8'h00;      memory[38311] <=  8'h00;      memory[38312] <=  8'h00;      memory[38313] <=  8'h00;      memory[38314] <=  8'h00;      memory[38315] <=  8'h00;      memory[38316] <=  8'h00;      memory[38317] <=  8'h00;      memory[38318] <=  8'h00;      memory[38319] <=  8'h00;      memory[38320] <=  8'h00;      memory[38321] <=  8'h00;      memory[38322] <=  8'h00;      memory[38323] <=  8'h00;      memory[38324] <=  8'h00;      memory[38325] <=  8'h00;      memory[38326] <=  8'h00;      memory[38327] <=  8'h00;      memory[38328] <=  8'h00;      memory[38329] <=  8'h00;      memory[38330] <=  8'h00;      memory[38331] <=  8'h00;      memory[38332] <=  8'h00;      memory[38333] <=  8'h00;      memory[38334] <=  8'h00;      memory[38335] <=  8'h00;      memory[38336] <=  8'h00;      memory[38337] <=  8'h00;      memory[38338] <=  8'h00;      memory[38339] <=  8'h00;      memory[38340] <=  8'h00;      memory[38341] <=  8'h00;      memory[38342] <=  8'h00;      memory[38343] <=  8'h00;      memory[38344] <=  8'h00;      memory[38345] <=  8'h00;      memory[38346] <=  8'h00;      memory[38347] <=  8'h00;      memory[38348] <=  8'h00;      memory[38349] <=  8'h00;      memory[38350] <=  8'h00;      memory[38351] <=  8'h00;      memory[38352] <=  8'h00;      memory[38353] <=  8'h00;      memory[38354] <=  8'h00;      memory[38355] <=  8'h00;      memory[38356] <=  8'h00;      memory[38357] <=  8'h00;      memory[38358] <=  8'h00;      memory[38359] <=  8'h00;      memory[38360] <=  8'h00;      memory[38361] <=  8'h00;      memory[38362] <=  8'h00;      memory[38363] <=  8'h00;      memory[38364] <=  8'h00;      memory[38365] <=  8'h00;      memory[38366] <=  8'h00;      memory[38367] <=  8'h00;      memory[38368] <=  8'h00;      memory[38369] <=  8'h00;      memory[38370] <=  8'h00;      memory[38371] <=  8'h00;      memory[38372] <=  8'h00;      memory[38373] <=  8'h00;      memory[38374] <=  8'h00;      memory[38375] <=  8'h00;      memory[38376] <=  8'h00;      memory[38377] <=  8'h00;      memory[38378] <=  8'h00;      memory[38379] <=  8'h00;      memory[38380] <=  8'h00;      memory[38381] <=  8'h00;      memory[38382] <=  8'h00;      memory[38383] <=  8'h00;      memory[38384] <=  8'h00;      memory[38385] <=  8'h00;      memory[38386] <=  8'h00;      memory[38387] <=  8'h00;      memory[38388] <=  8'h00;      memory[38389] <=  8'h00;      memory[38390] <=  8'h00;      memory[38391] <=  8'h00;      memory[38392] <=  8'h00;      memory[38393] <=  8'h00;      memory[38394] <=  8'h00;      memory[38395] <=  8'h00;      memory[38396] <=  8'h00;      memory[38397] <=  8'h00;      memory[38398] <=  8'h00;      memory[38399] <=  8'h00;      memory[38400] <=  8'h00;      memory[38401] <=  8'h00;      memory[38402] <=  8'h00;      memory[38403] <=  8'h00;      memory[38404] <=  8'h00;      memory[38405] <=  8'h00;      memory[38406] <=  8'h00;      memory[38407] <=  8'h00;      memory[38408] <=  8'h00;      memory[38409] <=  8'h00;      memory[38410] <=  8'h00;      memory[38411] <=  8'h00;      memory[38412] <=  8'h00;      memory[38413] <=  8'h00;      memory[38414] <=  8'h00;      memory[38415] <=  8'h00;      memory[38416] <=  8'h00;      memory[38417] <=  8'h00;      memory[38418] <=  8'h00;      memory[38419] <=  8'h00;      memory[38420] <=  8'h00;      memory[38421] <=  8'h00;      memory[38422] <=  8'h00;      memory[38423] <=  8'h00;      memory[38424] <=  8'h00;      memory[38425] <=  8'h00;      memory[38426] <=  8'h00;      memory[38427] <=  8'h00;      memory[38428] <=  8'h00;      memory[38429] <=  8'h00;      memory[38430] <=  8'h00;      memory[38431] <=  8'h00;      memory[38432] <=  8'h00;      memory[38433] <=  8'h00;      memory[38434] <=  8'h00;      memory[38435] <=  8'h00;      memory[38436] <=  8'h00;      memory[38437] <=  8'h00;      memory[38438] <=  8'h00;      memory[38439] <=  8'h00;      memory[38440] <=  8'h00;      memory[38441] <=  8'h00;      memory[38442] <=  8'h00;      memory[38443] <=  8'h00;      memory[38444] <=  8'h00;      memory[38445] <=  8'h00;      memory[38446] <=  8'h00;      memory[38447] <=  8'h00;      memory[38448] <=  8'h00;      memory[38449] <=  8'h00;      memory[38450] <=  8'h00;      memory[38451] <=  8'h00;      memory[38452] <=  8'h00;      memory[38453] <=  8'h00;      memory[38454] <=  8'h00;      memory[38455] <=  8'h00;      memory[38456] <=  8'h00;      memory[38457] <=  8'h00;      memory[38458] <=  8'h00;      memory[38459] <=  8'h00;      memory[38460] <=  8'h00;      memory[38461] <=  8'h00;      memory[38462] <=  8'h00;      memory[38463] <=  8'h00;      memory[38464] <=  8'h00;      memory[38465] <=  8'h00;      memory[38466] <=  8'h00;      memory[38467] <=  8'h00;      memory[38468] <=  8'h00;      memory[38469] <=  8'h00;      memory[38470] <=  8'h00;      memory[38471] <=  8'h00;      memory[38472] <=  8'h00;      memory[38473] <=  8'h00;      memory[38474] <=  8'h00;      memory[38475] <=  8'h00;      memory[38476] <=  8'h00;      memory[38477] <=  8'h00;      memory[38478] <=  8'h00;      memory[38479] <=  8'h00;      memory[38480] <=  8'h00;      memory[38481] <=  8'h00;      memory[38482] <=  8'h00;      memory[38483] <=  8'h00;      memory[38484] <=  8'h00;      memory[38485] <=  8'h00;      memory[38486] <=  8'h00;      memory[38487] <=  8'h00;      memory[38488] <=  8'h00;      memory[38489] <=  8'h00;      memory[38490] <=  8'h00;      memory[38491] <=  8'h00;      memory[38492] <=  8'h00;      memory[38493] <=  8'h00;      memory[38494] <=  8'h00;      memory[38495] <=  8'h00;      memory[38496] <=  8'h00;      memory[38497] <=  8'h00;      memory[38498] <=  8'h00;      memory[38499] <=  8'h00;      memory[38500] <=  8'h00;      memory[38501] <=  8'h00;      memory[38502] <=  8'h00;      memory[38503] <=  8'h00;      memory[38504] <=  8'h00;      memory[38505] <=  8'h00;      memory[38506] <=  8'h00;      memory[38507] <=  8'h00;      memory[38508] <=  8'h00;      memory[38509] <=  8'h00;      memory[38510] <=  8'h00;      memory[38511] <=  8'h00;      memory[38512] <=  8'h00;      memory[38513] <=  8'h00;      memory[38514] <=  8'h00;      memory[38515] <=  8'h00;      memory[38516] <=  8'h00;      memory[38517] <=  8'h00;      memory[38518] <=  8'h00;      memory[38519] <=  8'h00;      memory[38520] <=  8'h00;      memory[38521] <=  8'h00;      memory[38522] <=  8'h00;      memory[38523] <=  8'h00;      memory[38524] <=  8'h00;      memory[38525] <=  8'h00;      memory[38526] <=  8'h00;      memory[38527] <=  8'h00;      memory[38528] <=  8'h00;      memory[38529] <=  8'h00;      memory[38530] <=  8'h00;      memory[38531] <=  8'h00;      memory[38532] <=  8'h00;      memory[38533] <=  8'h00;      memory[38534] <=  8'h00;      memory[38535] <=  8'h00;      memory[38536] <=  8'h00;      memory[38537] <=  8'h00;      memory[38538] <=  8'h00;      memory[38539] <=  8'h00;      memory[38540] <=  8'h00;      memory[38541] <=  8'h00;      memory[38542] <=  8'h00;      memory[38543] <=  8'h00;      memory[38544] <=  8'h00;      memory[38545] <=  8'h00;      memory[38546] <=  8'h00;      memory[38547] <=  8'h00;      memory[38548] <=  8'h00;      memory[38549] <=  8'h00;      memory[38550] <=  8'h00;      memory[38551] <=  8'h00;      memory[38552] <=  8'h00;      memory[38553] <=  8'h00;      memory[38554] <=  8'h00;      memory[38555] <=  8'h00;      memory[38556] <=  8'h00;      memory[38557] <=  8'h00;      memory[38558] <=  8'h00;      memory[38559] <=  8'h00;      memory[38560] <=  8'h00;      memory[38561] <=  8'h00;      memory[38562] <=  8'h00;      memory[38563] <=  8'h00;      memory[38564] <=  8'h00;      memory[38565] <=  8'h00;      memory[38566] <=  8'h00;      memory[38567] <=  8'h00;      memory[38568] <=  8'h00;      memory[38569] <=  8'h00;      memory[38570] <=  8'h00;      memory[38571] <=  8'h00;      memory[38572] <=  8'h00;      memory[38573] <=  8'h00;      memory[38574] <=  8'h00;      memory[38575] <=  8'h00;      memory[38576] <=  8'h00;      memory[38577] <=  8'h00;      memory[38578] <=  8'h00;      memory[38579] <=  8'h00;      memory[38580] <=  8'h00;      memory[38581] <=  8'h00;      memory[38582] <=  8'h00;      memory[38583] <=  8'h00;      memory[38584] <=  8'h00;      memory[38585] <=  8'h00;      memory[38586] <=  8'h00;      memory[38587] <=  8'h00;      memory[38588] <=  8'h00;      memory[38589] <=  8'h00;      memory[38590] <=  8'h00;      memory[38591] <=  8'h00;      memory[38592] <=  8'h00;      memory[38593] <=  8'h00;      memory[38594] <=  8'h00;      memory[38595] <=  8'h00;      memory[38596] <=  8'h00;      memory[38597] <=  8'h00;      memory[38598] <=  8'h00;      memory[38599] <=  8'h00;      memory[38600] <=  8'h00;      memory[38601] <=  8'h00;      memory[38602] <=  8'h00;      memory[38603] <=  8'h00;      memory[38604] <=  8'h00;      memory[38605] <=  8'h00;      memory[38606] <=  8'h00;      memory[38607] <=  8'h00;      memory[38608] <=  8'h00;      memory[38609] <=  8'h00;      memory[38610] <=  8'h00;      memory[38611] <=  8'h00;      memory[38612] <=  8'h00;      memory[38613] <=  8'h00;      memory[38614] <=  8'h00;      memory[38615] <=  8'h00;      memory[38616] <=  8'h00;      memory[38617] <=  8'h00;      memory[38618] <=  8'h00;      memory[38619] <=  8'h00;      memory[38620] <=  8'h00;      memory[38621] <=  8'h00;      memory[38622] <=  8'h00;      memory[38623] <=  8'h00;      memory[38624] <=  8'h00;      memory[38625] <=  8'h00;      memory[38626] <=  8'h00;      memory[38627] <=  8'h00;      memory[38628] <=  8'h00;      memory[38629] <=  8'h00;      memory[38630] <=  8'h00;      memory[38631] <=  8'h00;      memory[38632] <=  8'h00;      memory[38633] <=  8'h00;      memory[38634] <=  8'h00;      memory[38635] <=  8'h00;      memory[38636] <=  8'h00;      memory[38637] <=  8'h00;      memory[38638] <=  8'h00;      memory[38639] <=  8'h00;      memory[38640] <=  8'h00;      memory[38641] <=  8'h00;      memory[38642] <=  8'h00;      memory[38643] <=  8'h00;      memory[38644] <=  8'h00;      memory[38645] <=  8'h00;      memory[38646] <=  8'h00;      memory[38647] <=  8'h00;      memory[38648] <=  8'h00;      memory[38649] <=  8'h00;      memory[38650] <=  8'h00;      memory[38651] <=  8'h00;      memory[38652] <=  8'h00;      memory[38653] <=  8'h00;      memory[38654] <=  8'h00;      memory[38655] <=  8'h00;      memory[38656] <=  8'h00;      memory[38657] <=  8'h00;      memory[38658] <=  8'h00;      memory[38659] <=  8'h00;      memory[38660] <=  8'h00;      memory[38661] <=  8'h00;      memory[38662] <=  8'h00;      memory[38663] <=  8'h00;      memory[38664] <=  8'h00;      memory[38665] <=  8'h00;      memory[38666] <=  8'h00;      memory[38667] <=  8'h00;      memory[38668] <=  8'h00;      memory[38669] <=  8'h00;      memory[38670] <=  8'h00;      memory[38671] <=  8'h00;      memory[38672] <=  8'h00;      memory[38673] <=  8'h00;      memory[38674] <=  8'h00;      memory[38675] <=  8'h00;      memory[38676] <=  8'h00;      memory[38677] <=  8'h00;      memory[38678] <=  8'h00;      memory[38679] <=  8'h00;      memory[38680] <=  8'h00;      memory[38681] <=  8'h00;      memory[38682] <=  8'h00;      memory[38683] <=  8'h00;      memory[38684] <=  8'h00;      memory[38685] <=  8'h00;      memory[38686] <=  8'h00;      memory[38687] <=  8'h00;      memory[38688] <=  8'h00;      memory[38689] <=  8'h00;      memory[38690] <=  8'h00;      memory[38691] <=  8'h00;      memory[38692] <=  8'h00;      memory[38693] <=  8'h00;      memory[38694] <=  8'h00;      memory[38695] <=  8'h00;      memory[38696] <=  8'h00;      memory[38697] <=  8'h00;      memory[38698] <=  8'h00;      memory[38699] <=  8'h00;      memory[38700] <=  8'h00;      memory[38701] <=  8'h00;      memory[38702] <=  8'h00;      memory[38703] <=  8'h00;      memory[38704] <=  8'h00;      memory[38705] <=  8'h00;      memory[38706] <=  8'h00;      memory[38707] <=  8'h00;      memory[38708] <=  8'h00;      memory[38709] <=  8'h00;      memory[38710] <=  8'h00;      memory[38711] <=  8'h00;      memory[38712] <=  8'h00;      memory[38713] <=  8'h00;      memory[38714] <=  8'h00;      memory[38715] <=  8'h00;      memory[38716] <=  8'h00;      memory[38717] <=  8'h00;      memory[38718] <=  8'h00;      memory[38719] <=  8'h00;      memory[38720] <=  8'h00;      memory[38721] <=  8'h00;      memory[38722] <=  8'h00;      memory[38723] <=  8'h00;      memory[38724] <=  8'h00;      memory[38725] <=  8'h00;      memory[38726] <=  8'h00;      memory[38727] <=  8'h00;      memory[38728] <=  8'h00;      memory[38729] <=  8'h00;      memory[38730] <=  8'h00;      memory[38731] <=  8'h00;      memory[38732] <=  8'h00;      memory[38733] <=  8'h00;      memory[38734] <=  8'h00;      memory[38735] <=  8'h00;      memory[38736] <=  8'h00;      memory[38737] <=  8'h00;      memory[38738] <=  8'h00;      memory[38739] <=  8'h00;      memory[38740] <=  8'h00;      memory[38741] <=  8'h00;      memory[38742] <=  8'h00;      memory[38743] <=  8'h00;      memory[38744] <=  8'h00;      memory[38745] <=  8'h00;      memory[38746] <=  8'h00;      memory[38747] <=  8'h00;      memory[38748] <=  8'h00;      memory[38749] <=  8'h00;      memory[38750] <=  8'h00;      memory[38751] <=  8'h00;      memory[38752] <=  8'h00;      memory[38753] <=  8'h00;      memory[38754] <=  8'h00;      memory[38755] <=  8'h00;      memory[38756] <=  8'h00;      memory[38757] <=  8'h00;      memory[38758] <=  8'h00;      memory[38759] <=  8'h00;      memory[38760] <=  8'h00;      memory[38761] <=  8'h00;      memory[38762] <=  8'h00;      memory[38763] <=  8'h00;      memory[38764] <=  8'h00;      memory[38765] <=  8'h00;      memory[38766] <=  8'h00;      memory[38767] <=  8'h00;      memory[38768] <=  8'h00;      memory[38769] <=  8'h00;      memory[38770] <=  8'h00;      memory[38771] <=  8'h00;      memory[38772] <=  8'h00;      memory[38773] <=  8'h00;      memory[38774] <=  8'h00;      memory[38775] <=  8'h00;      memory[38776] <=  8'h00;      memory[38777] <=  8'h00;      memory[38778] <=  8'h00;      memory[38779] <=  8'h00;      memory[38780] <=  8'h00;      memory[38781] <=  8'h00;      memory[38782] <=  8'h00;      memory[38783] <=  8'h00;      memory[38784] <=  8'h00;      memory[38785] <=  8'h00;      memory[38786] <=  8'h00;      memory[38787] <=  8'h00;      memory[38788] <=  8'h00;      memory[38789] <=  8'h00;      memory[38790] <=  8'h00;      memory[38791] <=  8'h00;      memory[38792] <=  8'h00;      memory[38793] <=  8'h00;      memory[38794] <=  8'h00;      memory[38795] <=  8'h00;      memory[38796] <=  8'h00;      memory[38797] <=  8'h00;      memory[38798] <=  8'h00;      memory[38799] <=  8'h00;      memory[38800] <=  8'h00;      memory[38801] <=  8'h00;      memory[38802] <=  8'h00;      memory[38803] <=  8'h00;      memory[38804] <=  8'h00;      memory[38805] <=  8'h00;      memory[38806] <=  8'h00;      memory[38807] <=  8'h00;      memory[38808] <=  8'h00;      memory[38809] <=  8'h00;      memory[38810] <=  8'h00;      memory[38811] <=  8'h00;      memory[38812] <=  8'h00;      memory[38813] <=  8'h00;      memory[38814] <=  8'h00;      memory[38815] <=  8'h00;      memory[38816] <=  8'h00;      memory[38817] <=  8'h00;      memory[38818] <=  8'h00;      memory[38819] <=  8'h00;      memory[38820] <=  8'h00;      memory[38821] <=  8'h00;      memory[38822] <=  8'h00;      memory[38823] <=  8'h00;      memory[38824] <=  8'h00;      memory[38825] <=  8'h00;      memory[38826] <=  8'h00;      memory[38827] <=  8'h00;      memory[38828] <=  8'h00;      memory[38829] <=  8'h00;      memory[38830] <=  8'h00;      memory[38831] <=  8'h00;      memory[38832] <=  8'h00;      memory[38833] <=  8'h00;      memory[38834] <=  8'h00;      memory[38835] <=  8'h00;      memory[38836] <=  8'h00;      memory[38837] <=  8'h00;      memory[38838] <=  8'h00;      memory[38839] <=  8'h00;      memory[38840] <=  8'h00;      memory[38841] <=  8'h00;      memory[38842] <=  8'h00;      memory[38843] <=  8'h00;      memory[38844] <=  8'h00;      memory[38845] <=  8'h00;      memory[38846] <=  8'h00;      memory[38847] <=  8'h00;      memory[38848] <=  8'h00;      memory[38849] <=  8'h00;      memory[38850] <=  8'h00;      memory[38851] <=  8'h00;      memory[38852] <=  8'h00;      memory[38853] <=  8'h00;      memory[38854] <=  8'h00;      memory[38855] <=  8'h00;      memory[38856] <=  8'h00;      memory[38857] <=  8'h00;      memory[38858] <=  8'h00;      memory[38859] <=  8'h00;      memory[38860] <=  8'h00;      memory[38861] <=  8'h00;      memory[38862] <=  8'h00;      memory[38863] <=  8'h00;      memory[38864] <=  8'h00;      memory[38865] <=  8'h00;      memory[38866] <=  8'h00;      memory[38867] <=  8'h00;      memory[38868] <=  8'h00;      memory[38869] <=  8'h00;      memory[38870] <=  8'h00;      memory[38871] <=  8'h00;      memory[38872] <=  8'h00;      memory[38873] <=  8'h00;      memory[38874] <=  8'h00;      memory[38875] <=  8'h00;      memory[38876] <=  8'h00;      memory[38877] <=  8'h00;      memory[38878] <=  8'h00;      memory[38879] <=  8'h00;      memory[38880] <=  8'h00;      memory[38881] <=  8'h00;      memory[38882] <=  8'h00;      memory[38883] <=  8'h00;      memory[38884] <=  8'h00;      memory[38885] <=  8'h00;      memory[38886] <=  8'h00;      memory[38887] <=  8'h00;      memory[38888] <=  8'h00;      memory[38889] <=  8'h00;      memory[38890] <=  8'h00;      memory[38891] <=  8'h00;      memory[38892] <=  8'h00;      memory[38893] <=  8'h00;      memory[38894] <=  8'h00;      memory[38895] <=  8'h00;      memory[38896] <=  8'h00;      memory[38897] <=  8'h00;      memory[38898] <=  8'h00;      memory[38899] <=  8'h00;      memory[38900] <=  8'h00;      memory[38901] <=  8'h00;      memory[38902] <=  8'h00;      memory[38903] <=  8'h00;      memory[38904] <=  8'h00;      memory[38905] <=  8'h00;      memory[38906] <=  8'h00;      memory[38907] <=  8'h00;      memory[38908] <=  8'h00;      memory[38909] <=  8'h00;      memory[38910] <=  8'h00;      memory[38911] <=  8'h00;      memory[38912] <=  8'h00;      memory[38913] <=  8'h00;      memory[38914] <=  8'h00;      memory[38915] <=  8'h00;      memory[38916] <=  8'h00;      memory[38917] <=  8'h00;      memory[38918] <=  8'h00;      memory[38919] <=  8'h00;      memory[38920] <=  8'h00;      memory[38921] <=  8'h00;      memory[38922] <=  8'h00;      memory[38923] <=  8'h00;      memory[38924] <=  8'h00;      memory[38925] <=  8'h00;      memory[38926] <=  8'h00;      memory[38927] <=  8'h00;      memory[38928] <=  8'h00;      memory[38929] <=  8'h00;      memory[38930] <=  8'h00;      memory[38931] <=  8'h00;      memory[38932] <=  8'h00;      memory[38933] <=  8'h00;      memory[38934] <=  8'h00;      memory[38935] <=  8'h00;      memory[38936] <=  8'h00;      memory[38937] <=  8'h00;      memory[38938] <=  8'h00;      memory[38939] <=  8'h00;      memory[38940] <=  8'h00;      memory[38941] <=  8'h00;      memory[38942] <=  8'h00;      memory[38943] <=  8'h00;      memory[38944] <=  8'h00;      memory[38945] <=  8'h00;      memory[38946] <=  8'h00;      memory[38947] <=  8'h00;      memory[38948] <=  8'h00;      memory[38949] <=  8'h00;      memory[38950] <=  8'h00;      memory[38951] <=  8'h00;      memory[38952] <=  8'h00;      memory[38953] <=  8'h00;      memory[38954] <=  8'h00;      memory[38955] <=  8'h00;      memory[38956] <=  8'h00;      memory[38957] <=  8'h00;      memory[38958] <=  8'h00;      memory[38959] <=  8'h00;      memory[38960] <=  8'h00;      memory[38961] <=  8'h00;      memory[38962] <=  8'h00;      memory[38963] <=  8'h00;      memory[38964] <=  8'h00;      memory[38965] <=  8'h00;      memory[38966] <=  8'h00;      memory[38967] <=  8'h00;      memory[38968] <=  8'h00;      memory[38969] <=  8'h00;      memory[38970] <=  8'h00;      memory[38971] <=  8'h00;      memory[38972] <=  8'h00;      memory[38973] <=  8'h00;      memory[38974] <=  8'h00;      memory[38975] <=  8'h00;      memory[38976] <=  8'h00;      memory[38977] <=  8'h00;      memory[38978] <=  8'h00;      memory[38979] <=  8'h00;      memory[38980] <=  8'h00;      memory[38981] <=  8'h00;      memory[38982] <=  8'h00;      memory[38983] <=  8'h00;      memory[38984] <=  8'h00;      memory[38985] <=  8'h00;      memory[38986] <=  8'h00;      memory[38987] <=  8'h00;      memory[38988] <=  8'h00;      memory[38989] <=  8'h00;      memory[38990] <=  8'h00;      memory[38991] <=  8'h00;      memory[38992] <=  8'h00;      memory[38993] <=  8'h00;      memory[38994] <=  8'h00;      memory[38995] <=  8'h00;      memory[38996] <=  8'h00;      memory[38997] <=  8'h00;      memory[38998] <=  8'h00;      memory[38999] <=  8'h00;      memory[39000] <=  8'h00;      memory[39001] <=  8'h00;      memory[39002] <=  8'h00;      memory[39003] <=  8'h00;      memory[39004] <=  8'h00;      memory[39005] <=  8'h00;      memory[39006] <=  8'h00;      memory[39007] <=  8'h00;      memory[39008] <=  8'h00;      memory[39009] <=  8'h00;      memory[39010] <=  8'h00;      memory[39011] <=  8'h00;      memory[39012] <=  8'h00;      memory[39013] <=  8'h00;      memory[39014] <=  8'h00;      memory[39015] <=  8'h00;      memory[39016] <=  8'h00;      memory[39017] <=  8'h00;      memory[39018] <=  8'h00;      memory[39019] <=  8'h00;      memory[39020] <=  8'h00;      memory[39021] <=  8'h00;      memory[39022] <=  8'h00;      memory[39023] <=  8'h00;      memory[39024] <=  8'h00;      memory[39025] <=  8'h00;      memory[39026] <=  8'h00;      memory[39027] <=  8'h00;      memory[39028] <=  8'h00;      memory[39029] <=  8'h00;      memory[39030] <=  8'h00;      memory[39031] <=  8'h00;      memory[39032] <=  8'h00;      memory[39033] <=  8'h00;      memory[39034] <=  8'h00;      memory[39035] <=  8'h00;      memory[39036] <=  8'h00;      memory[39037] <=  8'h00;      memory[39038] <=  8'h00;      memory[39039] <=  8'h00;      memory[39040] <=  8'h00;      memory[39041] <=  8'h00;      memory[39042] <=  8'h00;      memory[39043] <=  8'h00;      memory[39044] <=  8'h00;      memory[39045] <=  8'h00;      memory[39046] <=  8'h00;      memory[39047] <=  8'h00;      memory[39048] <=  8'h00;      memory[39049] <=  8'h00;      memory[39050] <=  8'h00;      memory[39051] <=  8'h00;      memory[39052] <=  8'h00;      memory[39053] <=  8'h00;      memory[39054] <=  8'h00;      memory[39055] <=  8'h00;      memory[39056] <=  8'h00;      memory[39057] <=  8'h00;      memory[39058] <=  8'h00;      memory[39059] <=  8'h00;      memory[39060] <=  8'h00;      memory[39061] <=  8'h00;      memory[39062] <=  8'h00;      memory[39063] <=  8'h00;      memory[39064] <=  8'h00;      memory[39065] <=  8'h00;      memory[39066] <=  8'h00;      memory[39067] <=  8'h00;      memory[39068] <=  8'h00;      memory[39069] <=  8'h00;      memory[39070] <=  8'h00;      memory[39071] <=  8'h00;      memory[39072] <=  8'h00;      memory[39073] <=  8'h00;      memory[39074] <=  8'h00;      memory[39075] <=  8'h00;      memory[39076] <=  8'h00;      memory[39077] <=  8'h00;      memory[39078] <=  8'h00;      memory[39079] <=  8'h00;      memory[39080] <=  8'h00;      memory[39081] <=  8'h00;      memory[39082] <=  8'h00;      memory[39083] <=  8'h00;      memory[39084] <=  8'h00;      memory[39085] <=  8'h00;      memory[39086] <=  8'h00;      memory[39087] <=  8'h00;      memory[39088] <=  8'h00;      memory[39089] <=  8'h00;      memory[39090] <=  8'h00;      memory[39091] <=  8'h00;      memory[39092] <=  8'h00;      memory[39093] <=  8'h00;      memory[39094] <=  8'h00;      memory[39095] <=  8'h00;      memory[39096] <=  8'h00;      memory[39097] <=  8'h00;      memory[39098] <=  8'h00;      memory[39099] <=  8'h00;      memory[39100] <=  8'h00;      memory[39101] <=  8'h00;      memory[39102] <=  8'h00;      memory[39103] <=  8'h00;      memory[39104] <=  8'h00;      memory[39105] <=  8'h00;      memory[39106] <=  8'h00;      memory[39107] <=  8'h00;      memory[39108] <=  8'h00;      memory[39109] <=  8'h00;      memory[39110] <=  8'h00;      memory[39111] <=  8'h00;      memory[39112] <=  8'h00;      memory[39113] <=  8'h00;      memory[39114] <=  8'h00;      memory[39115] <=  8'h00;      memory[39116] <=  8'h00;      memory[39117] <=  8'h00;      memory[39118] <=  8'h00;      memory[39119] <=  8'h00;      memory[39120] <=  8'h00;      memory[39121] <=  8'h00;      memory[39122] <=  8'h00;      memory[39123] <=  8'h00;      memory[39124] <=  8'h00;      memory[39125] <=  8'h00;      memory[39126] <=  8'h00;      memory[39127] <=  8'h00;      memory[39128] <=  8'h00;      memory[39129] <=  8'h00;      memory[39130] <=  8'h00;      memory[39131] <=  8'h00;      memory[39132] <=  8'h00;      memory[39133] <=  8'h00;      memory[39134] <=  8'h00;      memory[39135] <=  8'h00;      memory[39136] <=  8'h00;      memory[39137] <=  8'h00;      memory[39138] <=  8'h00;      memory[39139] <=  8'h00;      memory[39140] <=  8'h00;      memory[39141] <=  8'h00;      memory[39142] <=  8'h00;      memory[39143] <=  8'h00;      memory[39144] <=  8'h00;      memory[39145] <=  8'h00;      memory[39146] <=  8'h00;      memory[39147] <=  8'h00;      memory[39148] <=  8'h00;      memory[39149] <=  8'h00;      memory[39150] <=  8'h00;      memory[39151] <=  8'h00;      memory[39152] <=  8'h00;      memory[39153] <=  8'h00;      memory[39154] <=  8'h00;      memory[39155] <=  8'h00;      memory[39156] <=  8'h00;      memory[39157] <=  8'h00;      memory[39158] <=  8'h00;      memory[39159] <=  8'h00;      memory[39160] <=  8'h00;      memory[39161] <=  8'h00;      memory[39162] <=  8'h00;      memory[39163] <=  8'h00;      memory[39164] <=  8'h00;      memory[39165] <=  8'h00;      memory[39166] <=  8'h00;      memory[39167] <=  8'h00;      memory[39168] <=  8'h00;      memory[39169] <=  8'h00;      memory[39170] <=  8'h00;      memory[39171] <=  8'h00;      memory[39172] <=  8'h00;      memory[39173] <=  8'h00;      memory[39174] <=  8'h00;      memory[39175] <=  8'h00;      memory[39176] <=  8'h00;      memory[39177] <=  8'h00;      memory[39178] <=  8'h00;      memory[39179] <=  8'h00;      memory[39180] <=  8'h00;      memory[39181] <=  8'h00;      memory[39182] <=  8'h00;      memory[39183] <=  8'h00;      memory[39184] <=  8'h00;      memory[39185] <=  8'h00;      memory[39186] <=  8'h00;      memory[39187] <=  8'h00;      memory[39188] <=  8'h00;      memory[39189] <=  8'h00;      memory[39190] <=  8'h00;      memory[39191] <=  8'h00;      memory[39192] <=  8'h00;      memory[39193] <=  8'h00;      memory[39194] <=  8'h00;      memory[39195] <=  8'h00;      memory[39196] <=  8'h00;      memory[39197] <=  8'h00;      memory[39198] <=  8'h00;      memory[39199] <=  8'h00;      memory[39200] <=  8'h00;      memory[39201] <=  8'h00;      memory[39202] <=  8'h00;      memory[39203] <=  8'h00;      memory[39204] <=  8'h00;      memory[39205] <=  8'h00;      memory[39206] <=  8'h00;      memory[39207] <=  8'h00;      memory[39208] <=  8'h00;      memory[39209] <=  8'h00;      memory[39210] <=  8'h00;      memory[39211] <=  8'h00;      memory[39212] <=  8'h00;      memory[39213] <=  8'h00;      memory[39214] <=  8'h00;      memory[39215] <=  8'h00;      memory[39216] <=  8'h00;      memory[39217] <=  8'h00;      memory[39218] <=  8'h00;      memory[39219] <=  8'h00;      memory[39220] <=  8'h00;      memory[39221] <=  8'h00;      memory[39222] <=  8'h00;      memory[39223] <=  8'h00;      memory[39224] <=  8'h00;      memory[39225] <=  8'h00;      memory[39226] <=  8'h00;      memory[39227] <=  8'h00;      memory[39228] <=  8'h00;      memory[39229] <=  8'h00;      memory[39230] <=  8'h00;      memory[39231] <=  8'h00;      memory[39232] <=  8'h00;      memory[39233] <=  8'h00;      memory[39234] <=  8'h00;      memory[39235] <=  8'h00;      memory[39236] <=  8'h00;      memory[39237] <=  8'h00;      memory[39238] <=  8'h00;      memory[39239] <=  8'h00;      memory[39240] <=  8'h00;      memory[39241] <=  8'h00;      memory[39242] <=  8'h00;      memory[39243] <=  8'h00;      memory[39244] <=  8'h00;      memory[39245] <=  8'h00;      memory[39246] <=  8'h00;      memory[39247] <=  8'h00;      memory[39248] <=  8'h00;      memory[39249] <=  8'h00;      memory[39250] <=  8'h00;      memory[39251] <=  8'h00;      memory[39252] <=  8'h00;      memory[39253] <=  8'h00;      memory[39254] <=  8'h00;      memory[39255] <=  8'h00;      memory[39256] <=  8'h00;      memory[39257] <=  8'h00;      memory[39258] <=  8'h00;      memory[39259] <=  8'h00;      memory[39260] <=  8'h00;      memory[39261] <=  8'h00;      memory[39262] <=  8'h00;      memory[39263] <=  8'h00;      memory[39264] <=  8'h00;      memory[39265] <=  8'h00;      memory[39266] <=  8'h00;      memory[39267] <=  8'h00;      memory[39268] <=  8'h00;      memory[39269] <=  8'h00;      memory[39270] <=  8'h00;      memory[39271] <=  8'h00;      memory[39272] <=  8'h00;      memory[39273] <=  8'h00;      memory[39274] <=  8'h00;      memory[39275] <=  8'h00;      memory[39276] <=  8'h00;      memory[39277] <=  8'h00;      memory[39278] <=  8'h00;      memory[39279] <=  8'h00;      memory[39280] <=  8'h00;      memory[39281] <=  8'h00;      memory[39282] <=  8'h00;      memory[39283] <=  8'h00;      memory[39284] <=  8'h00;      memory[39285] <=  8'h00;      memory[39286] <=  8'h00;      memory[39287] <=  8'h00;      memory[39288] <=  8'h00;      memory[39289] <=  8'h00;      memory[39290] <=  8'h00;      memory[39291] <=  8'h00;      memory[39292] <=  8'h00;      memory[39293] <=  8'h00;      memory[39294] <=  8'h00;      memory[39295] <=  8'h00;      memory[39296] <=  8'h00;      memory[39297] <=  8'h00;      memory[39298] <=  8'h00;      memory[39299] <=  8'h00;      memory[39300] <=  8'h00;      memory[39301] <=  8'h00;      memory[39302] <=  8'h00;      memory[39303] <=  8'h00;      memory[39304] <=  8'h00;      memory[39305] <=  8'h00;      memory[39306] <=  8'h00;      memory[39307] <=  8'h00;      memory[39308] <=  8'h00;      memory[39309] <=  8'h00;      memory[39310] <=  8'h00;      memory[39311] <=  8'h00;      memory[39312] <=  8'h00;      memory[39313] <=  8'h00;      memory[39314] <=  8'h00;      memory[39315] <=  8'h00;      memory[39316] <=  8'h00;      memory[39317] <=  8'h00;      memory[39318] <=  8'h00;      memory[39319] <=  8'h00;      memory[39320] <=  8'h00;      memory[39321] <=  8'h00;      memory[39322] <=  8'h00;      memory[39323] <=  8'h00;      memory[39324] <=  8'h00;      memory[39325] <=  8'h00;      memory[39326] <=  8'h00;      memory[39327] <=  8'h00;      memory[39328] <=  8'h00;      memory[39329] <=  8'h00;      memory[39330] <=  8'h00;      memory[39331] <=  8'h00;      memory[39332] <=  8'h00;      memory[39333] <=  8'h00;      memory[39334] <=  8'h00;      memory[39335] <=  8'h00;      memory[39336] <=  8'h00;      memory[39337] <=  8'h00;      memory[39338] <=  8'h00;      memory[39339] <=  8'h00;      memory[39340] <=  8'h00;      memory[39341] <=  8'h00;      memory[39342] <=  8'h00;      memory[39343] <=  8'h00;      memory[39344] <=  8'h00;      memory[39345] <=  8'h00;      memory[39346] <=  8'h00;      memory[39347] <=  8'h00;      memory[39348] <=  8'h00;      memory[39349] <=  8'h00;      memory[39350] <=  8'h00;      memory[39351] <=  8'h00;      memory[39352] <=  8'h00;      memory[39353] <=  8'h00;      memory[39354] <=  8'h00;      memory[39355] <=  8'h00;      memory[39356] <=  8'h00;      memory[39357] <=  8'h00;      memory[39358] <=  8'h00;      memory[39359] <=  8'h00;      memory[39360] <=  8'h00;      memory[39361] <=  8'h00;      memory[39362] <=  8'h00;      memory[39363] <=  8'h00;      memory[39364] <=  8'h00;      memory[39365] <=  8'h00;      memory[39366] <=  8'h00;      memory[39367] <=  8'h00;      memory[39368] <=  8'h00;      memory[39369] <=  8'h00;      memory[39370] <=  8'h00;      memory[39371] <=  8'h00;      memory[39372] <=  8'h00;      memory[39373] <=  8'h00;      memory[39374] <=  8'h00;      memory[39375] <=  8'h00;      memory[39376] <=  8'h00;      memory[39377] <=  8'h00;      memory[39378] <=  8'h00;      memory[39379] <=  8'h00;      memory[39380] <=  8'h00;      memory[39381] <=  8'h00;      memory[39382] <=  8'h00;      memory[39383] <=  8'h00;      memory[39384] <=  8'h00;      memory[39385] <=  8'h00;      memory[39386] <=  8'h00;      memory[39387] <=  8'h00;      memory[39388] <=  8'h00;      memory[39389] <=  8'h00;      memory[39390] <=  8'h00;      memory[39391] <=  8'h00;      memory[39392] <=  8'h00;      memory[39393] <=  8'h00;      memory[39394] <=  8'h00;      memory[39395] <=  8'h00;      memory[39396] <=  8'h00;      memory[39397] <=  8'h00;      memory[39398] <=  8'h00;      memory[39399] <=  8'h00;      memory[39400] <=  8'h00;      memory[39401] <=  8'h00;      memory[39402] <=  8'h00;      memory[39403] <=  8'h00;      memory[39404] <=  8'h00;      memory[39405] <=  8'h00;      memory[39406] <=  8'h00;      memory[39407] <=  8'h00;      memory[39408] <=  8'h00;      memory[39409] <=  8'h00;      memory[39410] <=  8'h00;      memory[39411] <=  8'h00;      memory[39412] <=  8'h00;      memory[39413] <=  8'h00;      memory[39414] <=  8'h00;      memory[39415] <=  8'h00;      memory[39416] <=  8'h00;      memory[39417] <=  8'h00;      memory[39418] <=  8'h00;      memory[39419] <=  8'h00;      memory[39420] <=  8'h00;      memory[39421] <=  8'h00;      memory[39422] <=  8'h00;      memory[39423] <=  8'h00;      memory[39424] <=  8'h00;      memory[39425] <=  8'h00;      memory[39426] <=  8'h00;      memory[39427] <=  8'h00;      memory[39428] <=  8'h00;      memory[39429] <=  8'h00;      memory[39430] <=  8'h00;      memory[39431] <=  8'h00;      memory[39432] <=  8'h00;      memory[39433] <=  8'h00;      memory[39434] <=  8'h00;      memory[39435] <=  8'h00;      memory[39436] <=  8'h00;      memory[39437] <=  8'h00;      memory[39438] <=  8'h00;      memory[39439] <=  8'h00;      memory[39440] <=  8'h00;      memory[39441] <=  8'h00;      memory[39442] <=  8'h00;      memory[39443] <=  8'h00;      memory[39444] <=  8'h00;      memory[39445] <=  8'h00;      memory[39446] <=  8'h00;      memory[39447] <=  8'h00;      memory[39448] <=  8'h00;      memory[39449] <=  8'h00;      memory[39450] <=  8'h00;      memory[39451] <=  8'h00;      memory[39452] <=  8'h00;      memory[39453] <=  8'h00;      memory[39454] <=  8'h00;      memory[39455] <=  8'h00;      memory[39456] <=  8'h00;      memory[39457] <=  8'h00;      memory[39458] <=  8'h00;      memory[39459] <=  8'h00;      memory[39460] <=  8'h00;      memory[39461] <=  8'h00;      memory[39462] <=  8'h00;      memory[39463] <=  8'h00;      memory[39464] <=  8'h00;      memory[39465] <=  8'h00;      memory[39466] <=  8'h00;      memory[39467] <=  8'h00;      memory[39468] <=  8'h00;      memory[39469] <=  8'h00;      memory[39470] <=  8'h00;      memory[39471] <=  8'h00;      memory[39472] <=  8'h00;      memory[39473] <=  8'h00;      memory[39474] <=  8'h00;      memory[39475] <=  8'h00;      memory[39476] <=  8'h00;      memory[39477] <=  8'h00;      memory[39478] <=  8'h00;      memory[39479] <=  8'h00;      memory[39480] <=  8'h00;      memory[39481] <=  8'h00;      memory[39482] <=  8'h00;      memory[39483] <=  8'h00;      memory[39484] <=  8'h00;      memory[39485] <=  8'h00;      memory[39486] <=  8'h00;      memory[39487] <=  8'h00;      memory[39488] <=  8'h00;      memory[39489] <=  8'h00;      memory[39490] <=  8'h00;      memory[39491] <=  8'h00;      memory[39492] <=  8'h00;      memory[39493] <=  8'h00;      memory[39494] <=  8'h00;      memory[39495] <=  8'h00;      memory[39496] <=  8'h00;      memory[39497] <=  8'h00;      memory[39498] <=  8'h00;      memory[39499] <=  8'h00;      memory[39500] <=  8'h00;      memory[39501] <=  8'h00;      memory[39502] <=  8'h00;      memory[39503] <=  8'h00;      memory[39504] <=  8'h00;      memory[39505] <=  8'h00;      memory[39506] <=  8'h00;      memory[39507] <=  8'h00;      memory[39508] <=  8'h00;      memory[39509] <=  8'h00;      memory[39510] <=  8'h00;      memory[39511] <=  8'h00;      memory[39512] <=  8'h00;      memory[39513] <=  8'h00;      memory[39514] <=  8'h00;      memory[39515] <=  8'h00;      memory[39516] <=  8'h00;      memory[39517] <=  8'h00;      memory[39518] <=  8'h00;      memory[39519] <=  8'h00;      memory[39520] <=  8'h00;      memory[39521] <=  8'h00;      memory[39522] <=  8'h00;      memory[39523] <=  8'h00;      memory[39524] <=  8'h00;      memory[39525] <=  8'h00;      memory[39526] <=  8'h00;      memory[39527] <=  8'h00;      memory[39528] <=  8'h00;      memory[39529] <=  8'h00;      memory[39530] <=  8'h00;      memory[39531] <=  8'h00;      memory[39532] <=  8'h00;      memory[39533] <=  8'h00;      memory[39534] <=  8'h00;      memory[39535] <=  8'h00;      memory[39536] <=  8'h00;      memory[39537] <=  8'h00;      memory[39538] <=  8'h00;      memory[39539] <=  8'h00;      memory[39540] <=  8'h00;      memory[39541] <=  8'h00;      memory[39542] <=  8'h00;      memory[39543] <=  8'h00;      memory[39544] <=  8'h00;      memory[39545] <=  8'h00;      memory[39546] <=  8'h00;      memory[39547] <=  8'h00;      memory[39548] <=  8'h00;      memory[39549] <=  8'h00;      memory[39550] <=  8'h00;      memory[39551] <=  8'h00;      memory[39552] <=  8'h00;      memory[39553] <=  8'h00;      memory[39554] <=  8'h00;      memory[39555] <=  8'h00;      memory[39556] <=  8'h00;      memory[39557] <=  8'h00;      memory[39558] <=  8'h00;      memory[39559] <=  8'h00;      memory[39560] <=  8'h00;      memory[39561] <=  8'h00;      memory[39562] <=  8'h00;      memory[39563] <=  8'h00;      memory[39564] <=  8'h00;      memory[39565] <=  8'h00;      memory[39566] <=  8'h00;      memory[39567] <=  8'h00;      memory[39568] <=  8'h00;      memory[39569] <=  8'h00;      memory[39570] <=  8'h00;      memory[39571] <=  8'h00;      memory[39572] <=  8'h00;      memory[39573] <=  8'h00;      memory[39574] <=  8'h00;      memory[39575] <=  8'h00;      memory[39576] <=  8'h00;      memory[39577] <=  8'h00;      memory[39578] <=  8'h00;      memory[39579] <=  8'h00;      memory[39580] <=  8'h00;      memory[39581] <=  8'h00;      memory[39582] <=  8'h00;      memory[39583] <=  8'h00;      memory[39584] <=  8'h00;      memory[39585] <=  8'h00;      memory[39586] <=  8'h00;      memory[39587] <=  8'h00;      memory[39588] <=  8'h00;      memory[39589] <=  8'h00;      memory[39590] <=  8'h00;      memory[39591] <=  8'h00;      memory[39592] <=  8'h00;      memory[39593] <=  8'h00;      memory[39594] <=  8'h00;      memory[39595] <=  8'h00;      memory[39596] <=  8'h00;      memory[39597] <=  8'h00;      memory[39598] <=  8'h00;      memory[39599] <=  8'h00;      memory[39600] <=  8'h00;      memory[39601] <=  8'h00;      memory[39602] <=  8'h00;      memory[39603] <=  8'h00;      memory[39604] <=  8'h00;      memory[39605] <=  8'h00;      memory[39606] <=  8'h00;      memory[39607] <=  8'h00;      memory[39608] <=  8'h00;      memory[39609] <=  8'h00;      memory[39610] <=  8'h00;      memory[39611] <=  8'h00;      memory[39612] <=  8'h00;      memory[39613] <=  8'h00;      memory[39614] <=  8'h00;      memory[39615] <=  8'h00;      memory[39616] <=  8'h00;      memory[39617] <=  8'h00;      memory[39618] <=  8'h00;      memory[39619] <=  8'h00;      memory[39620] <=  8'h00;      memory[39621] <=  8'h00;      memory[39622] <=  8'h00;      memory[39623] <=  8'h00;      memory[39624] <=  8'h00;      memory[39625] <=  8'h00;      memory[39626] <=  8'h00;      memory[39627] <=  8'h00;      memory[39628] <=  8'h00;      memory[39629] <=  8'h00;      memory[39630] <=  8'h00;      memory[39631] <=  8'h00;      memory[39632] <=  8'h00;      memory[39633] <=  8'h00;      memory[39634] <=  8'h00;      memory[39635] <=  8'h00;      memory[39636] <=  8'h00;      memory[39637] <=  8'h00;      memory[39638] <=  8'h00;      memory[39639] <=  8'h00;      memory[39640] <=  8'h00;      memory[39641] <=  8'h00;      memory[39642] <=  8'h00;      memory[39643] <=  8'h00;      memory[39644] <=  8'h00;      memory[39645] <=  8'h00;      memory[39646] <=  8'h00;      memory[39647] <=  8'h00;      memory[39648] <=  8'h00;      memory[39649] <=  8'h00;      memory[39650] <=  8'h00;      memory[39651] <=  8'h00;      memory[39652] <=  8'h00;      memory[39653] <=  8'h00;      memory[39654] <=  8'h00;      memory[39655] <=  8'h00;      memory[39656] <=  8'h00;      memory[39657] <=  8'h00;      memory[39658] <=  8'h00;      memory[39659] <=  8'h00;      memory[39660] <=  8'h00;      memory[39661] <=  8'h00;      memory[39662] <=  8'h00;      memory[39663] <=  8'h00;      memory[39664] <=  8'h00;      memory[39665] <=  8'h00;      memory[39666] <=  8'h00;      memory[39667] <=  8'h00;      memory[39668] <=  8'h00;      memory[39669] <=  8'h00;      memory[39670] <=  8'h00;      memory[39671] <=  8'h00;      memory[39672] <=  8'h00;      memory[39673] <=  8'h00;      memory[39674] <=  8'h00;      memory[39675] <=  8'h00;      memory[39676] <=  8'h00;      memory[39677] <=  8'h00;      memory[39678] <=  8'h00;      memory[39679] <=  8'h00;      memory[39680] <=  8'h00;      memory[39681] <=  8'h00;      memory[39682] <=  8'h00;      memory[39683] <=  8'h00;      memory[39684] <=  8'h00;      memory[39685] <=  8'h00;      memory[39686] <=  8'h00;      memory[39687] <=  8'h00;      memory[39688] <=  8'h00;      memory[39689] <=  8'h00;      memory[39690] <=  8'h00;      memory[39691] <=  8'h00;      memory[39692] <=  8'h00;      memory[39693] <=  8'h00;      memory[39694] <=  8'h00;      memory[39695] <=  8'h00;      memory[39696] <=  8'h00;      memory[39697] <=  8'h00;      memory[39698] <=  8'h00;      memory[39699] <=  8'h00;      memory[39700] <=  8'h00;      memory[39701] <=  8'h00;      memory[39702] <=  8'h00;      memory[39703] <=  8'h00;      memory[39704] <=  8'h00;      memory[39705] <=  8'h00;      memory[39706] <=  8'h00;      memory[39707] <=  8'h00;      memory[39708] <=  8'h00;      memory[39709] <=  8'h00;      memory[39710] <=  8'h00;      memory[39711] <=  8'h00;      memory[39712] <=  8'h00;      memory[39713] <=  8'h00;      memory[39714] <=  8'h00;      memory[39715] <=  8'h00;      memory[39716] <=  8'h00;      memory[39717] <=  8'h00;      memory[39718] <=  8'h00;      memory[39719] <=  8'h00;      memory[39720] <=  8'h00;      memory[39721] <=  8'h00;      memory[39722] <=  8'h00;      memory[39723] <=  8'h00;      memory[39724] <=  8'h00;      memory[39725] <=  8'h00;      memory[39726] <=  8'h00;      memory[39727] <=  8'h00;      memory[39728] <=  8'h00;      memory[39729] <=  8'h00;      memory[39730] <=  8'h00;      memory[39731] <=  8'h00;      memory[39732] <=  8'h00;      memory[39733] <=  8'h00;      memory[39734] <=  8'h00;      memory[39735] <=  8'h00;      memory[39736] <=  8'h00;      memory[39737] <=  8'h00;      memory[39738] <=  8'h00;      memory[39739] <=  8'h00;      memory[39740] <=  8'h00;      memory[39741] <=  8'h00;      memory[39742] <=  8'h00;      memory[39743] <=  8'h00;      memory[39744] <=  8'h00;      memory[39745] <=  8'h00;      memory[39746] <=  8'h00;      memory[39747] <=  8'h00;      memory[39748] <=  8'h00;      memory[39749] <=  8'h00;      memory[39750] <=  8'h00;      memory[39751] <=  8'h00;      memory[39752] <=  8'h00;      memory[39753] <=  8'h00;      memory[39754] <=  8'h00;      memory[39755] <=  8'h00;      memory[39756] <=  8'h00;      memory[39757] <=  8'h00;      memory[39758] <=  8'h00;      memory[39759] <=  8'h00;      memory[39760] <=  8'h00;      memory[39761] <=  8'h00;      memory[39762] <=  8'h00;      memory[39763] <=  8'h00;      memory[39764] <=  8'h00;      memory[39765] <=  8'h00;      memory[39766] <=  8'h00;      memory[39767] <=  8'h00;      memory[39768] <=  8'h00;      memory[39769] <=  8'h00;      memory[39770] <=  8'h00;      memory[39771] <=  8'h00;      memory[39772] <=  8'h00;      memory[39773] <=  8'h00;      memory[39774] <=  8'h00;      memory[39775] <=  8'h00;      memory[39776] <=  8'h00;      memory[39777] <=  8'h00;      memory[39778] <=  8'h00;      memory[39779] <=  8'h00;      memory[39780] <=  8'h00;      memory[39781] <=  8'h00;      memory[39782] <=  8'h00;      memory[39783] <=  8'h00;      memory[39784] <=  8'h00;      memory[39785] <=  8'h00;      memory[39786] <=  8'h00;      memory[39787] <=  8'h00;      memory[39788] <=  8'h00;      memory[39789] <=  8'h00;      memory[39790] <=  8'h00;      memory[39791] <=  8'h00;      memory[39792] <=  8'h00;      memory[39793] <=  8'h00;      memory[39794] <=  8'h00;      memory[39795] <=  8'h00;      memory[39796] <=  8'h00;      memory[39797] <=  8'h00;      memory[39798] <=  8'h00;      memory[39799] <=  8'h00;      memory[39800] <=  8'h00;      memory[39801] <=  8'h00;      memory[39802] <=  8'h00;      memory[39803] <=  8'h00;      memory[39804] <=  8'h00;      memory[39805] <=  8'h00;      memory[39806] <=  8'h00;      memory[39807] <=  8'h00;      memory[39808] <=  8'h00;      memory[39809] <=  8'h00;      memory[39810] <=  8'h00;      memory[39811] <=  8'h00;      memory[39812] <=  8'h00;      memory[39813] <=  8'h00;      memory[39814] <=  8'h00;      memory[39815] <=  8'h00;      memory[39816] <=  8'h00;      memory[39817] <=  8'h00;      memory[39818] <=  8'h00;      memory[39819] <=  8'h00;      memory[39820] <=  8'h00;      memory[39821] <=  8'h00;      memory[39822] <=  8'h00;      memory[39823] <=  8'h00;      memory[39824] <=  8'h00;      memory[39825] <=  8'h00;      memory[39826] <=  8'h00;      memory[39827] <=  8'h00;      memory[39828] <=  8'h00;      memory[39829] <=  8'h00;      memory[39830] <=  8'h00;      memory[39831] <=  8'h00;      memory[39832] <=  8'h00;      memory[39833] <=  8'h00;      memory[39834] <=  8'h00;      memory[39835] <=  8'h00;      memory[39836] <=  8'h00;      memory[39837] <=  8'h00;      memory[39838] <=  8'h00;      memory[39839] <=  8'h00;      memory[39840] <=  8'h00;      memory[39841] <=  8'h00;      memory[39842] <=  8'h00;      memory[39843] <=  8'h00;      memory[39844] <=  8'h00;      memory[39845] <=  8'h00;      memory[39846] <=  8'h00;      memory[39847] <=  8'h00;      memory[39848] <=  8'h00;      memory[39849] <=  8'h00;      memory[39850] <=  8'h00;      memory[39851] <=  8'h00;      memory[39852] <=  8'h00;      memory[39853] <=  8'h00;      memory[39854] <=  8'h00;      memory[39855] <=  8'h00;      memory[39856] <=  8'h00;      memory[39857] <=  8'h00;      memory[39858] <=  8'h00;      memory[39859] <=  8'h00;      memory[39860] <=  8'h00;      memory[39861] <=  8'h00;      memory[39862] <=  8'h00;      memory[39863] <=  8'h00;      memory[39864] <=  8'h00;      memory[39865] <=  8'h00;      memory[39866] <=  8'h00;      memory[39867] <=  8'h00;      memory[39868] <=  8'h00;      memory[39869] <=  8'h00;      memory[39870] <=  8'h00;      memory[39871] <=  8'h00;      memory[39872] <=  8'h00;      memory[39873] <=  8'h00;      memory[39874] <=  8'h00;      memory[39875] <=  8'h00;      memory[39876] <=  8'h00;      memory[39877] <=  8'h00;      memory[39878] <=  8'h00;      memory[39879] <=  8'h00;      memory[39880] <=  8'h00;      memory[39881] <=  8'h00;      memory[39882] <=  8'h00;      memory[39883] <=  8'h00;      memory[39884] <=  8'h00;      memory[39885] <=  8'h00;      memory[39886] <=  8'h00;      memory[39887] <=  8'h00;      memory[39888] <=  8'h00;      memory[39889] <=  8'h00;      memory[39890] <=  8'h00;      memory[39891] <=  8'h00;      memory[39892] <=  8'h00;      memory[39893] <=  8'h00;      memory[39894] <=  8'h00;      memory[39895] <=  8'h00;      memory[39896] <=  8'h00;      memory[39897] <=  8'h00;      memory[39898] <=  8'h00;      memory[39899] <=  8'h00;      memory[39900] <=  8'h00;      memory[39901] <=  8'h00;      memory[39902] <=  8'h00;      memory[39903] <=  8'h00;      memory[39904] <=  8'h00;      memory[39905] <=  8'h00;      memory[39906] <=  8'h00;      memory[39907] <=  8'h00;      memory[39908] <=  8'h00;      memory[39909] <=  8'h00;      memory[39910] <=  8'h00;      memory[39911] <=  8'h00;      memory[39912] <=  8'h00;      memory[39913] <=  8'h00;      memory[39914] <=  8'h00;      memory[39915] <=  8'h00;      memory[39916] <=  8'h00;      memory[39917] <=  8'h00;      memory[39918] <=  8'h00;      memory[39919] <=  8'h00;      memory[39920] <=  8'h00;      memory[39921] <=  8'h00;      memory[39922] <=  8'h00;      memory[39923] <=  8'h00;      memory[39924] <=  8'h00;      memory[39925] <=  8'h00;      memory[39926] <=  8'h00;      memory[39927] <=  8'h00;      memory[39928] <=  8'h00;      memory[39929] <=  8'h00;      memory[39930] <=  8'h00;      memory[39931] <=  8'h00;      memory[39932] <=  8'h00;      memory[39933] <=  8'h00;      memory[39934] <=  8'h00;      memory[39935] <=  8'h00;      memory[39936] <=  8'h00;      memory[39937] <=  8'h00;      memory[39938] <=  8'h00;      memory[39939] <=  8'h00;      memory[39940] <=  8'h00;      memory[39941] <=  8'h00;      memory[39942] <=  8'h00;      memory[39943] <=  8'h00;      memory[39944] <=  8'h00;      memory[39945] <=  8'h00;      memory[39946] <=  8'h00;      memory[39947] <=  8'h00;      memory[39948] <=  8'h00;      memory[39949] <=  8'h00;      memory[39950] <=  8'h00;      memory[39951] <=  8'h00;      memory[39952] <=  8'h00;      memory[39953] <=  8'h00;      memory[39954] <=  8'h00;      memory[39955] <=  8'h00;      memory[39956] <=  8'h00;      memory[39957] <=  8'h00;      memory[39958] <=  8'h00;      memory[39959] <=  8'h00;      memory[39960] <=  8'h00;      memory[39961] <=  8'h00;      memory[39962] <=  8'h00;      memory[39963] <=  8'h00;      memory[39964] <=  8'h00;      memory[39965] <=  8'h00;      memory[39966] <=  8'h00;      memory[39967] <=  8'h00;      memory[39968] <=  8'h00;      memory[39969] <=  8'h00;      memory[39970] <=  8'h00;      memory[39971] <=  8'h00;      memory[39972] <=  8'h00;      memory[39973] <=  8'h00;      memory[39974] <=  8'h00;      memory[39975] <=  8'h00;      memory[39976] <=  8'h00;      memory[39977] <=  8'h00;      memory[39978] <=  8'h00;      memory[39979] <=  8'h00;      memory[39980] <=  8'h00;      memory[39981] <=  8'h00;      memory[39982] <=  8'h00;      memory[39983] <=  8'h00;      memory[39984] <=  8'h00;      memory[39985] <=  8'h00;      memory[39986] <=  8'h00;      memory[39987] <=  8'h00;      memory[39988] <=  8'h00;      memory[39989] <=  8'h00;      memory[39990] <=  8'h00;      memory[39991] <=  8'h00;      memory[39992] <=  8'h00;      memory[39993] <=  8'h00;      memory[39994] <=  8'h00;      memory[39995] <=  8'h00;      memory[39996] <=  8'h00;      memory[39997] <=  8'h00;      memory[39998] <=  8'h00;      memory[39999] <=  8'h00;      memory[40000] <=  8'h00;      memory[40001] <=  8'h00;      memory[40002] <=  8'h00;      memory[40003] <=  8'h00;      memory[40004] <=  8'h00;      memory[40005] <=  8'h00;      memory[40006] <=  8'h00;      memory[40007] <=  8'h00;      memory[40008] <=  8'h00;      memory[40009] <=  8'h00;      memory[40010] <=  8'h00;      memory[40011] <=  8'h00;      memory[40012] <=  8'h00;      memory[40013] <=  8'h00;      memory[40014] <=  8'h00;      memory[40015] <=  8'h00;      memory[40016] <=  8'h00;      memory[40017] <=  8'h00;      memory[40018] <=  8'h00;      memory[40019] <=  8'h00;      memory[40020] <=  8'h00;      memory[40021] <=  8'h00;      memory[40022] <=  8'h00;      memory[40023] <=  8'h00;      memory[40024] <=  8'h00;      memory[40025] <=  8'h00;      memory[40026] <=  8'h00;      memory[40027] <=  8'h00;      memory[40028] <=  8'h00;      memory[40029] <=  8'h00;      memory[40030] <=  8'h00;      memory[40031] <=  8'h00;      memory[40032] <=  8'h00;      memory[40033] <=  8'h00;      memory[40034] <=  8'h00;      memory[40035] <=  8'h00;      memory[40036] <=  8'h00;      memory[40037] <=  8'h00;      memory[40038] <=  8'h00;      memory[40039] <=  8'h00;      memory[40040] <=  8'h00;      memory[40041] <=  8'h00;      memory[40042] <=  8'h00;      memory[40043] <=  8'h00;      memory[40044] <=  8'h00;      memory[40045] <=  8'h00;      memory[40046] <=  8'h00;      memory[40047] <=  8'h00;      memory[40048] <=  8'h00;      memory[40049] <=  8'h00;      memory[40050] <=  8'h00;      memory[40051] <=  8'h00;      memory[40052] <=  8'h00;      memory[40053] <=  8'h00;      memory[40054] <=  8'h00;      memory[40055] <=  8'h00;      memory[40056] <=  8'h00;      memory[40057] <=  8'h00;      memory[40058] <=  8'h00;      memory[40059] <=  8'h00;      memory[40060] <=  8'h00;      memory[40061] <=  8'h00;      memory[40062] <=  8'h00;      memory[40063] <=  8'h00;      memory[40064] <=  8'h00;      memory[40065] <=  8'h00;      memory[40066] <=  8'h00;      memory[40067] <=  8'h00;      memory[40068] <=  8'h00;      memory[40069] <=  8'h00;      memory[40070] <=  8'h00;      memory[40071] <=  8'h00;      memory[40072] <=  8'h00;      memory[40073] <=  8'h00;      memory[40074] <=  8'h00;      memory[40075] <=  8'h00;      memory[40076] <=  8'h00;      memory[40077] <=  8'h00;      memory[40078] <=  8'h00;      memory[40079] <=  8'h00;      memory[40080] <=  8'h00;      memory[40081] <=  8'h00;      memory[40082] <=  8'h00;      memory[40083] <=  8'h00;      memory[40084] <=  8'h00;      memory[40085] <=  8'h00;      memory[40086] <=  8'h00;      memory[40087] <=  8'h00;      memory[40088] <=  8'h00;      memory[40089] <=  8'h00;      memory[40090] <=  8'h00;      memory[40091] <=  8'h00;      memory[40092] <=  8'h00;      memory[40093] <=  8'h00;      memory[40094] <=  8'h00;      memory[40095] <=  8'h00;      memory[40096] <=  8'h00;      memory[40097] <=  8'h00;      memory[40098] <=  8'h00;      memory[40099] <=  8'h00;      memory[40100] <=  8'h00;      memory[40101] <=  8'h00;      memory[40102] <=  8'h00;      memory[40103] <=  8'h00;      memory[40104] <=  8'h00;      memory[40105] <=  8'h00;      memory[40106] <=  8'h00;      memory[40107] <=  8'h00;      memory[40108] <=  8'h00;      memory[40109] <=  8'h00;      memory[40110] <=  8'h00;      memory[40111] <=  8'h00;      memory[40112] <=  8'h00;      memory[40113] <=  8'h00;      memory[40114] <=  8'h00;      memory[40115] <=  8'h00;      memory[40116] <=  8'h00;      memory[40117] <=  8'h00;      memory[40118] <=  8'h00;      memory[40119] <=  8'h00;      memory[40120] <=  8'h00;      memory[40121] <=  8'h00;      memory[40122] <=  8'h00;      memory[40123] <=  8'h00;      memory[40124] <=  8'h00;      memory[40125] <=  8'h00;      memory[40126] <=  8'h00;      memory[40127] <=  8'h00;      memory[40128] <=  8'h00;      memory[40129] <=  8'h00;      memory[40130] <=  8'h00;      memory[40131] <=  8'h00;      memory[40132] <=  8'h00;      memory[40133] <=  8'h00;      memory[40134] <=  8'h00;      memory[40135] <=  8'h00;      memory[40136] <=  8'h00;      memory[40137] <=  8'h00;      memory[40138] <=  8'h00;      memory[40139] <=  8'h00;      memory[40140] <=  8'h00;      memory[40141] <=  8'h00;      memory[40142] <=  8'h00;      memory[40143] <=  8'h00;      memory[40144] <=  8'h00;      memory[40145] <=  8'h00;      memory[40146] <=  8'h00;      memory[40147] <=  8'h00;      memory[40148] <=  8'h00;      memory[40149] <=  8'h00;      memory[40150] <=  8'h00;      memory[40151] <=  8'h00;      memory[40152] <=  8'h00;      memory[40153] <=  8'h00;      memory[40154] <=  8'h00;      memory[40155] <=  8'h00;      memory[40156] <=  8'h00;      memory[40157] <=  8'h00;      memory[40158] <=  8'h00;      memory[40159] <=  8'h00;      memory[40160] <=  8'h00;      memory[40161] <=  8'h00;      memory[40162] <=  8'h00;      memory[40163] <=  8'h00;      memory[40164] <=  8'h00;      memory[40165] <=  8'h00;      memory[40166] <=  8'h00;      memory[40167] <=  8'h00;      memory[40168] <=  8'h00;      memory[40169] <=  8'h00;      memory[40170] <=  8'h00;      memory[40171] <=  8'h00;      memory[40172] <=  8'h00;      memory[40173] <=  8'h00;      memory[40174] <=  8'h00;      memory[40175] <=  8'h00;      memory[40176] <=  8'h00;      memory[40177] <=  8'h00;      memory[40178] <=  8'h00;      memory[40179] <=  8'h00;      memory[40180] <=  8'h00;      memory[40181] <=  8'h00;      memory[40182] <=  8'h00;      memory[40183] <=  8'h00;      memory[40184] <=  8'h00;      memory[40185] <=  8'h00;      memory[40186] <=  8'h00;      memory[40187] <=  8'h00;      memory[40188] <=  8'h00;      memory[40189] <=  8'h00;      memory[40190] <=  8'h00;      memory[40191] <=  8'h00;      memory[40192] <=  8'h00;      memory[40193] <=  8'h00;      memory[40194] <=  8'h00;      memory[40195] <=  8'h00;      memory[40196] <=  8'h00;      memory[40197] <=  8'h00;      memory[40198] <=  8'h00;      memory[40199] <=  8'h00;      memory[40200] <=  8'h00;      memory[40201] <=  8'h00;      memory[40202] <=  8'h00;      memory[40203] <=  8'h00;      memory[40204] <=  8'h00;      memory[40205] <=  8'h00;      memory[40206] <=  8'h00;      memory[40207] <=  8'h00;      memory[40208] <=  8'h00;      memory[40209] <=  8'h00;      memory[40210] <=  8'h00;      memory[40211] <=  8'h00;      memory[40212] <=  8'h00;      memory[40213] <=  8'h00;      memory[40214] <=  8'h00;      memory[40215] <=  8'h00;      memory[40216] <=  8'h00;      memory[40217] <=  8'h00;      memory[40218] <=  8'h00;      memory[40219] <=  8'h00;      memory[40220] <=  8'h00;      memory[40221] <=  8'h00;      memory[40222] <=  8'h00;      memory[40223] <=  8'h00;      memory[40224] <=  8'h00;      memory[40225] <=  8'h00;      memory[40226] <=  8'h00;      memory[40227] <=  8'h00;      memory[40228] <=  8'h00;      memory[40229] <=  8'h00;      memory[40230] <=  8'h00;      memory[40231] <=  8'h00;      memory[40232] <=  8'h00;      memory[40233] <=  8'h00;      memory[40234] <=  8'h00;      memory[40235] <=  8'h00;      memory[40236] <=  8'h00;      memory[40237] <=  8'h00;      memory[40238] <=  8'h00;      memory[40239] <=  8'h00;      memory[40240] <=  8'h00;      memory[40241] <=  8'h00;      memory[40242] <=  8'h00;      memory[40243] <=  8'h00;      memory[40244] <=  8'h00;      memory[40245] <=  8'h00;      memory[40246] <=  8'h00;      memory[40247] <=  8'h00;      memory[40248] <=  8'h00;      memory[40249] <=  8'h00;      memory[40250] <=  8'h00;      memory[40251] <=  8'h00;      memory[40252] <=  8'h00;      memory[40253] <=  8'h00;      memory[40254] <=  8'h00;      memory[40255] <=  8'h00;      memory[40256] <=  8'h00;      memory[40257] <=  8'h00;      memory[40258] <=  8'h00;      memory[40259] <=  8'h00;      memory[40260] <=  8'h00;      memory[40261] <=  8'h00;      memory[40262] <=  8'h00;      memory[40263] <=  8'h00;      memory[40264] <=  8'h00;      memory[40265] <=  8'h00;      memory[40266] <=  8'h00;      memory[40267] <=  8'h00;      memory[40268] <=  8'h00;      memory[40269] <=  8'h00;      memory[40270] <=  8'h00;      memory[40271] <=  8'h00;      memory[40272] <=  8'h00;      memory[40273] <=  8'h00;      memory[40274] <=  8'h00;      memory[40275] <=  8'h00;      memory[40276] <=  8'h00;      memory[40277] <=  8'h00;      memory[40278] <=  8'h00;      memory[40279] <=  8'h00;      memory[40280] <=  8'h00;      memory[40281] <=  8'h00;      memory[40282] <=  8'h00;      memory[40283] <=  8'h00;      memory[40284] <=  8'h00;      memory[40285] <=  8'h00;      memory[40286] <=  8'h00;      memory[40287] <=  8'h00;      memory[40288] <=  8'h00;      memory[40289] <=  8'h00;      memory[40290] <=  8'h00;      memory[40291] <=  8'h00;      memory[40292] <=  8'h00;      memory[40293] <=  8'h00;      memory[40294] <=  8'h00;      memory[40295] <=  8'h00;      memory[40296] <=  8'h00;      memory[40297] <=  8'h00;      memory[40298] <=  8'h00;      memory[40299] <=  8'h00;      memory[40300] <=  8'h00;      memory[40301] <=  8'h00;      memory[40302] <=  8'h00;      memory[40303] <=  8'h00;      memory[40304] <=  8'h00;      memory[40305] <=  8'h00;      memory[40306] <=  8'h00;      memory[40307] <=  8'h00;      memory[40308] <=  8'h00;      memory[40309] <=  8'h00;      memory[40310] <=  8'h00;      memory[40311] <=  8'h00;      memory[40312] <=  8'h00;      memory[40313] <=  8'h00;      memory[40314] <=  8'h00;      memory[40315] <=  8'h00;      memory[40316] <=  8'h00;      memory[40317] <=  8'h00;      memory[40318] <=  8'h00;      memory[40319] <=  8'h00;      memory[40320] <=  8'h00;      memory[40321] <=  8'h00;      memory[40322] <=  8'h00;      memory[40323] <=  8'h00;      memory[40324] <=  8'h00;      memory[40325] <=  8'h00;      memory[40326] <=  8'h00;      memory[40327] <=  8'h00;      memory[40328] <=  8'h00;      memory[40329] <=  8'h00;      memory[40330] <=  8'h00;      memory[40331] <=  8'h00;      memory[40332] <=  8'h00;      memory[40333] <=  8'h00;      memory[40334] <=  8'h00;      memory[40335] <=  8'h00;      memory[40336] <=  8'h00;      memory[40337] <=  8'h00;      memory[40338] <=  8'h00;      memory[40339] <=  8'h00;      memory[40340] <=  8'h00;      memory[40341] <=  8'h00;      memory[40342] <=  8'h00;      memory[40343] <=  8'h00;      memory[40344] <=  8'h00;      memory[40345] <=  8'h00;      memory[40346] <=  8'h00;      memory[40347] <=  8'h00;      memory[40348] <=  8'h00;      memory[40349] <=  8'h00;      memory[40350] <=  8'h00;      memory[40351] <=  8'h00;      memory[40352] <=  8'h00;      memory[40353] <=  8'h00;      memory[40354] <=  8'h00;      memory[40355] <=  8'h00;      memory[40356] <=  8'h00;      memory[40357] <=  8'h00;      memory[40358] <=  8'h00;      memory[40359] <=  8'h00;      memory[40360] <=  8'h00;      memory[40361] <=  8'h00;      memory[40362] <=  8'h00;      memory[40363] <=  8'h00;      memory[40364] <=  8'h00;      memory[40365] <=  8'h00;      memory[40366] <=  8'h00;      memory[40367] <=  8'h00;      memory[40368] <=  8'h00;      memory[40369] <=  8'h00;      memory[40370] <=  8'h00;      memory[40371] <=  8'h00;      memory[40372] <=  8'h00;      memory[40373] <=  8'h00;      memory[40374] <=  8'h00;      memory[40375] <=  8'h00;      memory[40376] <=  8'h00;      memory[40377] <=  8'h00;      memory[40378] <=  8'h00;      memory[40379] <=  8'h00;      memory[40380] <=  8'h00;      memory[40381] <=  8'h00;      memory[40382] <=  8'h00;      memory[40383] <=  8'h00;      memory[40384] <=  8'h00;      memory[40385] <=  8'h00;      memory[40386] <=  8'h00;      memory[40387] <=  8'h00;      memory[40388] <=  8'h00;      memory[40389] <=  8'h00;      memory[40390] <=  8'h00;      memory[40391] <=  8'h00;      memory[40392] <=  8'h00;      memory[40393] <=  8'h00;      memory[40394] <=  8'h00;      memory[40395] <=  8'h00;      memory[40396] <=  8'h00;      memory[40397] <=  8'h00;      memory[40398] <=  8'h00;      memory[40399] <=  8'h00;      memory[40400] <=  8'h00;      memory[40401] <=  8'h00;      memory[40402] <=  8'h00;      memory[40403] <=  8'h00;      memory[40404] <=  8'h00;      memory[40405] <=  8'h00;      memory[40406] <=  8'h00;      memory[40407] <=  8'h00;      memory[40408] <=  8'h00;      memory[40409] <=  8'h00;      memory[40410] <=  8'h00;      memory[40411] <=  8'h00;      memory[40412] <=  8'h00;      memory[40413] <=  8'h00;      memory[40414] <=  8'h00;      memory[40415] <=  8'h00;      memory[40416] <=  8'h00;      memory[40417] <=  8'h00;      memory[40418] <=  8'h00;      memory[40419] <=  8'h00;      memory[40420] <=  8'h00;      memory[40421] <=  8'h00;      memory[40422] <=  8'h00;      memory[40423] <=  8'h00;      memory[40424] <=  8'h00;      memory[40425] <=  8'h00;      memory[40426] <=  8'h00;      memory[40427] <=  8'h00;      memory[40428] <=  8'h00;      memory[40429] <=  8'h00;      memory[40430] <=  8'h00;      memory[40431] <=  8'h00;      memory[40432] <=  8'h00;      memory[40433] <=  8'h00;      memory[40434] <=  8'h00;      memory[40435] <=  8'h00;      memory[40436] <=  8'h00;      memory[40437] <=  8'h00;      memory[40438] <=  8'h00;      memory[40439] <=  8'h00;      memory[40440] <=  8'h00;      memory[40441] <=  8'h00;      memory[40442] <=  8'h00;      memory[40443] <=  8'h00;      memory[40444] <=  8'h00;      memory[40445] <=  8'h00;      memory[40446] <=  8'h00;      memory[40447] <=  8'h00;      memory[40448] <=  8'h00;      memory[40449] <=  8'h00;      memory[40450] <=  8'h00;      memory[40451] <=  8'h00;      memory[40452] <=  8'h00;      memory[40453] <=  8'h00;      memory[40454] <=  8'h00;      memory[40455] <=  8'h00;      memory[40456] <=  8'h00;      memory[40457] <=  8'h00;      memory[40458] <=  8'h00;      memory[40459] <=  8'h00;      memory[40460] <=  8'h00;      memory[40461] <=  8'h00;      memory[40462] <=  8'h00;      memory[40463] <=  8'h00;      memory[40464] <=  8'h00;      memory[40465] <=  8'h00;      memory[40466] <=  8'h00;      memory[40467] <=  8'h00;      memory[40468] <=  8'h00;      memory[40469] <=  8'h00;      memory[40470] <=  8'h00;      memory[40471] <=  8'h00;      memory[40472] <=  8'h00;      memory[40473] <=  8'h00;      memory[40474] <=  8'h00;      memory[40475] <=  8'h00;      memory[40476] <=  8'h00;      memory[40477] <=  8'h00;      memory[40478] <=  8'h00;      memory[40479] <=  8'h00;      memory[40480] <=  8'h00;      memory[40481] <=  8'h00;      memory[40482] <=  8'h00;      memory[40483] <=  8'h00;      memory[40484] <=  8'h00;      memory[40485] <=  8'h00;      memory[40486] <=  8'h00;      memory[40487] <=  8'h00;      memory[40488] <=  8'h00;      memory[40489] <=  8'h00;      memory[40490] <=  8'h00;      memory[40491] <=  8'h00;      memory[40492] <=  8'h00;      memory[40493] <=  8'h00;      memory[40494] <=  8'h00;      memory[40495] <=  8'h00;      memory[40496] <=  8'h00;      memory[40497] <=  8'h00;      memory[40498] <=  8'h00;      memory[40499] <=  8'h00;      memory[40500] <=  8'h00;      memory[40501] <=  8'h00;      memory[40502] <=  8'h00;      memory[40503] <=  8'h00;      memory[40504] <=  8'h00;      memory[40505] <=  8'h00;      memory[40506] <=  8'h00;      memory[40507] <=  8'h00;      memory[40508] <=  8'h00;      memory[40509] <=  8'h00;      memory[40510] <=  8'h00;      memory[40511] <=  8'h00;      memory[40512] <=  8'h00;      memory[40513] <=  8'h00;      memory[40514] <=  8'h00;      memory[40515] <=  8'h00;      memory[40516] <=  8'h00;      memory[40517] <=  8'h00;      memory[40518] <=  8'h00;      memory[40519] <=  8'h00;      memory[40520] <=  8'h00;      memory[40521] <=  8'h00;      memory[40522] <=  8'h00;      memory[40523] <=  8'h00;      memory[40524] <=  8'h00;      memory[40525] <=  8'h00;      memory[40526] <=  8'h00;      memory[40527] <=  8'h00;      memory[40528] <=  8'h00;      memory[40529] <=  8'h00;      memory[40530] <=  8'h00;      memory[40531] <=  8'h00;      memory[40532] <=  8'h00;      memory[40533] <=  8'h00;      memory[40534] <=  8'h00;      memory[40535] <=  8'h00;      memory[40536] <=  8'h00;      memory[40537] <=  8'h00;      memory[40538] <=  8'h00;      memory[40539] <=  8'h00;      memory[40540] <=  8'h00;      memory[40541] <=  8'h00;      memory[40542] <=  8'h00;      memory[40543] <=  8'h00;      memory[40544] <=  8'h00;      memory[40545] <=  8'h00;      memory[40546] <=  8'h00;      memory[40547] <=  8'h00;      memory[40548] <=  8'h00;      memory[40549] <=  8'h00;      memory[40550] <=  8'h00;      memory[40551] <=  8'h00;      memory[40552] <=  8'h00;      memory[40553] <=  8'h00;      memory[40554] <=  8'h00;      memory[40555] <=  8'h00;      memory[40556] <=  8'h00;      memory[40557] <=  8'h00;      memory[40558] <=  8'h00;      memory[40559] <=  8'h00;      memory[40560] <=  8'h00;      memory[40561] <=  8'h00;      memory[40562] <=  8'h00;      memory[40563] <=  8'h00;      memory[40564] <=  8'h00;      memory[40565] <=  8'h00;      memory[40566] <=  8'h00;      memory[40567] <=  8'h00;      memory[40568] <=  8'h00;      memory[40569] <=  8'h00;      memory[40570] <=  8'h00;      memory[40571] <=  8'h00;      memory[40572] <=  8'h00;      memory[40573] <=  8'h00;      memory[40574] <=  8'h00;      memory[40575] <=  8'h00;      memory[40576] <=  8'h00;      memory[40577] <=  8'h00;      memory[40578] <=  8'h00;      memory[40579] <=  8'h00;      memory[40580] <=  8'h00;      memory[40581] <=  8'h00;      memory[40582] <=  8'h00;      memory[40583] <=  8'h00;      memory[40584] <=  8'h00;      memory[40585] <=  8'h00;      memory[40586] <=  8'h00;      memory[40587] <=  8'h00;      memory[40588] <=  8'h00;      memory[40589] <=  8'h00;      memory[40590] <=  8'h00;      memory[40591] <=  8'h00;      memory[40592] <=  8'h00;      memory[40593] <=  8'h00;      memory[40594] <=  8'h00;      memory[40595] <=  8'h00;      memory[40596] <=  8'h00;      memory[40597] <=  8'h00;      memory[40598] <=  8'h00;      memory[40599] <=  8'h00;      memory[40600] <=  8'h00;      memory[40601] <=  8'h00;      memory[40602] <=  8'h00;      memory[40603] <=  8'h00;      memory[40604] <=  8'h00;      memory[40605] <=  8'h00;      memory[40606] <=  8'h00;      memory[40607] <=  8'h00;      memory[40608] <=  8'h00;      memory[40609] <=  8'h00;      memory[40610] <=  8'h00;      memory[40611] <=  8'h00;      memory[40612] <=  8'h00;      memory[40613] <=  8'h00;      memory[40614] <=  8'h00;      memory[40615] <=  8'h00;      memory[40616] <=  8'h00;      memory[40617] <=  8'h00;      memory[40618] <=  8'h00;      memory[40619] <=  8'h00;      memory[40620] <=  8'h00;      memory[40621] <=  8'h00;      memory[40622] <=  8'h00;      memory[40623] <=  8'h00;      memory[40624] <=  8'h00;      memory[40625] <=  8'h00;      memory[40626] <=  8'h00;      memory[40627] <=  8'h00;      memory[40628] <=  8'h00;      memory[40629] <=  8'h00;      memory[40630] <=  8'h00;      memory[40631] <=  8'h00;      memory[40632] <=  8'h00;      memory[40633] <=  8'h00;      memory[40634] <=  8'h00;      memory[40635] <=  8'h00;      memory[40636] <=  8'h00;      memory[40637] <=  8'h00;      memory[40638] <=  8'h00;      memory[40639] <=  8'h00;      memory[40640] <=  8'h00;      memory[40641] <=  8'h00;      memory[40642] <=  8'h00;      memory[40643] <=  8'h00;      memory[40644] <=  8'h00;      memory[40645] <=  8'h00;      memory[40646] <=  8'h00;      memory[40647] <=  8'h00;      memory[40648] <=  8'h00;      memory[40649] <=  8'h00;      memory[40650] <=  8'h00;      memory[40651] <=  8'h00;      memory[40652] <=  8'h00;      memory[40653] <=  8'h00;      memory[40654] <=  8'h00;      memory[40655] <=  8'h00;      memory[40656] <=  8'h00;      memory[40657] <=  8'h00;      memory[40658] <=  8'h00;      memory[40659] <=  8'h00;      memory[40660] <=  8'h00;      memory[40661] <=  8'h00;      memory[40662] <=  8'h00;      memory[40663] <=  8'h00;      memory[40664] <=  8'h00;      memory[40665] <=  8'h00;      memory[40666] <=  8'h00;      memory[40667] <=  8'h00;      memory[40668] <=  8'h00;      memory[40669] <=  8'h00;      memory[40670] <=  8'h00;      memory[40671] <=  8'h00;      memory[40672] <=  8'h00;      memory[40673] <=  8'h00;      memory[40674] <=  8'h00;      memory[40675] <=  8'h00;      memory[40676] <=  8'h00;      memory[40677] <=  8'h00;      memory[40678] <=  8'h00;      memory[40679] <=  8'h00;      memory[40680] <=  8'h00;      memory[40681] <=  8'h00;      memory[40682] <=  8'h00;      memory[40683] <=  8'h00;      memory[40684] <=  8'h00;      memory[40685] <=  8'h00;      memory[40686] <=  8'h00;      memory[40687] <=  8'h00;      memory[40688] <=  8'h00;      memory[40689] <=  8'h00;      memory[40690] <=  8'h00;      memory[40691] <=  8'h00;      memory[40692] <=  8'h00;      memory[40693] <=  8'h00;      memory[40694] <=  8'h00;      memory[40695] <=  8'h00;      memory[40696] <=  8'h00;      memory[40697] <=  8'h00;      memory[40698] <=  8'h00;      memory[40699] <=  8'h00;      memory[40700] <=  8'h00;      memory[40701] <=  8'h00;      memory[40702] <=  8'h00;      memory[40703] <=  8'h00;      memory[40704] <=  8'h00;      memory[40705] <=  8'h00;      memory[40706] <=  8'h00;      memory[40707] <=  8'h00;      memory[40708] <=  8'h00;      memory[40709] <=  8'h00;      memory[40710] <=  8'h00;      memory[40711] <=  8'h00;      memory[40712] <=  8'h00;      memory[40713] <=  8'h00;      memory[40714] <=  8'h00;      memory[40715] <=  8'h00;      memory[40716] <=  8'h00;      memory[40717] <=  8'h00;      memory[40718] <=  8'h00;      memory[40719] <=  8'h00;      memory[40720] <=  8'h00;      memory[40721] <=  8'h00;      memory[40722] <=  8'h00;      memory[40723] <=  8'h00;      memory[40724] <=  8'h00;      memory[40725] <=  8'h00;      memory[40726] <=  8'h00;      memory[40727] <=  8'h00;      memory[40728] <=  8'h00;      memory[40729] <=  8'h00;      memory[40730] <=  8'h00;      memory[40731] <=  8'h00;      memory[40732] <=  8'h00;      memory[40733] <=  8'h00;      memory[40734] <=  8'h00;      memory[40735] <=  8'h00;      memory[40736] <=  8'h00;      memory[40737] <=  8'h00;      memory[40738] <=  8'h00;      memory[40739] <=  8'h00;      memory[40740] <=  8'h00;      memory[40741] <=  8'h00;      memory[40742] <=  8'h00;      memory[40743] <=  8'h00;      memory[40744] <=  8'h00;      memory[40745] <=  8'h00;      memory[40746] <=  8'h00;      memory[40747] <=  8'h00;      memory[40748] <=  8'h00;      memory[40749] <=  8'h00;      memory[40750] <=  8'h00;      memory[40751] <=  8'h00;      memory[40752] <=  8'h00;      memory[40753] <=  8'h00;      memory[40754] <=  8'h00;      memory[40755] <=  8'h00;      memory[40756] <=  8'h00;      memory[40757] <=  8'h00;      memory[40758] <=  8'h00;      memory[40759] <=  8'h00;      memory[40760] <=  8'h00;      memory[40761] <=  8'h00;      memory[40762] <=  8'h00;      memory[40763] <=  8'h00;      memory[40764] <=  8'h00;      memory[40765] <=  8'h00;      memory[40766] <=  8'h00;      memory[40767] <=  8'h00;      memory[40768] <=  8'h00;      memory[40769] <=  8'h00;      memory[40770] <=  8'h00;      memory[40771] <=  8'h00;      memory[40772] <=  8'h00;      memory[40773] <=  8'h00;      memory[40774] <=  8'h00;      memory[40775] <=  8'h00;      memory[40776] <=  8'h00;      memory[40777] <=  8'h00;      memory[40778] <=  8'h00;      memory[40779] <=  8'h00;      memory[40780] <=  8'h00;      memory[40781] <=  8'h00;      memory[40782] <=  8'h00;      memory[40783] <=  8'h00;      memory[40784] <=  8'h00;      memory[40785] <=  8'h00;      memory[40786] <=  8'h00;      memory[40787] <=  8'h00;      memory[40788] <=  8'h00;      memory[40789] <=  8'h00;      memory[40790] <=  8'h00;      memory[40791] <=  8'h00;      memory[40792] <=  8'h00;      memory[40793] <=  8'h00;      memory[40794] <=  8'h00;      memory[40795] <=  8'h00;      memory[40796] <=  8'h00;      memory[40797] <=  8'h00;      memory[40798] <=  8'h00;      memory[40799] <=  8'h00;      memory[40800] <=  8'h00;      memory[40801] <=  8'h00;      memory[40802] <=  8'h00;      memory[40803] <=  8'h00;      memory[40804] <=  8'h00;      memory[40805] <=  8'h00;      memory[40806] <=  8'h00;      memory[40807] <=  8'h00;      memory[40808] <=  8'h00;      memory[40809] <=  8'h00;      memory[40810] <=  8'h00;      memory[40811] <=  8'h00;      memory[40812] <=  8'h00;      memory[40813] <=  8'h00;      memory[40814] <=  8'h00;      memory[40815] <=  8'h00;      memory[40816] <=  8'h00;      memory[40817] <=  8'h00;      memory[40818] <=  8'h00;      memory[40819] <=  8'h00;      memory[40820] <=  8'h00;      memory[40821] <=  8'h00;      memory[40822] <=  8'h00;      memory[40823] <=  8'h00;      memory[40824] <=  8'h00;      memory[40825] <=  8'h00;      memory[40826] <=  8'h00;      memory[40827] <=  8'h00;      memory[40828] <=  8'h00;      memory[40829] <=  8'h00;      memory[40830] <=  8'h00;      memory[40831] <=  8'h00;      memory[40832] <=  8'h00;      memory[40833] <=  8'h00;      memory[40834] <=  8'h00;      memory[40835] <=  8'h00;      memory[40836] <=  8'h00;      memory[40837] <=  8'h00;      memory[40838] <=  8'h00;      memory[40839] <=  8'h00;      memory[40840] <=  8'h00;      memory[40841] <=  8'h00;      memory[40842] <=  8'h00;      memory[40843] <=  8'h00;      memory[40844] <=  8'h00;      memory[40845] <=  8'h00;      memory[40846] <=  8'h00;      memory[40847] <=  8'h00;      memory[40848] <=  8'h00;      memory[40849] <=  8'h00;      memory[40850] <=  8'h00;      memory[40851] <=  8'h00;      memory[40852] <=  8'h00;      memory[40853] <=  8'h00;      memory[40854] <=  8'h00;      memory[40855] <=  8'h00;      memory[40856] <=  8'h00;      memory[40857] <=  8'h00;      memory[40858] <=  8'h00;      memory[40859] <=  8'h00;      memory[40860] <=  8'h00;      memory[40861] <=  8'h00;      memory[40862] <=  8'h00;      memory[40863] <=  8'h00;      memory[40864] <=  8'h00;      memory[40865] <=  8'h00;      memory[40866] <=  8'h00;      memory[40867] <=  8'h00;      memory[40868] <=  8'h00;      memory[40869] <=  8'h00;      memory[40870] <=  8'h00;      memory[40871] <=  8'h00;      memory[40872] <=  8'h00;      memory[40873] <=  8'h00;      memory[40874] <=  8'h00;      memory[40875] <=  8'h00;      memory[40876] <=  8'h00;      memory[40877] <=  8'h00;      memory[40878] <=  8'h00;      memory[40879] <=  8'h00;      memory[40880] <=  8'h00;      memory[40881] <=  8'h00;      memory[40882] <=  8'h00;      memory[40883] <=  8'h00;      memory[40884] <=  8'h00;      memory[40885] <=  8'h00;      memory[40886] <=  8'h00;      memory[40887] <=  8'h00;      memory[40888] <=  8'h00;      memory[40889] <=  8'h00;      memory[40890] <=  8'h00;      memory[40891] <=  8'h00;      memory[40892] <=  8'h00;      memory[40893] <=  8'h00;      memory[40894] <=  8'h00;      memory[40895] <=  8'h00;      memory[40896] <=  8'h00;      memory[40897] <=  8'h00;      memory[40898] <=  8'h00;      memory[40899] <=  8'h00;      memory[40900] <=  8'h00;      memory[40901] <=  8'h00;      memory[40902] <=  8'h00;      memory[40903] <=  8'h00;      memory[40904] <=  8'h00;      memory[40905] <=  8'h00;      memory[40906] <=  8'h00;      memory[40907] <=  8'h00;      memory[40908] <=  8'h00;      memory[40909] <=  8'h00;      memory[40910] <=  8'h00;      memory[40911] <=  8'h00;      memory[40912] <=  8'h00;      memory[40913] <=  8'h00;      memory[40914] <=  8'h00;      memory[40915] <=  8'h00;      memory[40916] <=  8'h00;      memory[40917] <=  8'h00;      memory[40918] <=  8'h00;      memory[40919] <=  8'h00;      memory[40920] <=  8'h00;      memory[40921] <=  8'h00;      memory[40922] <=  8'h00;      memory[40923] <=  8'h00;      memory[40924] <=  8'h00;      memory[40925] <=  8'h00;      memory[40926] <=  8'h00;      memory[40927] <=  8'h00;      memory[40928] <=  8'h00;      memory[40929] <=  8'h00;      memory[40930] <=  8'h00;      memory[40931] <=  8'h00;      memory[40932] <=  8'h00;      memory[40933] <=  8'h00;      memory[40934] <=  8'h00;      memory[40935] <=  8'h00;      memory[40936] <=  8'h00;      memory[40937] <=  8'h00;      memory[40938] <=  8'h00;      memory[40939] <=  8'h00;      memory[40940] <=  8'h00;      memory[40941] <=  8'h00;      memory[40942] <=  8'h00;      memory[40943] <=  8'h00;      memory[40944] <=  8'h00;      memory[40945] <=  8'h00;      memory[40946] <=  8'h00;      memory[40947] <=  8'h00;      memory[40948] <=  8'h00;      memory[40949] <=  8'h00;      memory[40950] <=  8'h00;      memory[40951] <=  8'h00;      memory[40952] <=  8'h00;      memory[40953] <=  8'h00;      memory[40954] <=  8'h00;      memory[40955] <=  8'h00;      memory[40956] <=  8'h00;      memory[40957] <=  8'h00;      memory[40958] <=  8'h00;      memory[40959] <=  8'h00;      memory[40960] <=  8'h00;      memory[40961] <=  8'h00;      memory[40962] <=  8'h00;      memory[40963] <=  8'h00;      memory[40964] <=  8'h00;      memory[40965] <=  8'h00;      memory[40966] <=  8'h00;      memory[40967] <=  8'h00;      memory[40968] <=  8'h00;      memory[40969] <=  8'h00;      memory[40970] <=  8'h00;      memory[40971] <=  8'h00;      memory[40972] <=  8'h00;      memory[40973] <=  8'h00;      memory[40974] <=  8'h00;      memory[40975] <=  8'h00;      memory[40976] <=  8'h00;      memory[40977] <=  8'h00;      memory[40978] <=  8'h00;      memory[40979] <=  8'h00;      memory[40980] <=  8'h00;      memory[40981] <=  8'h00;      memory[40982] <=  8'h00;      memory[40983] <=  8'h00;      memory[40984] <=  8'h00;      memory[40985] <=  8'h00;      memory[40986] <=  8'h00;      memory[40987] <=  8'h00;      memory[40988] <=  8'h00;      memory[40989] <=  8'h00;      memory[40990] <=  8'h00;      memory[40991] <=  8'h00;      memory[40992] <=  8'h00;      memory[40993] <=  8'h00;      memory[40994] <=  8'h00;      memory[40995] <=  8'h00;      memory[40996] <=  8'h00;      memory[40997] <=  8'h00;      memory[40998] <=  8'h00;      memory[40999] <=  8'h00;      memory[41000] <=  8'h00;      memory[41001] <=  8'h00;      memory[41002] <=  8'h00;      memory[41003] <=  8'h00;      memory[41004] <=  8'h00;      memory[41005] <=  8'h00;      memory[41006] <=  8'h00;      memory[41007] <=  8'h00;      memory[41008] <=  8'h00;      memory[41009] <=  8'h00;      memory[41010] <=  8'h00;      memory[41011] <=  8'h00;      memory[41012] <=  8'h00;      memory[41013] <=  8'h00;      memory[41014] <=  8'h00;      memory[41015] <=  8'h00;      memory[41016] <=  8'h00;      memory[41017] <=  8'h00;      memory[41018] <=  8'h00;      memory[41019] <=  8'h00;      memory[41020] <=  8'h00;      memory[41021] <=  8'h00;      memory[41022] <=  8'h00;      memory[41023] <=  8'h00;      memory[41024] <=  8'h00;      memory[41025] <=  8'h00;      memory[41026] <=  8'h00;      memory[41027] <=  8'h00;      memory[41028] <=  8'h00;      memory[41029] <=  8'h00;      memory[41030] <=  8'h00;      memory[41031] <=  8'h00;      memory[41032] <=  8'h00;      memory[41033] <=  8'h00;      memory[41034] <=  8'h00;      memory[41035] <=  8'h00;      memory[41036] <=  8'h00;      memory[41037] <=  8'h00;      memory[41038] <=  8'h00;      memory[41039] <=  8'h00;      memory[41040] <=  8'h00;      memory[41041] <=  8'h00;      memory[41042] <=  8'h00;      memory[41043] <=  8'h00;      memory[41044] <=  8'h00;      memory[41045] <=  8'h00;      memory[41046] <=  8'h00;      memory[41047] <=  8'h00;      memory[41048] <=  8'h00;      memory[41049] <=  8'h00;      memory[41050] <=  8'h00;      memory[41051] <=  8'h00;      memory[41052] <=  8'h00;      memory[41053] <=  8'h00;      memory[41054] <=  8'h00;      memory[41055] <=  8'h00;      memory[41056] <=  8'h00;      memory[41057] <=  8'h00;      memory[41058] <=  8'h00;      memory[41059] <=  8'h00;      memory[41060] <=  8'h00;      memory[41061] <=  8'h00;      memory[41062] <=  8'h00;      memory[41063] <=  8'h00;      memory[41064] <=  8'h00;      memory[41065] <=  8'h00;      memory[41066] <=  8'h00;      memory[41067] <=  8'h00;      memory[41068] <=  8'h00;      memory[41069] <=  8'h00;      memory[41070] <=  8'h00;      memory[41071] <=  8'h00;      memory[41072] <=  8'h00;      memory[41073] <=  8'h00;      memory[41074] <=  8'h00;      memory[41075] <=  8'h00;      memory[41076] <=  8'h00;      memory[41077] <=  8'h00;      memory[41078] <=  8'h00;      memory[41079] <=  8'h00;      memory[41080] <=  8'h00;      memory[41081] <=  8'h00;      memory[41082] <=  8'h00;      memory[41083] <=  8'h00;      memory[41084] <=  8'h00;      memory[41085] <=  8'h00;      memory[41086] <=  8'h00;      memory[41087] <=  8'h00;      memory[41088] <=  8'h00;      memory[41089] <=  8'h00;      memory[41090] <=  8'h00;      memory[41091] <=  8'h00;      memory[41092] <=  8'h00;      memory[41093] <=  8'h00;      memory[41094] <=  8'h00;      memory[41095] <=  8'h00;      memory[41096] <=  8'h00;      memory[41097] <=  8'h00;      memory[41098] <=  8'h00;      memory[41099] <=  8'h00;      memory[41100] <=  8'h00;      memory[41101] <=  8'h00;      memory[41102] <=  8'h00;      memory[41103] <=  8'h00;      memory[41104] <=  8'h00;      memory[41105] <=  8'h00;      memory[41106] <=  8'h00;      memory[41107] <=  8'h00;      memory[41108] <=  8'h00;      memory[41109] <=  8'h00;      memory[41110] <=  8'h00;      memory[41111] <=  8'h00;      memory[41112] <=  8'h00;      memory[41113] <=  8'h00;      memory[41114] <=  8'h00;      memory[41115] <=  8'h00;      memory[41116] <=  8'h00;      memory[41117] <=  8'h00;      memory[41118] <=  8'h00;      memory[41119] <=  8'h00;      memory[41120] <=  8'h00;      memory[41121] <=  8'h00;      memory[41122] <=  8'h00;      memory[41123] <=  8'h00;      memory[41124] <=  8'h00;      memory[41125] <=  8'h00;      memory[41126] <=  8'h00;      memory[41127] <=  8'h00;      memory[41128] <=  8'h00;      memory[41129] <=  8'h00;      memory[41130] <=  8'h00;      memory[41131] <=  8'h00;      memory[41132] <=  8'h00;      memory[41133] <=  8'h00;      memory[41134] <=  8'h00;      memory[41135] <=  8'h00;      memory[41136] <=  8'h00;      memory[41137] <=  8'h00;      memory[41138] <=  8'h00;      memory[41139] <=  8'h00;      memory[41140] <=  8'h00;      memory[41141] <=  8'h00;      memory[41142] <=  8'h00;      memory[41143] <=  8'h00;      memory[41144] <=  8'h00;      memory[41145] <=  8'h00;      memory[41146] <=  8'h00;      memory[41147] <=  8'h00;      memory[41148] <=  8'h00;      memory[41149] <=  8'h00;      memory[41150] <=  8'h00;      memory[41151] <=  8'h00;      memory[41152] <=  8'h00;      memory[41153] <=  8'h00;      memory[41154] <=  8'h00;      memory[41155] <=  8'h00;      memory[41156] <=  8'h00;      memory[41157] <=  8'h00;      memory[41158] <=  8'h00;      memory[41159] <=  8'h00;      memory[41160] <=  8'h00;      memory[41161] <=  8'h00;      memory[41162] <=  8'h00;      memory[41163] <=  8'h00;      memory[41164] <=  8'h00;      memory[41165] <=  8'h00;      memory[41166] <=  8'h00;      memory[41167] <=  8'h00;      memory[41168] <=  8'h00;      memory[41169] <=  8'h00;      memory[41170] <=  8'h00;      memory[41171] <=  8'h00;      memory[41172] <=  8'h00;      memory[41173] <=  8'h00;      memory[41174] <=  8'h00;      memory[41175] <=  8'h00;      memory[41176] <=  8'h00;      memory[41177] <=  8'h00;      memory[41178] <=  8'h00;      memory[41179] <=  8'h00;      memory[41180] <=  8'h00;      memory[41181] <=  8'h00;      memory[41182] <=  8'h00;      memory[41183] <=  8'h00;      memory[41184] <=  8'h00;      memory[41185] <=  8'h00;      memory[41186] <=  8'h00;      memory[41187] <=  8'h00;      memory[41188] <=  8'h00;      memory[41189] <=  8'h00;      memory[41190] <=  8'h00;      memory[41191] <=  8'h00;      memory[41192] <=  8'h00;      memory[41193] <=  8'h00;      memory[41194] <=  8'h00;      memory[41195] <=  8'h00;      memory[41196] <=  8'h00;      memory[41197] <=  8'h00;      memory[41198] <=  8'h00;      memory[41199] <=  8'h00;      memory[41200] <=  8'h00;      memory[41201] <=  8'h00;      memory[41202] <=  8'h00;      memory[41203] <=  8'h00;      memory[41204] <=  8'h00;      memory[41205] <=  8'h00;      memory[41206] <=  8'h00;      memory[41207] <=  8'h00;      memory[41208] <=  8'h00;      memory[41209] <=  8'h00;      memory[41210] <=  8'h00;      memory[41211] <=  8'h00;      memory[41212] <=  8'h00;      memory[41213] <=  8'h00;      memory[41214] <=  8'h00;      memory[41215] <=  8'h00;      memory[41216] <=  8'h00;      memory[41217] <=  8'h00;      memory[41218] <=  8'h00;      memory[41219] <=  8'h00;      memory[41220] <=  8'h00;      memory[41221] <=  8'h00;      memory[41222] <=  8'h00;      memory[41223] <=  8'h00;      memory[41224] <=  8'h00;      memory[41225] <=  8'h00;      memory[41226] <=  8'h00;      memory[41227] <=  8'h00;      memory[41228] <=  8'h00;      memory[41229] <=  8'h00;      memory[41230] <=  8'h00;      memory[41231] <=  8'h00;      memory[41232] <=  8'h00;      memory[41233] <=  8'h00;      memory[41234] <=  8'h00;      memory[41235] <=  8'h00;      memory[41236] <=  8'h00;      memory[41237] <=  8'h00;      memory[41238] <=  8'h00;      memory[41239] <=  8'h00;      memory[41240] <=  8'h00;      memory[41241] <=  8'h00;      memory[41242] <=  8'h00;      memory[41243] <=  8'h00;      memory[41244] <=  8'h00;      memory[41245] <=  8'h00;      memory[41246] <=  8'h00;      memory[41247] <=  8'h00;      memory[41248] <=  8'h00;      memory[41249] <=  8'h00;      memory[41250] <=  8'h00;      memory[41251] <=  8'h00;      memory[41252] <=  8'h00;      memory[41253] <=  8'h00;      memory[41254] <=  8'h00;      memory[41255] <=  8'h00;      memory[41256] <=  8'h00;      memory[41257] <=  8'h00;      memory[41258] <=  8'h00;      memory[41259] <=  8'h00;      memory[41260] <=  8'h00;      memory[41261] <=  8'h00;      memory[41262] <=  8'h00;      memory[41263] <=  8'h00;      memory[41264] <=  8'h00;      memory[41265] <=  8'h00;      memory[41266] <=  8'h00;      memory[41267] <=  8'h00;      memory[41268] <=  8'h00;      memory[41269] <=  8'h00;      memory[41270] <=  8'h00;      memory[41271] <=  8'h00;      memory[41272] <=  8'h00;      memory[41273] <=  8'h00;      memory[41274] <=  8'h00;      memory[41275] <=  8'h00;      memory[41276] <=  8'h00;      memory[41277] <=  8'h00;      memory[41278] <=  8'h00;      memory[41279] <=  8'h00;      memory[41280] <=  8'h00;      memory[41281] <=  8'h00;      memory[41282] <=  8'h00;      memory[41283] <=  8'h00;      memory[41284] <=  8'h00;      memory[41285] <=  8'h00;      memory[41286] <=  8'h00;      memory[41287] <=  8'h00;      memory[41288] <=  8'h00;      memory[41289] <=  8'h00;      memory[41290] <=  8'h00;      memory[41291] <=  8'h00;      memory[41292] <=  8'h00;      memory[41293] <=  8'h00;      memory[41294] <=  8'h00;      memory[41295] <=  8'h00;      memory[41296] <=  8'h00;      memory[41297] <=  8'h00;      memory[41298] <=  8'h00;      memory[41299] <=  8'h00;      memory[41300] <=  8'h00;      memory[41301] <=  8'h00;      memory[41302] <=  8'h00;      memory[41303] <=  8'h00;      memory[41304] <=  8'h00;      memory[41305] <=  8'h00;      memory[41306] <=  8'h00;      memory[41307] <=  8'h00;      memory[41308] <=  8'h00;      memory[41309] <=  8'h00;      memory[41310] <=  8'h00;      memory[41311] <=  8'h00;      memory[41312] <=  8'h00;      memory[41313] <=  8'h00;      memory[41314] <=  8'h00;      memory[41315] <=  8'h00;      memory[41316] <=  8'h00;      memory[41317] <=  8'h00;      memory[41318] <=  8'h00;      memory[41319] <=  8'h00;      memory[41320] <=  8'h00;      memory[41321] <=  8'h00;      memory[41322] <=  8'h00;      memory[41323] <=  8'h00;      memory[41324] <=  8'h00;      memory[41325] <=  8'h00;      memory[41326] <=  8'h00;      memory[41327] <=  8'h00;      memory[41328] <=  8'h00;      memory[41329] <=  8'h00;      memory[41330] <=  8'h00;      memory[41331] <=  8'h00;      memory[41332] <=  8'h00;      memory[41333] <=  8'h00;      memory[41334] <=  8'h00;      memory[41335] <=  8'h00;      memory[41336] <=  8'h00;      memory[41337] <=  8'h00;      memory[41338] <=  8'h00;      memory[41339] <=  8'h00;      memory[41340] <=  8'h00;      memory[41341] <=  8'h00;      memory[41342] <=  8'h00;      memory[41343] <=  8'h00;      memory[41344] <=  8'h00;      memory[41345] <=  8'h00;      memory[41346] <=  8'h00;      memory[41347] <=  8'h00;      memory[41348] <=  8'h00;      memory[41349] <=  8'h00;      memory[41350] <=  8'h00;      memory[41351] <=  8'h00;      memory[41352] <=  8'h00;      memory[41353] <=  8'h00;      memory[41354] <=  8'h00;      memory[41355] <=  8'h00;      memory[41356] <=  8'h00;      memory[41357] <=  8'h00;      memory[41358] <=  8'h00;      memory[41359] <=  8'h00;      memory[41360] <=  8'h00;      memory[41361] <=  8'h00;      memory[41362] <=  8'h00;      memory[41363] <=  8'h00;      memory[41364] <=  8'h00;      memory[41365] <=  8'h00;      memory[41366] <=  8'h00;      memory[41367] <=  8'h00;      memory[41368] <=  8'h00;      memory[41369] <=  8'h00;      memory[41370] <=  8'h00;      memory[41371] <=  8'h00;      memory[41372] <=  8'h00;      memory[41373] <=  8'h00;      memory[41374] <=  8'h00;      memory[41375] <=  8'h00;      memory[41376] <=  8'h00;      memory[41377] <=  8'h00;      memory[41378] <=  8'h00;      memory[41379] <=  8'h00;      memory[41380] <=  8'h00;      memory[41381] <=  8'h00;      memory[41382] <=  8'h00;      memory[41383] <=  8'h00;      memory[41384] <=  8'h00;      memory[41385] <=  8'h00;      memory[41386] <=  8'h00;      memory[41387] <=  8'h00;      memory[41388] <=  8'h00;      memory[41389] <=  8'h00;      memory[41390] <=  8'h00;      memory[41391] <=  8'h00;      memory[41392] <=  8'h00;      memory[41393] <=  8'h00;      memory[41394] <=  8'h00;      memory[41395] <=  8'h00;      memory[41396] <=  8'h00;      memory[41397] <=  8'h00;      memory[41398] <=  8'h00;      memory[41399] <=  8'h00;      memory[41400] <=  8'h00;      memory[41401] <=  8'h00;      memory[41402] <=  8'h00;      memory[41403] <=  8'h00;      memory[41404] <=  8'h00;      memory[41405] <=  8'h00;      memory[41406] <=  8'h00;      memory[41407] <=  8'h00;      memory[41408] <=  8'h00;      memory[41409] <=  8'h00;      memory[41410] <=  8'h00;      memory[41411] <=  8'h00;      memory[41412] <=  8'h00;      memory[41413] <=  8'h00;      memory[41414] <=  8'h00;      memory[41415] <=  8'h00;      memory[41416] <=  8'h00;      memory[41417] <=  8'h00;      memory[41418] <=  8'h00;      memory[41419] <=  8'h00;      memory[41420] <=  8'h00;      memory[41421] <=  8'h00;      memory[41422] <=  8'h00;      memory[41423] <=  8'h00;      memory[41424] <=  8'h00;      memory[41425] <=  8'h00;      memory[41426] <=  8'h00;      memory[41427] <=  8'h00;      memory[41428] <=  8'h00;      memory[41429] <=  8'h00;      memory[41430] <=  8'h00;      memory[41431] <=  8'h00;      memory[41432] <=  8'h00;      memory[41433] <=  8'h00;      memory[41434] <=  8'h00;      memory[41435] <=  8'h00;      memory[41436] <=  8'h00;      memory[41437] <=  8'h00;      memory[41438] <=  8'h00;      memory[41439] <=  8'h00;      memory[41440] <=  8'h00;      memory[41441] <=  8'h00;      memory[41442] <=  8'h00;      memory[41443] <=  8'h00;      memory[41444] <=  8'h00;      memory[41445] <=  8'h00;      memory[41446] <=  8'h00;      memory[41447] <=  8'h00;      memory[41448] <=  8'h00;      memory[41449] <=  8'h00;      memory[41450] <=  8'h00;      memory[41451] <=  8'h00;      memory[41452] <=  8'h00;      memory[41453] <=  8'h00;      memory[41454] <=  8'h00;      memory[41455] <=  8'h00;      memory[41456] <=  8'h00;      memory[41457] <=  8'h00;      memory[41458] <=  8'h00;      memory[41459] <=  8'h00;      memory[41460] <=  8'h00;      memory[41461] <=  8'h00;      memory[41462] <=  8'h00;      memory[41463] <=  8'h00;      memory[41464] <=  8'h00;      memory[41465] <=  8'h00;      memory[41466] <=  8'h00;      memory[41467] <=  8'h00;      memory[41468] <=  8'h00;      memory[41469] <=  8'h00;      memory[41470] <=  8'h00;      memory[41471] <=  8'h00;      memory[41472] <=  8'h00;      memory[41473] <=  8'h00;      memory[41474] <=  8'h00;      memory[41475] <=  8'h00;      memory[41476] <=  8'h00;      memory[41477] <=  8'h00;      memory[41478] <=  8'h00;      memory[41479] <=  8'h00;      memory[41480] <=  8'h00;      memory[41481] <=  8'h00;      memory[41482] <=  8'h00;      memory[41483] <=  8'h00;      memory[41484] <=  8'h00;      memory[41485] <=  8'h00;      memory[41486] <=  8'h00;      memory[41487] <=  8'h00;      memory[41488] <=  8'h00;      memory[41489] <=  8'h00;      memory[41490] <=  8'h00;      memory[41491] <=  8'h00;      memory[41492] <=  8'h00;      memory[41493] <=  8'h00;      memory[41494] <=  8'h00;      memory[41495] <=  8'h00;      memory[41496] <=  8'h00;      memory[41497] <=  8'h00;      memory[41498] <=  8'h00;      memory[41499] <=  8'h00;      memory[41500] <=  8'h00;      memory[41501] <=  8'h00;      memory[41502] <=  8'h00;      memory[41503] <=  8'h00;      memory[41504] <=  8'h00;      memory[41505] <=  8'h00;      memory[41506] <=  8'h00;      memory[41507] <=  8'h00;      memory[41508] <=  8'h00;      memory[41509] <=  8'h00;      memory[41510] <=  8'h00;      memory[41511] <=  8'h00;      memory[41512] <=  8'h00;      memory[41513] <=  8'h00;      memory[41514] <=  8'h00;      memory[41515] <=  8'h00;      memory[41516] <=  8'h00;      memory[41517] <=  8'h00;      memory[41518] <=  8'h00;      memory[41519] <=  8'h00;      memory[41520] <=  8'h00;      memory[41521] <=  8'h00;      memory[41522] <=  8'h00;      memory[41523] <=  8'h00;      memory[41524] <=  8'h00;      memory[41525] <=  8'h00;      memory[41526] <=  8'h00;      memory[41527] <=  8'h00;      memory[41528] <=  8'h00;      memory[41529] <=  8'h00;      memory[41530] <=  8'h00;      memory[41531] <=  8'h00;      memory[41532] <=  8'h00;      memory[41533] <=  8'h00;      memory[41534] <=  8'h00;      memory[41535] <=  8'h00;      memory[41536] <=  8'h00;      memory[41537] <=  8'h00;      memory[41538] <=  8'h00;      memory[41539] <=  8'h00;      memory[41540] <=  8'h00;      memory[41541] <=  8'h00;      memory[41542] <=  8'h00;      memory[41543] <=  8'h00;      memory[41544] <=  8'h00;      memory[41545] <=  8'h00;      memory[41546] <=  8'h00;      memory[41547] <=  8'h00;      memory[41548] <=  8'h00;      memory[41549] <=  8'h00;      memory[41550] <=  8'h00;      memory[41551] <=  8'h00;      memory[41552] <=  8'h00;      memory[41553] <=  8'h00;      memory[41554] <=  8'h00;      memory[41555] <=  8'h00;      memory[41556] <=  8'h00;      memory[41557] <=  8'h00;      memory[41558] <=  8'h00;      memory[41559] <=  8'h00;      memory[41560] <=  8'h00;      memory[41561] <=  8'h00;      memory[41562] <=  8'h00;      memory[41563] <=  8'h00;      memory[41564] <=  8'h00;      memory[41565] <=  8'h00;      memory[41566] <=  8'h00;      memory[41567] <=  8'h00;      memory[41568] <=  8'h00;      memory[41569] <=  8'h00;      memory[41570] <=  8'h00;      memory[41571] <=  8'h00;      memory[41572] <=  8'h00;      memory[41573] <=  8'h00;      memory[41574] <=  8'h00;      memory[41575] <=  8'h00;      memory[41576] <=  8'h00;      memory[41577] <=  8'h00;      memory[41578] <=  8'h00;      memory[41579] <=  8'h00;      memory[41580] <=  8'h00;      memory[41581] <=  8'h00;      memory[41582] <=  8'h00;      memory[41583] <=  8'h00;      memory[41584] <=  8'h00;      memory[41585] <=  8'h00;      memory[41586] <=  8'h00;      memory[41587] <=  8'h00;      memory[41588] <=  8'h00;      memory[41589] <=  8'h00;      memory[41590] <=  8'h00;      memory[41591] <=  8'h00;      memory[41592] <=  8'h00;      memory[41593] <=  8'h00;      memory[41594] <=  8'h00;      memory[41595] <=  8'h00;      memory[41596] <=  8'h00;      memory[41597] <=  8'h00;      memory[41598] <=  8'h00;      memory[41599] <=  8'h00;      memory[41600] <=  8'h00;      memory[41601] <=  8'h00;      memory[41602] <=  8'h00;      memory[41603] <=  8'h00;      memory[41604] <=  8'h00;      memory[41605] <=  8'h00;      memory[41606] <=  8'h00;      memory[41607] <=  8'h00;      memory[41608] <=  8'h00;      memory[41609] <=  8'h00;      memory[41610] <=  8'h00;      memory[41611] <=  8'h00;      memory[41612] <=  8'h00;      memory[41613] <=  8'h00;      memory[41614] <=  8'h00;      memory[41615] <=  8'h00;      memory[41616] <=  8'h00;      memory[41617] <=  8'h00;      memory[41618] <=  8'h00;      memory[41619] <=  8'h00;      memory[41620] <=  8'h00;      memory[41621] <=  8'h00;      memory[41622] <=  8'h00;      memory[41623] <=  8'h00;      memory[41624] <=  8'h00;      memory[41625] <=  8'h00;      memory[41626] <=  8'h00;      memory[41627] <=  8'h00;      memory[41628] <=  8'h00;      memory[41629] <=  8'h00;      memory[41630] <=  8'h00;      memory[41631] <=  8'h00;      memory[41632] <=  8'h00;      memory[41633] <=  8'h00;      memory[41634] <=  8'h00;      memory[41635] <=  8'h00;      memory[41636] <=  8'h00;      memory[41637] <=  8'h00;      memory[41638] <=  8'h00;      memory[41639] <=  8'h00;      memory[41640] <=  8'h00;      memory[41641] <=  8'h00;      memory[41642] <=  8'h00;      memory[41643] <=  8'h00;      memory[41644] <=  8'h00;      memory[41645] <=  8'h00;      memory[41646] <=  8'h00;      memory[41647] <=  8'h00;      memory[41648] <=  8'h00;      memory[41649] <=  8'h00;      memory[41650] <=  8'h00;      memory[41651] <=  8'h00;      memory[41652] <=  8'h00;      memory[41653] <=  8'h00;      memory[41654] <=  8'h00;      memory[41655] <=  8'h00;      memory[41656] <=  8'h00;      memory[41657] <=  8'h00;      memory[41658] <=  8'h00;      memory[41659] <=  8'h00;      memory[41660] <=  8'h00;      memory[41661] <=  8'h00;      memory[41662] <=  8'h00;      memory[41663] <=  8'h00;      memory[41664] <=  8'h00;      memory[41665] <=  8'h00;      memory[41666] <=  8'h00;      memory[41667] <=  8'h00;      memory[41668] <=  8'h00;      memory[41669] <=  8'h00;      memory[41670] <=  8'h00;      memory[41671] <=  8'h00;      memory[41672] <=  8'h00;      memory[41673] <=  8'h00;      memory[41674] <=  8'h00;      memory[41675] <=  8'h00;      memory[41676] <=  8'h00;      memory[41677] <=  8'h00;      memory[41678] <=  8'h00;      memory[41679] <=  8'h00;      memory[41680] <=  8'h00;      memory[41681] <=  8'h00;      memory[41682] <=  8'h00;      memory[41683] <=  8'h00;      memory[41684] <=  8'h00;      memory[41685] <=  8'h00;      memory[41686] <=  8'h00;      memory[41687] <=  8'h00;      memory[41688] <=  8'h00;      memory[41689] <=  8'h00;      memory[41690] <=  8'h00;      memory[41691] <=  8'h00;      memory[41692] <=  8'h00;      memory[41693] <=  8'h00;      memory[41694] <=  8'h00;      memory[41695] <=  8'h00;      memory[41696] <=  8'h00;      memory[41697] <=  8'h00;      memory[41698] <=  8'h00;      memory[41699] <=  8'h00;      memory[41700] <=  8'h00;      memory[41701] <=  8'h00;      memory[41702] <=  8'h00;      memory[41703] <=  8'h00;      memory[41704] <=  8'h00;      memory[41705] <=  8'h00;      memory[41706] <=  8'h00;      memory[41707] <=  8'h00;      memory[41708] <=  8'h00;      memory[41709] <=  8'h00;      memory[41710] <=  8'h00;      memory[41711] <=  8'h00;      memory[41712] <=  8'h00;      memory[41713] <=  8'h00;      memory[41714] <=  8'h00;      memory[41715] <=  8'h00;      memory[41716] <=  8'h00;      memory[41717] <=  8'h00;      memory[41718] <=  8'h00;      memory[41719] <=  8'h00;      memory[41720] <=  8'h00;      memory[41721] <=  8'h00;      memory[41722] <=  8'h00;      memory[41723] <=  8'h00;      memory[41724] <=  8'h00;      memory[41725] <=  8'h00;      memory[41726] <=  8'h00;      memory[41727] <=  8'h00;      memory[41728] <=  8'h00;      memory[41729] <=  8'h00;      memory[41730] <=  8'h00;      memory[41731] <=  8'h00;      memory[41732] <=  8'h00;      memory[41733] <=  8'h00;      memory[41734] <=  8'h00;      memory[41735] <=  8'h00;      memory[41736] <=  8'h00;      memory[41737] <=  8'h00;      memory[41738] <=  8'h00;      memory[41739] <=  8'h00;      memory[41740] <=  8'h00;      memory[41741] <=  8'h00;      memory[41742] <=  8'h00;      memory[41743] <=  8'h00;      memory[41744] <=  8'h00;      memory[41745] <=  8'h00;      memory[41746] <=  8'h00;      memory[41747] <=  8'h00;      memory[41748] <=  8'h00;      memory[41749] <=  8'h00;      memory[41750] <=  8'h00;      memory[41751] <=  8'h00;      memory[41752] <=  8'h00;      memory[41753] <=  8'h00;      memory[41754] <=  8'h00;      memory[41755] <=  8'h00;      memory[41756] <=  8'h00;      memory[41757] <=  8'h00;      memory[41758] <=  8'h00;      memory[41759] <=  8'h00;      memory[41760] <=  8'h00;      memory[41761] <=  8'h00;      memory[41762] <=  8'h00;      memory[41763] <=  8'h00;      memory[41764] <=  8'h00;      memory[41765] <=  8'h00;      memory[41766] <=  8'h00;      memory[41767] <=  8'h00;      memory[41768] <=  8'h00;      memory[41769] <=  8'h00;      memory[41770] <=  8'h00;      memory[41771] <=  8'h00;      memory[41772] <=  8'h00;      memory[41773] <=  8'h00;      memory[41774] <=  8'h00;      memory[41775] <=  8'h00;      memory[41776] <=  8'h00;      memory[41777] <=  8'h00;      memory[41778] <=  8'h00;      memory[41779] <=  8'h00;      memory[41780] <=  8'h00;      memory[41781] <=  8'h00;      memory[41782] <=  8'h00;      memory[41783] <=  8'h00;      memory[41784] <=  8'h00;      memory[41785] <=  8'h00;      memory[41786] <=  8'h00;      memory[41787] <=  8'h00;      memory[41788] <=  8'h00;      memory[41789] <=  8'h00;      memory[41790] <=  8'h00;      memory[41791] <=  8'h00;      memory[41792] <=  8'h00;      memory[41793] <=  8'h00;      memory[41794] <=  8'h00;      memory[41795] <=  8'h00;      memory[41796] <=  8'h00;      memory[41797] <=  8'h00;      memory[41798] <=  8'h00;      memory[41799] <=  8'h00;      memory[41800] <=  8'h00;      memory[41801] <=  8'h00;      memory[41802] <=  8'h00;      memory[41803] <=  8'h00;      memory[41804] <=  8'h00;      memory[41805] <=  8'h00;      memory[41806] <=  8'h00;      memory[41807] <=  8'h00;      memory[41808] <=  8'h00;      memory[41809] <=  8'h00;      memory[41810] <=  8'h00;      memory[41811] <=  8'h00;      memory[41812] <=  8'h00;      memory[41813] <=  8'h00;      memory[41814] <=  8'h00;      memory[41815] <=  8'h00;      memory[41816] <=  8'h00;      memory[41817] <=  8'h00;      memory[41818] <=  8'h00;      memory[41819] <=  8'h00;      memory[41820] <=  8'h00;      memory[41821] <=  8'h00;      memory[41822] <=  8'h00;      memory[41823] <=  8'h00;      memory[41824] <=  8'h00;      memory[41825] <=  8'h00;      memory[41826] <=  8'h00;      memory[41827] <=  8'h00;      memory[41828] <=  8'h00;      memory[41829] <=  8'h00;      memory[41830] <=  8'h00;      memory[41831] <=  8'h00;      memory[41832] <=  8'h00;      memory[41833] <=  8'h00;      memory[41834] <=  8'h00;      memory[41835] <=  8'h00;      memory[41836] <=  8'h00;      memory[41837] <=  8'h00;      memory[41838] <=  8'h00;      memory[41839] <=  8'h00;      memory[41840] <=  8'h00;      memory[41841] <=  8'h00;      memory[41842] <=  8'h00;      memory[41843] <=  8'h00;      memory[41844] <=  8'h00;      memory[41845] <=  8'h00;      memory[41846] <=  8'h00;      memory[41847] <=  8'h00;      memory[41848] <=  8'h00;      memory[41849] <=  8'h00;      memory[41850] <=  8'h00;      memory[41851] <=  8'h00;      memory[41852] <=  8'h00;      memory[41853] <=  8'h00;      memory[41854] <=  8'h00;      memory[41855] <=  8'h00;      memory[41856] <=  8'h00;      memory[41857] <=  8'h00;      memory[41858] <=  8'h00;      memory[41859] <=  8'h00;      memory[41860] <=  8'h00;      memory[41861] <=  8'h00;      memory[41862] <=  8'h00;      memory[41863] <=  8'h00;      memory[41864] <=  8'h00;      memory[41865] <=  8'h00;      memory[41866] <=  8'h00;      memory[41867] <=  8'h00;      memory[41868] <=  8'h00;      memory[41869] <=  8'h00;      memory[41870] <=  8'h00;      memory[41871] <=  8'h00;      memory[41872] <=  8'h00;      memory[41873] <=  8'h00;      memory[41874] <=  8'h00;      memory[41875] <=  8'h00;      memory[41876] <=  8'h00;      memory[41877] <=  8'h00;      memory[41878] <=  8'h00;      memory[41879] <=  8'h00;      memory[41880] <=  8'h00;      memory[41881] <=  8'h00;      memory[41882] <=  8'h00;      memory[41883] <=  8'h00;      memory[41884] <=  8'h00;      memory[41885] <=  8'h00;      memory[41886] <=  8'h00;      memory[41887] <=  8'h00;      memory[41888] <=  8'h00;      memory[41889] <=  8'h00;      memory[41890] <=  8'h00;      memory[41891] <=  8'h00;      memory[41892] <=  8'h00;      memory[41893] <=  8'h00;      memory[41894] <=  8'h00;      memory[41895] <=  8'h00;      memory[41896] <=  8'h00;      memory[41897] <=  8'h00;      memory[41898] <=  8'h00;      memory[41899] <=  8'h00;      memory[41900] <=  8'h00;      memory[41901] <=  8'h00;      memory[41902] <=  8'h00;      memory[41903] <=  8'h00;      memory[41904] <=  8'h00;      memory[41905] <=  8'h00;      memory[41906] <=  8'h00;      memory[41907] <=  8'h00;      memory[41908] <=  8'h00;      memory[41909] <=  8'h00;      memory[41910] <=  8'h00;      memory[41911] <=  8'h00;      memory[41912] <=  8'h00;      memory[41913] <=  8'h00;      memory[41914] <=  8'h00;      memory[41915] <=  8'h00;      memory[41916] <=  8'h00;      memory[41917] <=  8'h00;      memory[41918] <=  8'h00;      memory[41919] <=  8'h00;      memory[41920] <=  8'h00;      memory[41921] <=  8'h00;      memory[41922] <=  8'h00;      memory[41923] <=  8'h00;      memory[41924] <=  8'h00;      memory[41925] <=  8'h00;      memory[41926] <=  8'h00;      memory[41927] <=  8'h00;      memory[41928] <=  8'h00;      memory[41929] <=  8'h00;      memory[41930] <=  8'h00;      memory[41931] <=  8'h00;      memory[41932] <=  8'h00;      memory[41933] <=  8'h00;      memory[41934] <=  8'h00;      memory[41935] <=  8'h00;      memory[41936] <=  8'h00;      memory[41937] <=  8'h00;      memory[41938] <=  8'h00;      memory[41939] <=  8'h00;      memory[41940] <=  8'h00;      memory[41941] <=  8'h00;      memory[41942] <=  8'h00;      memory[41943] <=  8'h00;      memory[41944] <=  8'h00;      memory[41945] <=  8'h00;      memory[41946] <=  8'h00;      memory[41947] <=  8'h00;      memory[41948] <=  8'h00;      memory[41949] <=  8'h00;      memory[41950] <=  8'h00;      memory[41951] <=  8'h00;      memory[41952] <=  8'h00;      memory[41953] <=  8'h00;      memory[41954] <=  8'h00;      memory[41955] <=  8'h00;      memory[41956] <=  8'h00;      memory[41957] <=  8'h00;      memory[41958] <=  8'h00;      memory[41959] <=  8'h00;      memory[41960] <=  8'h00;      memory[41961] <=  8'h00;      memory[41962] <=  8'h00;      memory[41963] <=  8'h00;      memory[41964] <=  8'h00;      memory[41965] <=  8'h00;      memory[41966] <=  8'h00;      memory[41967] <=  8'h00;      memory[41968] <=  8'h00;      memory[41969] <=  8'h00;      memory[41970] <=  8'h00;      memory[41971] <=  8'h00;      memory[41972] <=  8'h00;      memory[41973] <=  8'h00;      memory[41974] <=  8'h00;      memory[41975] <=  8'h00;      memory[41976] <=  8'h00;      memory[41977] <=  8'h00;      memory[41978] <=  8'h00;      memory[41979] <=  8'h00;      memory[41980] <=  8'h00;      memory[41981] <=  8'h00;      memory[41982] <=  8'h00;      memory[41983] <=  8'h00;      memory[41984] <=  8'h00;      memory[41985] <=  8'h00;      memory[41986] <=  8'h00;      memory[41987] <=  8'h00;      memory[41988] <=  8'h00;      memory[41989] <=  8'h00;      memory[41990] <=  8'h00;      memory[41991] <=  8'h00;      memory[41992] <=  8'h00;      memory[41993] <=  8'h00;      memory[41994] <=  8'h00;      memory[41995] <=  8'h00;      memory[41996] <=  8'h00;      memory[41997] <=  8'h00;      memory[41998] <=  8'h00;      memory[41999] <=  8'h00;      memory[42000] <=  8'h00;      memory[42001] <=  8'h00;      memory[42002] <=  8'h00;      memory[42003] <=  8'h00;      memory[42004] <=  8'h00;      memory[42005] <=  8'h00;      memory[42006] <=  8'h00;      memory[42007] <=  8'h00;      memory[42008] <=  8'h00;      memory[42009] <=  8'h00;      memory[42010] <=  8'h00;      memory[42011] <=  8'h00;      memory[42012] <=  8'h00;      memory[42013] <=  8'h00;      memory[42014] <=  8'h00;      memory[42015] <=  8'h00;      memory[42016] <=  8'h00;      memory[42017] <=  8'h00;      memory[42018] <=  8'h00;      memory[42019] <=  8'h00;      memory[42020] <=  8'h00;      memory[42021] <=  8'h00;      memory[42022] <=  8'h00;      memory[42023] <=  8'h00;      memory[42024] <=  8'h00;      memory[42025] <=  8'h00;      memory[42026] <=  8'h00;      memory[42027] <=  8'h00;      memory[42028] <=  8'h00;      memory[42029] <=  8'h00;      memory[42030] <=  8'h00;      memory[42031] <=  8'h00;      memory[42032] <=  8'h00;      memory[42033] <=  8'h00;      memory[42034] <=  8'h00;      memory[42035] <=  8'h00;      memory[42036] <=  8'h00;      memory[42037] <=  8'h00;      memory[42038] <=  8'h00;      memory[42039] <=  8'h00;      memory[42040] <=  8'h00;      memory[42041] <=  8'h00;      memory[42042] <=  8'h00;      memory[42043] <=  8'h00;      memory[42044] <=  8'h00;      memory[42045] <=  8'h00;      memory[42046] <=  8'h00;      memory[42047] <=  8'h00;      memory[42048] <=  8'h00;      memory[42049] <=  8'h00;      memory[42050] <=  8'h00;      memory[42051] <=  8'h00;      memory[42052] <=  8'h00;      memory[42053] <=  8'h00;      memory[42054] <=  8'h00;      memory[42055] <=  8'h00;      memory[42056] <=  8'h00;      memory[42057] <=  8'h00;      memory[42058] <=  8'h00;      memory[42059] <=  8'h00;      memory[42060] <=  8'h00;      memory[42061] <=  8'h00;      memory[42062] <=  8'h00;      memory[42063] <=  8'h00;      memory[42064] <=  8'h00;      memory[42065] <=  8'h00;      memory[42066] <=  8'h00;      memory[42067] <=  8'h00;      memory[42068] <=  8'h00;      memory[42069] <=  8'h00;      memory[42070] <=  8'h00;      memory[42071] <=  8'h00;      memory[42072] <=  8'h00;      memory[42073] <=  8'h00;      memory[42074] <=  8'h00;      memory[42075] <=  8'h00;      memory[42076] <=  8'h00;      memory[42077] <=  8'h00;      memory[42078] <=  8'h00;      memory[42079] <=  8'h00;      memory[42080] <=  8'h00;      memory[42081] <=  8'h00;      memory[42082] <=  8'h00;      memory[42083] <=  8'h00;      memory[42084] <=  8'h00;      memory[42085] <=  8'h00;      memory[42086] <=  8'h00;      memory[42087] <=  8'h00;      memory[42088] <=  8'h00;      memory[42089] <=  8'h00;      memory[42090] <=  8'h00;      memory[42091] <=  8'h00;      memory[42092] <=  8'h00;      memory[42093] <=  8'h00;      memory[42094] <=  8'h00;      memory[42095] <=  8'h00;      memory[42096] <=  8'h00;      memory[42097] <=  8'h00;      memory[42098] <=  8'h00;      memory[42099] <=  8'h00;      memory[42100] <=  8'h00;      memory[42101] <=  8'h00;      memory[42102] <=  8'h00;      memory[42103] <=  8'h00;      memory[42104] <=  8'h00;      memory[42105] <=  8'h00;      memory[42106] <=  8'h00;      memory[42107] <=  8'h00;      memory[42108] <=  8'h00;      memory[42109] <=  8'h00;      memory[42110] <=  8'h00;      memory[42111] <=  8'h00;      memory[42112] <=  8'h00;      memory[42113] <=  8'h00;      memory[42114] <=  8'h00;      memory[42115] <=  8'h00;      memory[42116] <=  8'h00;      memory[42117] <=  8'h00;      memory[42118] <=  8'h00;      memory[42119] <=  8'h00;      memory[42120] <=  8'h00;      memory[42121] <=  8'h00;      memory[42122] <=  8'h00;      memory[42123] <=  8'h00;      memory[42124] <=  8'h00;      memory[42125] <=  8'h00;      memory[42126] <=  8'h00;      memory[42127] <=  8'h00;      memory[42128] <=  8'h00;      memory[42129] <=  8'h00;      memory[42130] <=  8'h00;      memory[42131] <=  8'h00;      memory[42132] <=  8'h00;      memory[42133] <=  8'h00;      memory[42134] <=  8'h00;      memory[42135] <=  8'h00;      memory[42136] <=  8'h00;      memory[42137] <=  8'h00;      memory[42138] <=  8'h00;      memory[42139] <=  8'h00;      memory[42140] <=  8'h00;      memory[42141] <=  8'h00;      memory[42142] <=  8'h00;      memory[42143] <=  8'h00;      memory[42144] <=  8'h00;      memory[42145] <=  8'h00;      memory[42146] <=  8'h00;      memory[42147] <=  8'h00;      memory[42148] <=  8'h00;      memory[42149] <=  8'h00;      memory[42150] <=  8'h00;      memory[42151] <=  8'h00;      memory[42152] <=  8'h00;      memory[42153] <=  8'h00;      memory[42154] <=  8'h00;      memory[42155] <=  8'h00;      memory[42156] <=  8'h00;      memory[42157] <=  8'h00;      memory[42158] <=  8'h00;      memory[42159] <=  8'h00;      memory[42160] <=  8'h00;      memory[42161] <=  8'h00;      memory[42162] <=  8'h00;      memory[42163] <=  8'h00;      memory[42164] <=  8'h00;      memory[42165] <=  8'h00;      memory[42166] <=  8'h00;      memory[42167] <=  8'h00;      memory[42168] <=  8'h00;      memory[42169] <=  8'h00;      memory[42170] <=  8'h00;      memory[42171] <=  8'h00;      memory[42172] <=  8'h00;      memory[42173] <=  8'h00;      memory[42174] <=  8'h00;      memory[42175] <=  8'h00;      memory[42176] <=  8'h00;      memory[42177] <=  8'h00;      memory[42178] <=  8'h00;      memory[42179] <=  8'h00;      memory[42180] <=  8'h00;      memory[42181] <=  8'h00;      memory[42182] <=  8'h00;      memory[42183] <=  8'h00;      memory[42184] <=  8'h00;      memory[42185] <=  8'h00;      memory[42186] <=  8'h00;      memory[42187] <=  8'h00;      memory[42188] <=  8'h00;      memory[42189] <=  8'h00;      memory[42190] <=  8'h00;      memory[42191] <=  8'h00;      memory[42192] <=  8'h00;      memory[42193] <=  8'h00;      memory[42194] <=  8'h00;      memory[42195] <=  8'h00;      memory[42196] <=  8'h00;      memory[42197] <=  8'h00;      memory[42198] <=  8'h00;      memory[42199] <=  8'h00;      memory[42200] <=  8'h00;      memory[42201] <=  8'h00;      memory[42202] <=  8'h00;      memory[42203] <=  8'h00;      memory[42204] <=  8'h00;      memory[42205] <=  8'h00;      memory[42206] <=  8'h00;      memory[42207] <=  8'h00;      memory[42208] <=  8'h00;      memory[42209] <=  8'h00;      memory[42210] <=  8'h00;      memory[42211] <=  8'h00;      memory[42212] <=  8'h00;      memory[42213] <=  8'h00;      memory[42214] <=  8'h00;      memory[42215] <=  8'h00;      memory[42216] <=  8'h00;      memory[42217] <=  8'h00;      memory[42218] <=  8'h00;      memory[42219] <=  8'h00;      memory[42220] <=  8'h00;      memory[42221] <=  8'h00;      memory[42222] <=  8'h00;      memory[42223] <=  8'h00;      memory[42224] <=  8'h00;      memory[42225] <=  8'h00;      memory[42226] <=  8'h00;      memory[42227] <=  8'h00;      memory[42228] <=  8'h00;      memory[42229] <=  8'h00;      memory[42230] <=  8'h00;      memory[42231] <=  8'h00;      memory[42232] <=  8'h00;      memory[42233] <=  8'h00;      memory[42234] <=  8'h00;      memory[42235] <=  8'h00;      memory[42236] <=  8'h00;      memory[42237] <=  8'h00;      memory[42238] <=  8'h00;      memory[42239] <=  8'h00;      memory[42240] <=  8'h00;      memory[42241] <=  8'h00;      memory[42242] <=  8'h00;      memory[42243] <=  8'h00;      memory[42244] <=  8'h00;      memory[42245] <=  8'h00;      memory[42246] <=  8'h00;      memory[42247] <=  8'h00;      memory[42248] <=  8'h00;      memory[42249] <=  8'h00;      memory[42250] <=  8'h00;      memory[42251] <=  8'h00;      memory[42252] <=  8'h00;      memory[42253] <=  8'h00;      memory[42254] <=  8'h00;      memory[42255] <=  8'h00;      memory[42256] <=  8'h00;      memory[42257] <=  8'h00;      memory[42258] <=  8'h00;      memory[42259] <=  8'h00;      memory[42260] <=  8'h00;      memory[42261] <=  8'h00;      memory[42262] <=  8'h00;      memory[42263] <=  8'h00;      memory[42264] <=  8'h00;      memory[42265] <=  8'h00;      memory[42266] <=  8'h00;      memory[42267] <=  8'h00;      memory[42268] <=  8'h00;      memory[42269] <=  8'h00;      memory[42270] <=  8'h00;      memory[42271] <=  8'h00;      memory[42272] <=  8'h00;      memory[42273] <=  8'h00;      memory[42274] <=  8'h00;      memory[42275] <=  8'h00;      memory[42276] <=  8'h00;      memory[42277] <=  8'h00;      memory[42278] <=  8'h00;      memory[42279] <=  8'h00;      memory[42280] <=  8'h00;      memory[42281] <=  8'h00;      memory[42282] <=  8'h00;      memory[42283] <=  8'h00;      memory[42284] <=  8'h00;      memory[42285] <=  8'h00;      memory[42286] <=  8'h00;      memory[42287] <=  8'h00;      memory[42288] <=  8'h00;      memory[42289] <=  8'h00;      memory[42290] <=  8'h00;      memory[42291] <=  8'h00;      memory[42292] <=  8'h00;      memory[42293] <=  8'h00;      memory[42294] <=  8'h00;      memory[42295] <=  8'h00;      memory[42296] <=  8'h00;      memory[42297] <=  8'h00;      memory[42298] <=  8'h00;      memory[42299] <=  8'h00;      memory[42300] <=  8'h00;      memory[42301] <=  8'h00;      memory[42302] <=  8'h00;      memory[42303] <=  8'h00;      memory[42304] <=  8'h00;      memory[42305] <=  8'h00;      memory[42306] <=  8'h00;      memory[42307] <=  8'h00;      memory[42308] <=  8'h00;      memory[42309] <=  8'h00;      memory[42310] <=  8'h00;      memory[42311] <=  8'h00;      memory[42312] <=  8'h00;      memory[42313] <=  8'h00;      memory[42314] <=  8'h00;      memory[42315] <=  8'h00;      memory[42316] <=  8'h00;      memory[42317] <=  8'h00;      memory[42318] <=  8'h00;      memory[42319] <=  8'h00;      memory[42320] <=  8'h00;      memory[42321] <=  8'h00;      memory[42322] <=  8'h00;      memory[42323] <=  8'h00;      memory[42324] <=  8'h00;      memory[42325] <=  8'h00;      memory[42326] <=  8'h00;      memory[42327] <=  8'h00;      memory[42328] <=  8'h00;      memory[42329] <=  8'h00;      memory[42330] <=  8'h00;      memory[42331] <=  8'h00;      memory[42332] <=  8'h00;      memory[42333] <=  8'h00;      memory[42334] <=  8'h00;      memory[42335] <=  8'h00;      memory[42336] <=  8'h00;      memory[42337] <=  8'h00;      memory[42338] <=  8'h00;      memory[42339] <=  8'h00;      memory[42340] <=  8'h00;      memory[42341] <=  8'h00;      memory[42342] <=  8'h00;      memory[42343] <=  8'h00;      memory[42344] <=  8'h00;      memory[42345] <=  8'h00;      memory[42346] <=  8'h00;      memory[42347] <=  8'h00;      memory[42348] <=  8'h00;      memory[42349] <=  8'h00;      memory[42350] <=  8'h00;      memory[42351] <=  8'h00;      memory[42352] <=  8'h00;      memory[42353] <=  8'h00;      memory[42354] <=  8'h00;      memory[42355] <=  8'h00;      memory[42356] <=  8'h00;      memory[42357] <=  8'h00;      memory[42358] <=  8'h00;      memory[42359] <=  8'h00;      memory[42360] <=  8'h00;      memory[42361] <=  8'h00;      memory[42362] <=  8'h00;      memory[42363] <=  8'h00;      memory[42364] <=  8'h00;      memory[42365] <=  8'h00;      memory[42366] <=  8'h00;      memory[42367] <=  8'h00;      memory[42368] <=  8'h00;      memory[42369] <=  8'h00;      memory[42370] <=  8'h00;      memory[42371] <=  8'h00;      memory[42372] <=  8'h00;      memory[42373] <=  8'h00;      memory[42374] <=  8'h00;      memory[42375] <=  8'h00;      memory[42376] <=  8'h00;      memory[42377] <=  8'h00;      memory[42378] <=  8'h00;      memory[42379] <=  8'h00;      memory[42380] <=  8'h00;      memory[42381] <=  8'h00;      memory[42382] <=  8'h00;      memory[42383] <=  8'h00;      memory[42384] <=  8'h00;      memory[42385] <=  8'h00;      memory[42386] <=  8'h00;      memory[42387] <=  8'h00;      memory[42388] <=  8'h00;      memory[42389] <=  8'h00;      memory[42390] <=  8'h00;      memory[42391] <=  8'h00;      memory[42392] <=  8'h00;      memory[42393] <=  8'h00;      memory[42394] <=  8'h00;      memory[42395] <=  8'h00;      memory[42396] <=  8'h00;      memory[42397] <=  8'h00;      memory[42398] <=  8'h00;      memory[42399] <=  8'h00;      memory[42400] <=  8'h00;      memory[42401] <=  8'h00;      memory[42402] <=  8'h00;      memory[42403] <=  8'h00;      memory[42404] <=  8'h00;      memory[42405] <=  8'h00;      memory[42406] <=  8'h00;      memory[42407] <=  8'h00;      memory[42408] <=  8'h00;      memory[42409] <=  8'h00;      memory[42410] <=  8'h00;      memory[42411] <=  8'h00;      memory[42412] <=  8'h00;      memory[42413] <=  8'h00;      memory[42414] <=  8'h00;      memory[42415] <=  8'h00;      memory[42416] <=  8'h00;      memory[42417] <=  8'h00;      memory[42418] <=  8'h00;      memory[42419] <=  8'h00;      memory[42420] <=  8'h00;      memory[42421] <=  8'h00;      memory[42422] <=  8'h00;      memory[42423] <=  8'h00;      memory[42424] <=  8'h00;      memory[42425] <=  8'h00;      memory[42426] <=  8'h00;      memory[42427] <=  8'h00;      memory[42428] <=  8'h00;      memory[42429] <=  8'h00;      memory[42430] <=  8'h00;      memory[42431] <=  8'h00;      memory[42432] <=  8'h00;      memory[42433] <=  8'h00;      memory[42434] <=  8'h00;      memory[42435] <=  8'h00;      memory[42436] <=  8'h00;      memory[42437] <=  8'h00;      memory[42438] <=  8'h00;      memory[42439] <=  8'h00;      memory[42440] <=  8'h00;      memory[42441] <=  8'h00;      memory[42442] <=  8'h00;      memory[42443] <=  8'h00;      memory[42444] <=  8'h00;      memory[42445] <=  8'h00;      memory[42446] <=  8'h00;      memory[42447] <=  8'h00;      memory[42448] <=  8'h00;      memory[42449] <=  8'h00;      memory[42450] <=  8'h00;      memory[42451] <=  8'h00;      memory[42452] <=  8'h00;      memory[42453] <=  8'h00;      memory[42454] <=  8'h00;      memory[42455] <=  8'h00;      memory[42456] <=  8'h00;      memory[42457] <=  8'h00;      memory[42458] <=  8'h00;      memory[42459] <=  8'h00;      memory[42460] <=  8'h00;      memory[42461] <=  8'h00;      memory[42462] <=  8'h00;      memory[42463] <=  8'h00;      memory[42464] <=  8'h00;      memory[42465] <=  8'h00;      memory[42466] <=  8'h00;      memory[42467] <=  8'h00;      memory[42468] <=  8'h00;      memory[42469] <=  8'h00;      memory[42470] <=  8'h00;      memory[42471] <=  8'h00;      memory[42472] <=  8'h00;      memory[42473] <=  8'h00;      memory[42474] <=  8'h00;      memory[42475] <=  8'h00;      memory[42476] <=  8'h00;      memory[42477] <=  8'h00;      memory[42478] <=  8'h00;      memory[42479] <=  8'h00;      memory[42480] <=  8'h00;      memory[42481] <=  8'h00;      memory[42482] <=  8'h00;      memory[42483] <=  8'h00;      memory[42484] <=  8'h00;      memory[42485] <=  8'h00;      memory[42486] <=  8'h00;      memory[42487] <=  8'h00;      memory[42488] <=  8'h00;      memory[42489] <=  8'h00;      memory[42490] <=  8'h00;      memory[42491] <=  8'h00;      memory[42492] <=  8'h00;      memory[42493] <=  8'h00;      memory[42494] <=  8'h00;      memory[42495] <=  8'h00;      memory[42496] <=  8'h00;      memory[42497] <=  8'h00;      memory[42498] <=  8'h00;      memory[42499] <=  8'h00;      memory[42500] <=  8'h00;      memory[42501] <=  8'h00;      memory[42502] <=  8'h00;      memory[42503] <=  8'h00;      memory[42504] <=  8'h00;      memory[42505] <=  8'h00;      memory[42506] <=  8'h00;      memory[42507] <=  8'h00;      memory[42508] <=  8'h00;      memory[42509] <=  8'h00;      memory[42510] <=  8'h00;      memory[42511] <=  8'h00;      memory[42512] <=  8'h00;      memory[42513] <=  8'h00;      memory[42514] <=  8'h00;      memory[42515] <=  8'h00;      memory[42516] <=  8'h00;      memory[42517] <=  8'h00;      memory[42518] <=  8'h00;      memory[42519] <=  8'h00;      memory[42520] <=  8'h00;      memory[42521] <=  8'h00;      memory[42522] <=  8'h00;      memory[42523] <=  8'h00;      memory[42524] <=  8'h00;      memory[42525] <=  8'h00;      memory[42526] <=  8'h00;      memory[42527] <=  8'h00;      memory[42528] <=  8'h00;      memory[42529] <=  8'h00;      memory[42530] <=  8'h00;      memory[42531] <=  8'h00;      memory[42532] <=  8'h00;      memory[42533] <=  8'h00;      memory[42534] <=  8'h00;      memory[42535] <=  8'h00;      memory[42536] <=  8'h00;      memory[42537] <=  8'h00;      memory[42538] <=  8'h00;      memory[42539] <=  8'h00;      memory[42540] <=  8'h00;      memory[42541] <=  8'h00;      memory[42542] <=  8'h00;      memory[42543] <=  8'h00;      memory[42544] <=  8'h00;      memory[42545] <=  8'h00;      memory[42546] <=  8'h00;      memory[42547] <=  8'h00;      memory[42548] <=  8'h00;      memory[42549] <=  8'h00;      memory[42550] <=  8'h00;      memory[42551] <=  8'h00;      memory[42552] <=  8'h00;      memory[42553] <=  8'h00;      memory[42554] <=  8'h00;      memory[42555] <=  8'h00;      memory[42556] <=  8'h00;      memory[42557] <=  8'h00;      memory[42558] <=  8'h00;      memory[42559] <=  8'h00;      memory[42560] <=  8'h00;      memory[42561] <=  8'h00;      memory[42562] <=  8'h00;      memory[42563] <=  8'h00;      memory[42564] <=  8'h00;      memory[42565] <=  8'h00;      memory[42566] <=  8'h00;      memory[42567] <=  8'h00;      memory[42568] <=  8'h00;      memory[42569] <=  8'h00;      memory[42570] <=  8'h00;      memory[42571] <=  8'h00;      memory[42572] <=  8'h00;      memory[42573] <=  8'h00;      memory[42574] <=  8'h00;      memory[42575] <=  8'h00;      memory[42576] <=  8'h00;      memory[42577] <=  8'h00;      memory[42578] <=  8'h00;      memory[42579] <=  8'h00;      memory[42580] <=  8'h00;      memory[42581] <=  8'h00;      memory[42582] <=  8'h00;      memory[42583] <=  8'h00;      memory[42584] <=  8'h00;      memory[42585] <=  8'h00;      memory[42586] <=  8'h00;      memory[42587] <=  8'h00;      memory[42588] <=  8'h00;      memory[42589] <=  8'h00;      memory[42590] <=  8'h00;      memory[42591] <=  8'h00;      memory[42592] <=  8'h00;      memory[42593] <=  8'h00;      memory[42594] <=  8'h00;      memory[42595] <=  8'h00;      memory[42596] <=  8'h00;      memory[42597] <=  8'h00;      memory[42598] <=  8'h00;      memory[42599] <=  8'h00;      memory[42600] <=  8'h00;      memory[42601] <=  8'h00;      memory[42602] <=  8'h00;      memory[42603] <=  8'h00;      memory[42604] <=  8'h00;      memory[42605] <=  8'h00;      memory[42606] <=  8'h00;      memory[42607] <=  8'h00;      memory[42608] <=  8'h00;      memory[42609] <=  8'h00;      memory[42610] <=  8'h00;      memory[42611] <=  8'h00;      memory[42612] <=  8'h00;      memory[42613] <=  8'h00;      memory[42614] <=  8'h00;      memory[42615] <=  8'h00;      memory[42616] <=  8'h00;      memory[42617] <=  8'h00;      memory[42618] <=  8'h00;      memory[42619] <=  8'h00;      memory[42620] <=  8'h00;      memory[42621] <=  8'h00;      memory[42622] <=  8'h00;      memory[42623] <=  8'h00;      memory[42624] <=  8'h00;      memory[42625] <=  8'h00;      memory[42626] <=  8'h00;      memory[42627] <=  8'h00;      memory[42628] <=  8'h00;      memory[42629] <=  8'h00;      memory[42630] <=  8'h00;      memory[42631] <=  8'h00;      memory[42632] <=  8'h00;      memory[42633] <=  8'h00;      memory[42634] <=  8'h00;      memory[42635] <=  8'h00;      memory[42636] <=  8'h00;      memory[42637] <=  8'h00;      memory[42638] <=  8'h00;      memory[42639] <=  8'h00;      memory[42640] <=  8'h00;      memory[42641] <=  8'h00;      memory[42642] <=  8'h00;      memory[42643] <=  8'h00;      memory[42644] <=  8'h00;      memory[42645] <=  8'h00;      memory[42646] <=  8'h00;      memory[42647] <=  8'h00;      memory[42648] <=  8'h00;      memory[42649] <=  8'h00;      memory[42650] <=  8'h00;      memory[42651] <=  8'h00;      memory[42652] <=  8'h00;      memory[42653] <=  8'h00;      memory[42654] <=  8'h00;      memory[42655] <=  8'h00;      memory[42656] <=  8'h00;      memory[42657] <=  8'h00;      memory[42658] <=  8'h00;      memory[42659] <=  8'h00;      memory[42660] <=  8'h00;      memory[42661] <=  8'h00;      memory[42662] <=  8'h00;      memory[42663] <=  8'h00;      memory[42664] <=  8'h00;      memory[42665] <=  8'h00;      memory[42666] <=  8'h00;      memory[42667] <=  8'h00;      memory[42668] <=  8'h00;      memory[42669] <=  8'h00;      memory[42670] <=  8'h00;      memory[42671] <=  8'h00;      memory[42672] <=  8'h00;      memory[42673] <=  8'h00;      memory[42674] <=  8'h00;      memory[42675] <=  8'h00;      memory[42676] <=  8'h00;      memory[42677] <=  8'h00;      memory[42678] <=  8'h00;      memory[42679] <=  8'h00;      memory[42680] <=  8'h00;      memory[42681] <=  8'h00;      memory[42682] <=  8'h00;      memory[42683] <=  8'h00;      memory[42684] <=  8'h00;      memory[42685] <=  8'h00;      memory[42686] <=  8'h00;      memory[42687] <=  8'h00;      memory[42688] <=  8'h00;      memory[42689] <=  8'h00;      memory[42690] <=  8'h00;      memory[42691] <=  8'h00;      memory[42692] <=  8'h00;      memory[42693] <=  8'h00;      memory[42694] <=  8'h00;      memory[42695] <=  8'h00;      memory[42696] <=  8'h00;      memory[42697] <=  8'h00;      memory[42698] <=  8'h00;      memory[42699] <=  8'h00;      memory[42700] <=  8'h00;      memory[42701] <=  8'h00;      memory[42702] <=  8'h00;      memory[42703] <=  8'h00;      memory[42704] <=  8'h00;      memory[42705] <=  8'h00;      memory[42706] <=  8'h00;      memory[42707] <=  8'h00;      memory[42708] <=  8'h00;      memory[42709] <=  8'h00;      memory[42710] <=  8'h00;      memory[42711] <=  8'h00;      memory[42712] <=  8'h00;      memory[42713] <=  8'h00;      memory[42714] <=  8'h00;      memory[42715] <=  8'h00;      memory[42716] <=  8'h00;      memory[42717] <=  8'h00;      memory[42718] <=  8'h00;      memory[42719] <=  8'h00;      memory[42720] <=  8'h00;      memory[42721] <=  8'h00;      memory[42722] <=  8'h00;      memory[42723] <=  8'h00;      memory[42724] <=  8'h00;      memory[42725] <=  8'h00;      memory[42726] <=  8'h00;      memory[42727] <=  8'h00;      memory[42728] <=  8'h00;      memory[42729] <=  8'h00;      memory[42730] <=  8'h00;      memory[42731] <=  8'h00;      memory[42732] <=  8'h00;      memory[42733] <=  8'h00;      memory[42734] <=  8'h00;      memory[42735] <=  8'h00;      memory[42736] <=  8'h00;      memory[42737] <=  8'h00;      memory[42738] <=  8'h00;      memory[42739] <=  8'h00;      memory[42740] <=  8'h00;      memory[42741] <=  8'h00;      memory[42742] <=  8'h00;      memory[42743] <=  8'h00;      memory[42744] <=  8'h00;      memory[42745] <=  8'h00;      memory[42746] <=  8'h00;      memory[42747] <=  8'h00;      memory[42748] <=  8'h00;      memory[42749] <=  8'h00;      memory[42750] <=  8'h00;      memory[42751] <=  8'h00;      memory[42752] <=  8'h00;      memory[42753] <=  8'h00;      memory[42754] <=  8'h00;      memory[42755] <=  8'h00;      memory[42756] <=  8'h00;      memory[42757] <=  8'h00;      memory[42758] <=  8'h00;      memory[42759] <=  8'h00;      memory[42760] <=  8'h00;      memory[42761] <=  8'h00;      memory[42762] <=  8'h00;      memory[42763] <=  8'h00;      memory[42764] <=  8'h00;      memory[42765] <=  8'h00;      memory[42766] <=  8'h00;      memory[42767] <=  8'h00;      memory[42768] <=  8'h00;      memory[42769] <=  8'h00;      memory[42770] <=  8'h00;      memory[42771] <=  8'h00;      memory[42772] <=  8'h00;      memory[42773] <=  8'h00;      memory[42774] <=  8'h00;      memory[42775] <=  8'h00;      memory[42776] <=  8'h00;      memory[42777] <=  8'h00;      memory[42778] <=  8'h00;      memory[42779] <=  8'h00;      memory[42780] <=  8'h00;      memory[42781] <=  8'h00;      memory[42782] <=  8'h00;      memory[42783] <=  8'h00;      memory[42784] <=  8'h00;      memory[42785] <=  8'h00;      memory[42786] <=  8'h00;      memory[42787] <=  8'h00;      memory[42788] <=  8'h00;      memory[42789] <=  8'h00;      memory[42790] <=  8'h00;      memory[42791] <=  8'h00;      memory[42792] <=  8'h00;      memory[42793] <=  8'h00;      memory[42794] <=  8'h00;      memory[42795] <=  8'h00;      memory[42796] <=  8'h00;      memory[42797] <=  8'h00;      memory[42798] <=  8'h00;      memory[42799] <=  8'h00;      memory[42800] <=  8'h00;      memory[42801] <=  8'h00;      memory[42802] <=  8'h00;      memory[42803] <=  8'h00;      memory[42804] <=  8'h00;      memory[42805] <=  8'h00;      memory[42806] <=  8'h00;      memory[42807] <=  8'h00;      memory[42808] <=  8'h00;      memory[42809] <=  8'h00;      memory[42810] <=  8'h00;      memory[42811] <=  8'h00;      memory[42812] <=  8'h00;      memory[42813] <=  8'h00;      memory[42814] <=  8'h00;      memory[42815] <=  8'h00;      memory[42816] <=  8'h00;      memory[42817] <=  8'h00;      memory[42818] <=  8'h00;      memory[42819] <=  8'h00;      memory[42820] <=  8'h00;      memory[42821] <=  8'h00;      memory[42822] <=  8'h00;      memory[42823] <=  8'h00;      memory[42824] <=  8'h00;      memory[42825] <=  8'h00;      memory[42826] <=  8'h00;      memory[42827] <=  8'h00;      memory[42828] <=  8'h00;      memory[42829] <=  8'h00;      memory[42830] <=  8'h00;      memory[42831] <=  8'h00;      memory[42832] <=  8'h00;      memory[42833] <=  8'h00;      memory[42834] <=  8'h00;      memory[42835] <=  8'h00;      memory[42836] <=  8'h00;      memory[42837] <=  8'h00;      memory[42838] <=  8'h00;      memory[42839] <=  8'h00;      memory[42840] <=  8'h00;      memory[42841] <=  8'h00;      memory[42842] <=  8'h00;      memory[42843] <=  8'h00;      memory[42844] <=  8'h00;      memory[42845] <=  8'h00;      memory[42846] <=  8'h00;      memory[42847] <=  8'h00;      memory[42848] <=  8'h00;      memory[42849] <=  8'h00;      memory[42850] <=  8'h00;      memory[42851] <=  8'h00;      memory[42852] <=  8'h00;      memory[42853] <=  8'h00;      memory[42854] <=  8'h00;      memory[42855] <=  8'h00;      memory[42856] <=  8'h00;      memory[42857] <=  8'h00;      memory[42858] <=  8'h00;      memory[42859] <=  8'h00;      memory[42860] <=  8'h00;      memory[42861] <=  8'h00;      memory[42862] <=  8'h00;      memory[42863] <=  8'h00;      memory[42864] <=  8'h00;      memory[42865] <=  8'h00;      memory[42866] <=  8'h00;      memory[42867] <=  8'h00;      memory[42868] <=  8'h00;      memory[42869] <=  8'h00;      memory[42870] <=  8'h00;      memory[42871] <=  8'h00;      memory[42872] <=  8'h00;      memory[42873] <=  8'h00;      memory[42874] <=  8'h00;      memory[42875] <=  8'h00;      memory[42876] <=  8'h00;      memory[42877] <=  8'h00;      memory[42878] <=  8'h00;      memory[42879] <=  8'h00;      memory[42880] <=  8'h00;      memory[42881] <=  8'h00;      memory[42882] <=  8'h00;      memory[42883] <=  8'h00;      memory[42884] <=  8'h00;      memory[42885] <=  8'h00;      memory[42886] <=  8'h00;      memory[42887] <=  8'h00;      memory[42888] <=  8'h00;      memory[42889] <=  8'h00;      memory[42890] <=  8'h00;      memory[42891] <=  8'h00;      memory[42892] <=  8'h00;      memory[42893] <=  8'h00;      memory[42894] <=  8'h00;      memory[42895] <=  8'h00;      memory[42896] <=  8'h00;      memory[42897] <=  8'h00;      memory[42898] <=  8'h00;      memory[42899] <=  8'h00;      memory[42900] <=  8'h00;      memory[42901] <=  8'h00;      memory[42902] <=  8'h00;      memory[42903] <=  8'h00;      memory[42904] <=  8'h00;      memory[42905] <=  8'h00;      memory[42906] <=  8'h00;      memory[42907] <=  8'h00;      memory[42908] <=  8'h00;      memory[42909] <=  8'h00;      memory[42910] <=  8'h00;      memory[42911] <=  8'h00;      memory[42912] <=  8'h00;      memory[42913] <=  8'h00;      memory[42914] <=  8'h00;      memory[42915] <=  8'h00;      memory[42916] <=  8'h00;      memory[42917] <=  8'h00;      memory[42918] <=  8'h00;      memory[42919] <=  8'h00;      memory[42920] <=  8'h00;      memory[42921] <=  8'h00;      memory[42922] <=  8'h00;      memory[42923] <=  8'h00;      memory[42924] <=  8'h00;      memory[42925] <=  8'h00;      memory[42926] <=  8'h00;      memory[42927] <=  8'h00;      memory[42928] <=  8'h00;      memory[42929] <=  8'h00;      memory[42930] <=  8'h00;      memory[42931] <=  8'h00;      memory[42932] <=  8'h00;      memory[42933] <=  8'h00;      memory[42934] <=  8'h00;      memory[42935] <=  8'h00;      memory[42936] <=  8'h00;      memory[42937] <=  8'h00;      memory[42938] <=  8'h00;      memory[42939] <=  8'h00;      memory[42940] <=  8'h00;      memory[42941] <=  8'h00;      memory[42942] <=  8'h00;      memory[42943] <=  8'h00;      memory[42944] <=  8'h00;      memory[42945] <=  8'h00;      memory[42946] <=  8'h00;      memory[42947] <=  8'h00;      memory[42948] <=  8'h00;      memory[42949] <=  8'h00;      memory[42950] <=  8'h00;      memory[42951] <=  8'h00;      memory[42952] <=  8'h00;      memory[42953] <=  8'h00;      memory[42954] <=  8'h00;      memory[42955] <=  8'h00;      memory[42956] <=  8'h00;      memory[42957] <=  8'h00;      memory[42958] <=  8'h00;      memory[42959] <=  8'h00;      memory[42960] <=  8'h00;      memory[42961] <=  8'h00;      memory[42962] <=  8'h00;      memory[42963] <=  8'h00;      memory[42964] <=  8'h00;      memory[42965] <=  8'h00;      memory[42966] <=  8'h00;      memory[42967] <=  8'h00;      memory[42968] <=  8'h00;      memory[42969] <=  8'h00;      memory[42970] <=  8'h00;      memory[42971] <=  8'h00;      memory[42972] <=  8'h00;      memory[42973] <=  8'h00;      memory[42974] <=  8'h00;      memory[42975] <=  8'h00;      memory[42976] <=  8'h00;      memory[42977] <=  8'h00;      memory[42978] <=  8'h00;      memory[42979] <=  8'h00;      memory[42980] <=  8'h00;      memory[42981] <=  8'h00;      memory[42982] <=  8'h00;      memory[42983] <=  8'h00;      memory[42984] <=  8'h00;      memory[42985] <=  8'h00;      memory[42986] <=  8'h00;      memory[42987] <=  8'h00;      memory[42988] <=  8'h00;      memory[42989] <=  8'h00;      memory[42990] <=  8'h00;      memory[42991] <=  8'h00;      memory[42992] <=  8'h00;      memory[42993] <=  8'h00;      memory[42994] <=  8'h00;      memory[42995] <=  8'h00;      memory[42996] <=  8'h00;      memory[42997] <=  8'h00;      memory[42998] <=  8'h00;      memory[42999] <=  8'h00;      memory[43000] <=  8'h00;      memory[43001] <=  8'h00;      memory[43002] <=  8'h00;      memory[43003] <=  8'h00;      memory[43004] <=  8'h00;      memory[43005] <=  8'h00;      memory[43006] <=  8'h00;      memory[43007] <=  8'h00;      memory[43008] <=  8'h00;      memory[43009] <=  8'h00;      memory[43010] <=  8'h00;      memory[43011] <=  8'h00;      memory[43012] <=  8'h00;      memory[43013] <=  8'h00;      memory[43014] <=  8'h00;      memory[43015] <=  8'h00;      memory[43016] <=  8'h00;      memory[43017] <=  8'h00;      memory[43018] <=  8'h00;      memory[43019] <=  8'h00;      memory[43020] <=  8'h00;      memory[43021] <=  8'h00;      memory[43022] <=  8'h00;      memory[43023] <=  8'h00;      memory[43024] <=  8'h00;      memory[43025] <=  8'h00;      memory[43026] <=  8'h00;      memory[43027] <=  8'h00;      memory[43028] <=  8'h00;      memory[43029] <=  8'h00;      memory[43030] <=  8'h00;      memory[43031] <=  8'h00;      memory[43032] <=  8'h00;      memory[43033] <=  8'h00;      memory[43034] <=  8'h00;      memory[43035] <=  8'h00;      memory[43036] <=  8'h00;      memory[43037] <=  8'h00;      memory[43038] <=  8'h00;      memory[43039] <=  8'h00;      memory[43040] <=  8'h00;      memory[43041] <=  8'h00;      memory[43042] <=  8'h00;      memory[43043] <=  8'h00;      memory[43044] <=  8'h00;      memory[43045] <=  8'h00;      memory[43046] <=  8'h00;      memory[43047] <=  8'h00;      memory[43048] <=  8'h00;      memory[43049] <=  8'h00;      memory[43050] <=  8'h00;      memory[43051] <=  8'h00;      memory[43052] <=  8'h00;      memory[43053] <=  8'h00;      memory[43054] <=  8'h00;      memory[43055] <=  8'h00;      memory[43056] <=  8'h00;      memory[43057] <=  8'h00;      memory[43058] <=  8'h00;      memory[43059] <=  8'h00;      memory[43060] <=  8'h00;      memory[43061] <=  8'h00;      memory[43062] <=  8'h00;      memory[43063] <=  8'h00;      memory[43064] <=  8'h00;      memory[43065] <=  8'h00;      memory[43066] <=  8'h00;      memory[43067] <=  8'h00;      memory[43068] <=  8'h00;      memory[43069] <=  8'h00;      memory[43070] <=  8'h00;      memory[43071] <=  8'h00;      memory[43072] <=  8'h00;      memory[43073] <=  8'h00;      memory[43074] <=  8'h00;      memory[43075] <=  8'h00;      memory[43076] <=  8'h00;      memory[43077] <=  8'h00;      memory[43078] <=  8'h00;      memory[43079] <=  8'h00;      memory[43080] <=  8'h00;      memory[43081] <=  8'h00;      memory[43082] <=  8'h00;      memory[43083] <=  8'h00;      memory[43084] <=  8'h00;      memory[43085] <=  8'h00;      memory[43086] <=  8'h00;      memory[43087] <=  8'h00;      memory[43088] <=  8'h00;      memory[43089] <=  8'h00;      memory[43090] <=  8'h00;      memory[43091] <=  8'h00;      memory[43092] <=  8'h00;      memory[43093] <=  8'h00;      memory[43094] <=  8'h00;      memory[43095] <=  8'h00;      memory[43096] <=  8'h00;      memory[43097] <=  8'h00;      memory[43098] <=  8'h00;      memory[43099] <=  8'h00;      memory[43100] <=  8'h00;      memory[43101] <=  8'h00;      memory[43102] <=  8'h00;      memory[43103] <=  8'h00;      memory[43104] <=  8'h00;      memory[43105] <=  8'h00;      memory[43106] <=  8'h00;      memory[43107] <=  8'h00;      memory[43108] <=  8'h00;      memory[43109] <=  8'h00;      memory[43110] <=  8'h00;      memory[43111] <=  8'h00;      memory[43112] <=  8'h00;      memory[43113] <=  8'h00;      memory[43114] <=  8'h00;      memory[43115] <=  8'h00;      memory[43116] <=  8'h00;      memory[43117] <=  8'h00;      memory[43118] <=  8'h00;      memory[43119] <=  8'h00;      memory[43120] <=  8'h00;      memory[43121] <=  8'h00;      memory[43122] <=  8'h00;      memory[43123] <=  8'h00;      memory[43124] <=  8'h00;      memory[43125] <=  8'h00;      memory[43126] <=  8'h00;      memory[43127] <=  8'h00;      memory[43128] <=  8'h00;      memory[43129] <=  8'h00;      memory[43130] <=  8'h00;      memory[43131] <=  8'h00;      memory[43132] <=  8'h00;      memory[43133] <=  8'h00;      memory[43134] <=  8'h00;      memory[43135] <=  8'h00;      memory[43136] <=  8'h00;      memory[43137] <=  8'h00;      memory[43138] <=  8'h00;      memory[43139] <=  8'h00;      memory[43140] <=  8'h00;      memory[43141] <=  8'h00;      memory[43142] <=  8'h00;      memory[43143] <=  8'h00;      memory[43144] <=  8'h00;      memory[43145] <=  8'h00;      memory[43146] <=  8'h00;      memory[43147] <=  8'h00;      memory[43148] <=  8'h00;      memory[43149] <=  8'h00;      memory[43150] <=  8'h00;      memory[43151] <=  8'h00;      memory[43152] <=  8'h00;      memory[43153] <=  8'h00;      memory[43154] <=  8'h00;      memory[43155] <=  8'h00;      memory[43156] <=  8'h00;      memory[43157] <=  8'h00;      memory[43158] <=  8'h00;      memory[43159] <=  8'h00;      memory[43160] <=  8'h00;      memory[43161] <=  8'h00;      memory[43162] <=  8'h00;      memory[43163] <=  8'h00;      memory[43164] <=  8'h00;      memory[43165] <=  8'h00;      memory[43166] <=  8'h00;      memory[43167] <=  8'h00;      memory[43168] <=  8'h00;      memory[43169] <=  8'h00;      memory[43170] <=  8'h00;      memory[43171] <=  8'h00;      memory[43172] <=  8'h00;      memory[43173] <=  8'h00;      memory[43174] <=  8'h00;      memory[43175] <=  8'h00;      memory[43176] <=  8'h00;      memory[43177] <=  8'h00;      memory[43178] <=  8'h00;      memory[43179] <=  8'h00;      memory[43180] <=  8'h00;      memory[43181] <=  8'h00;      memory[43182] <=  8'h00;      memory[43183] <=  8'h00;      memory[43184] <=  8'h00;      memory[43185] <=  8'h00;      memory[43186] <=  8'h00;      memory[43187] <=  8'h00;      memory[43188] <=  8'h00;      memory[43189] <=  8'h00;      memory[43190] <=  8'h00;      memory[43191] <=  8'h00;      memory[43192] <=  8'h00;      memory[43193] <=  8'h00;      memory[43194] <=  8'h00;      memory[43195] <=  8'h00;      memory[43196] <=  8'h00;      memory[43197] <=  8'h00;      memory[43198] <=  8'h00;      memory[43199] <=  8'h00;      memory[43200] <=  8'h00;      memory[43201] <=  8'h00;      memory[43202] <=  8'h00;      memory[43203] <=  8'h00;      memory[43204] <=  8'h00;      memory[43205] <=  8'h00;      memory[43206] <=  8'h00;      memory[43207] <=  8'h00;      memory[43208] <=  8'h00;      memory[43209] <=  8'h00;      memory[43210] <=  8'h00;      memory[43211] <=  8'h00;      memory[43212] <=  8'h00;      memory[43213] <=  8'h00;      memory[43214] <=  8'h00;      memory[43215] <=  8'h00;      memory[43216] <=  8'h00;      memory[43217] <=  8'h00;      memory[43218] <=  8'h00;      memory[43219] <=  8'h00;      memory[43220] <=  8'h00;      memory[43221] <=  8'h00;      memory[43222] <=  8'h00;      memory[43223] <=  8'h00;      memory[43224] <=  8'h00;      memory[43225] <=  8'h00;      memory[43226] <=  8'h00;      memory[43227] <=  8'h00;      memory[43228] <=  8'h00;      memory[43229] <=  8'h00;      memory[43230] <=  8'h00;      memory[43231] <=  8'h00;      memory[43232] <=  8'h00;      memory[43233] <=  8'h00;      memory[43234] <=  8'h00;      memory[43235] <=  8'h00;      memory[43236] <=  8'h00;      memory[43237] <=  8'h00;      memory[43238] <=  8'h00;      memory[43239] <=  8'h00;      memory[43240] <=  8'h00;      memory[43241] <=  8'h00;      memory[43242] <=  8'h00;      memory[43243] <=  8'h00;      memory[43244] <=  8'h00;      memory[43245] <=  8'h00;      memory[43246] <=  8'h00;      memory[43247] <=  8'h00;      memory[43248] <=  8'h00;      memory[43249] <=  8'h00;      memory[43250] <=  8'h00;      memory[43251] <=  8'h00;      memory[43252] <=  8'h00;      memory[43253] <=  8'h00;      memory[43254] <=  8'h00;      memory[43255] <=  8'h00;      memory[43256] <=  8'h00;      memory[43257] <=  8'h00;      memory[43258] <=  8'h00;      memory[43259] <=  8'h00;      memory[43260] <=  8'h00;      memory[43261] <=  8'h00;      memory[43262] <=  8'h00;      memory[43263] <=  8'h00;      memory[43264] <=  8'h00;      memory[43265] <=  8'h00;      memory[43266] <=  8'h00;      memory[43267] <=  8'h00;      memory[43268] <=  8'h00;      memory[43269] <=  8'h00;      memory[43270] <=  8'h00;      memory[43271] <=  8'h00;      memory[43272] <=  8'h00;      memory[43273] <=  8'h00;      memory[43274] <=  8'h00;      memory[43275] <=  8'h00;      memory[43276] <=  8'h00;      memory[43277] <=  8'h00;      memory[43278] <=  8'h00;      memory[43279] <=  8'h00;      memory[43280] <=  8'h00;      memory[43281] <=  8'h00;      memory[43282] <=  8'h00;      memory[43283] <=  8'h00;      memory[43284] <=  8'h00;      memory[43285] <=  8'h00;      memory[43286] <=  8'h00;      memory[43287] <=  8'h00;      memory[43288] <=  8'h00;      memory[43289] <=  8'h00;      memory[43290] <=  8'h00;      memory[43291] <=  8'h00;      memory[43292] <=  8'h00;      memory[43293] <=  8'h00;      memory[43294] <=  8'h00;      memory[43295] <=  8'h00;      memory[43296] <=  8'h00;      memory[43297] <=  8'h00;      memory[43298] <=  8'h00;      memory[43299] <=  8'h00;      memory[43300] <=  8'h00;      memory[43301] <=  8'h00;      memory[43302] <=  8'h00;      memory[43303] <=  8'h00;      memory[43304] <=  8'h00;      memory[43305] <=  8'h00;      memory[43306] <=  8'h00;      memory[43307] <=  8'h00;      memory[43308] <=  8'h00;      memory[43309] <=  8'h00;      memory[43310] <=  8'h00;      memory[43311] <=  8'h00;      memory[43312] <=  8'h00;      memory[43313] <=  8'h00;      memory[43314] <=  8'h00;      memory[43315] <=  8'h00;      memory[43316] <=  8'h00;      memory[43317] <=  8'h00;      memory[43318] <=  8'h00;      memory[43319] <=  8'h00;      memory[43320] <=  8'h00;      memory[43321] <=  8'h00;      memory[43322] <=  8'h00;      memory[43323] <=  8'h00;      memory[43324] <=  8'h00;      memory[43325] <=  8'h00;      memory[43326] <=  8'h00;      memory[43327] <=  8'h00;      memory[43328] <=  8'h00;      memory[43329] <=  8'h00;      memory[43330] <=  8'h00;      memory[43331] <=  8'h00;      memory[43332] <=  8'h00;      memory[43333] <=  8'h00;      memory[43334] <=  8'h00;      memory[43335] <=  8'h00;      memory[43336] <=  8'h00;      memory[43337] <=  8'h00;      memory[43338] <=  8'h00;      memory[43339] <=  8'h00;      memory[43340] <=  8'h00;      memory[43341] <=  8'h00;      memory[43342] <=  8'h00;      memory[43343] <=  8'h00;      memory[43344] <=  8'h00;      memory[43345] <=  8'h00;      memory[43346] <=  8'h00;      memory[43347] <=  8'h00;      memory[43348] <=  8'h00;      memory[43349] <=  8'h00;      memory[43350] <=  8'h00;      memory[43351] <=  8'h00;      memory[43352] <=  8'h00;      memory[43353] <=  8'h00;      memory[43354] <=  8'h00;      memory[43355] <=  8'h00;      memory[43356] <=  8'h00;      memory[43357] <=  8'h00;      memory[43358] <=  8'h00;      memory[43359] <=  8'h00;      memory[43360] <=  8'h00;      memory[43361] <=  8'h00;      memory[43362] <=  8'h00;      memory[43363] <=  8'h00;      memory[43364] <=  8'h00;      memory[43365] <=  8'h00;      memory[43366] <=  8'h00;      memory[43367] <=  8'h00;      memory[43368] <=  8'h00;      memory[43369] <=  8'h00;      memory[43370] <=  8'h00;      memory[43371] <=  8'h00;      memory[43372] <=  8'h00;      memory[43373] <=  8'h00;      memory[43374] <=  8'h00;      memory[43375] <=  8'h00;      memory[43376] <=  8'h00;      memory[43377] <=  8'h00;      memory[43378] <=  8'h00;      memory[43379] <=  8'h00;      memory[43380] <=  8'h00;      memory[43381] <=  8'h00;      memory[43382] <=  8'h00;      memory[43383] <=  8'h00;      memory[43384] <=  8'h00;      memory[43385] <=  8'h00;      memory[43386] <=  8'h00;      memory[43387] <=  8'h00;      memory[43388] <=  8'h00;      memory[43389] <=  8'h00;      memory[43390] <=  8'h00;      memory[43391] <=  8'h00;      memory[43392] <=  8'h00;      memory[43393] <=  8'h00;      memory[43394] <=  8'h00;      memory[43395] <=  8'h00;      memory[43396] <=  8'h00;      memory[43397] <=  8'h00;      memory[43398] <=  8'h00;      memory[43399] <=  8'h00;      memory[43400] <=  8'h00;      memory[43401] <=  8'h00;      memory[43402] <=  8'h00;      memory[43403] <=  8'h00;      memory[43404] <=  8'h00;      memory[43405] <=  8'h00;      memory[43406] <=  8'h00;      memory[43407] <=  8'h00;      memory[43408] <=  8'h00;      memory[43409] <=  8'h00;      memory[43410] <=  8'h00;      memory[43411] <=  8'h00;      memory[43412] <=  8'h00;      memory[43413] <=  8'h00;      memory[43414] <=  8'h00;      memory[43415] <=  8'h00;      memory[43416] <=  8'h00;      memory[43417] <=  8'h00;      memory[43418] <=  8'h00;      memory[43419] <=  8'h00;      memory[43420] <=  8'h00;      memory[43421] <=  8'h00;      memory[43422] <=  8'h00;      memory[43423] <=  8'h00;      memory[43424] <=  8'h00;      memory[43425] <=  8'h00;      memory[43426] <=  8'h00;      memory[43427] <=  8'h00;      memory[43428] <=  8'h00;      memory[43429] <=  8'h00;      memory[43430] <=  8'h00;      memory[43431] <=  8'h00;      memory[43432] <=  8'h00;      memory[43433] <=  8'h00;      memory[43434] <=  8'h00;      memory[43435] <=  8'h00;      memory[43436] <=  8'h00;      memory[43437] <=  8'h00;      memory[43438] <=  8'h00;      memory[43439] <=  8'h00;      memory[43440] <=  8'h00;      memory[43441] <=  8'h00;      memory[43442] <=  8'h00;      memory[43443] <=  8'h00;      memory[43444] <=  8'h00;      memory[43445] <=  8'h00;      memory[43446] <=  8'h00;      memory[43447] <=  8'h00;      memory[43448] <=  8'h00;      memory[43449] <=  8'h00;      memory[43450] <=  8'h00;      memory[43451] <=  8'h00;      memory[43452] <=  8'h00;      memory[43453] <=  8'h00;      memory[43454] <=  8'h00;      memory[43455] <=  8'h00;      memory[43456] <=  8'h00;      memory[43457] <=  8'h00;      memory[43458] <=  8'h00;      memory[43459] <=  8'h00;      memory[43460] <=  8'h00;      memory[43461] <=  8'h00;      memory[43462] <=  8'h00;      memory[43463] <=  8'h00;      memory[43464] <=  8'h00;      memory[43465] <=  8'h00;      memory[43466] <=  8'h00;      memory[43467] <=  8'h00;      memory[43468] <=  8'h00;      memory[43469] <=  8'h00;      memory[43470] <=  8'h00;      memory[43471] <=  8'h00;      memory[43472] <=  8'h00;      memory[43473] <=  8'h00;      memory[43474] <=  8'h00;      memory[43475] <=  8'h00;      memory[43476] <=  8'h00;      memory[43477] <=  8'h00;      memory[43478] <=  8'h00;      memory[43479] <=  8'h00;      memory[43480] <=  8'h00;      memory[43481] <=  8'h00;      memory[43482] <=  8'h00;      memory[43483] <=  8'h00;      memory[43484] <=  8'h00;      memory[43485] <=  8'h00;      memory[43486] <=  8'h00;      memory[43487] <=  8'h00;      memory[43488] <=  8'h00;      memory[43489] <=  8'h00;      memory[43490] <=  8'h00;      memory[43491] <=  8'h00;      memory[43492] <=  8'h00;      memory[43493] <=  8'h00;      memory[43494] <=  8'h00;      memory[43495] <=  8'h00;      memory[43496] <=  8'h00;      memory[43497] <=  8'h00;      memory[43498] <=  8'h00;      memory[43499] <=  8'h00;      memory[43500] <=  8'h00;      memory[43501] <=  8'h00;      memory[43502] <=  8'h00;      memory[43503] <=  8'h00;      memory[43504] <=  8'h00;      memory[43505] <=  8'h00;      memory[43506] <=  8'h00;      memory[43507] <=  8'h00;      memory[43508] <=  8'h00;      memory[43509] <=  8'h00;      memory[43510] <=  8'h00;      memory[43511] <=  8'h00;      memory[43512] <=  8'h00;      memory[43513] <=  8'h00;      memory[43514] <=  8'h00;      memory[43515] <=  8'h00;      memory[43516] <=  8'h00;      memory[43517] <=  8'h00;      memory[43518] <=  8'h00;      memory[43519] <=  8'h00;      memory[43520] <=  8'h00;      memory[43521] <=  8'h00;      memory[43522] <=  8'h00;      memory[43523] <=  8'h00;      memory[43524] <=  8'h00;      memory[43525] <=  8'h00;      memory[43526] <=  8'h00;      memory[43527] <=  8'h00;      memory[43528] <=  8'h00;      memory[43529] <=  8'h00;      memory[43530] <=  8'h00;      memory[43531] <=  8'h00;      memory[43532] <=  8'h00;      memory[43533] <=  8'h00;      memory[43534] <=  8'h00;      memory[43535] <=  8'h00;      memory[43536] <=  8'h00;      memory[43537] <=  8'h00;      memory[43538] <=  8'h00;      memory[43539] <=  8'h00;      memory[43540] <=  8'h00;      memory[43541] <=  8'h00;      memory[43542] <=  8'h00;      memory[43543] <=  8'h00;      memory[43544] <=  8'h00;      memory[43545] <=  8'h00;      memory[43546] <=  8'h00;      memory[43547] <=  8'h00;      memory[43548] <=  8'h00;      memory[43549] <=  8'h00;      memory[43550] <=  8'h00;      memory[43551] <=  8'h00;      memory[43552] <=  8'h00;      memory[43553] <=  8'h00;      memory[43554] <=  8'h00;      memory[43555] <=  8'h00;      memory[43556] <=  8'h00;      memory[43557] <=  8'h00;      memory[43558] <=  8'h00;      memory[43559] <=  8'h00;      memory[43560] <=  8'h00;      memory[43561] <=  8'h00;      memory[43562] <=  8'h00;      memory[43563] <=  8'h00;      memory[43564] <=  8'h00;      memory[43565] <=  8'h00;      memory[43566] <=  8'h00;      memory[43567] <=  8'h00;      memory[43568] <=  8'h00;      memory[43569] <=  8'h00;      memory[43570] <=  8'h00;      memory[43571] <=  8'h00;      memory[43572] <=  8'h00;      memory[43573] <=  8'h00;      memory[43574] <=  8'h00;      memory[43575] <=  8'h00;      memory[43576] <=  8'h00;      memory[43577] <=  8'h00;      memory[43578] <=  8'h00;      memory[43579] <=  8'h00;      memory[43580] <=  8'h00;      memory[43581] <=  8'h00;      memory[43582] <=  8'h00;      memory[43583] <=  8'h00;      memory[43584] <=  8'h00;      memory[43585] <=  8'h00;      memory[43586] <=  8'h00;      memory[43587] <=  8'h00;      memory[43588] <=  8'h00;      memory[43589] <=  8'h00;      memory[43590] <=  8'h00;      memory[43591] <=  8'h00;      memory[43592] <=  8'h00;      memory[43593] <=  8'h00;      memory[43594] <=  8'h00;      memory[43595] <=  8'h00;      memory[43596] <=  8'h00;      memory[43597] <=  8'h00;      memory[43598] <=  8'h00;      memory[43599] <=  8'h00;      memory[43600] <=  8'h00;      memory[43601] <=  8'h00;      memory[43602] <=  8'h00;      memory[43603] <=  8'h00;      memory[43604] <=  8'h00;      memory[43605] <=  8'h00;      memory[43606] <=  8'h00;      memory[43607] <=  8'h00;      memory[43608] <=  8'h00;      memory[43609] <=  8'h00;      memory[43610] <=  8'h00;      memory[43611] <=  8'h00;      memory[43612] <=  8'h00;      memory[43613] <=  8'h00;      memory[43614] <=  8'h00;      memory[43615] <=  8'h00;      memory[43616] <=  8'h00;      memory[43617] <=  8'h00;      memory[43618] <=  8'h00;      memory[43619] <=  8'h00;      memory[43620] <=  8'h00;      memory[43621] <=  8'h00;      memory[43622] <=  8'h00;      memory[43623] <=  8'h00;      memory[43624] <=  8'h00;      memory[43625] <=  8'h00;      memory[43626] <=  8'h00;      memory[43627] <=  8'h00;      memory[43628] <=  8'h00;      memory[43629] <=  8'h00;      memory[43630] <=  8'h00;      memory[43631] <=  8'h00;      memory[43632] <=  8'h00;      memory[43633] <=  8'h00;      memory[43634] <=  8'h00;      memory[43635] <=  8'h00;      memory[43636] <=  8'h00;      memory[43637] <=  8'h00;      memory[43638] <=  8'h00;      memory[43639] <=  8'h00;      memory[43640] <=  8'h00;      memory[43641] <=  8'h00;      memory[43642] <=  8'h00;      memory[43643] <=  8'h00;      memory[43644] <=  8'h00;      memory[43645] <=  8'h00;      memory[43646] <=  8'h00;      memory[43647] <=  8'h00;      memory[43648] <=  8'h00;      memory[43649] <=  8'h00;      memory[43650] <=  8'h00;      memory[43651] <=  8'h00;      memory[43652] <=  8'h00;      memory[43653] <=  8'h00;      memory[43654] <=  8'h00;      memory[43655] <=  8'h00;      memory[43656] <=  8'h00;      memory[43657] <=  8'h00;      memory[43658] <=  8'h00;      memory[43659] <=  8'h00;      memory[43660] <=  8'h00;      memory[43661] <=  8'h00;      memory[43662] <=  8'h00;      memory[43663] <=  8'h00;      memory[43664] <=  8'h00;      memory[43665] <=  8'h00;      memory[43666] <=  8'h00;      memory[43667] <=  8'h00;      memory[43668] <=  8'h00;      memory[43669] <=  8'h00;      memory[43670] <=  8'h00;      memory[43671] <=  8'h00;      memory[43672] <=  8'h00;      memory[43673] <=  8'h00;      memory[43674] <=  8'h00;      memory[43675] <=  8'h00;      memory[43676] <=  8'h00;      memory[43677] <=  8'h00;      memory[43678] <=  8'h00;      memory[43679] <=  8'h00;      memory[43680] <=  8'h00;      memory[43681] <=  8'h00;      memory[43682] <=  8'h00;      memory[43683] <=  8'h00;      memory[43684] <=  8'h00;      memory[43685] <=  8'h00;      memory[43686] <=  8'h00;      memory[43687] <=  8'h00;      memory[43688] <=  8'h00;      memory[43689] <=  8'h00;      memory[43690] <=  8'h00;      memory[43691] <=  8'h00;      memory[43692] <=  8'h00;      memory[43693] <=  8'h00;      memory[43694] <=  8'h00;      memory[43695] <=  8'h00;      memory[43696] <=  8'h00;      memory[43697] <=  8'h00;      memory[43698] <=  8'h00;      memory[43699] <=  8'h00;      memory[43700] <=  8'h00;      memory[43701] <=  8'h00;      memory[43702] <=  8'h00;      memory[43703] <=  8'h00;      memory[43704] <=  8'h00;      memory[43705] <=  8'h00;      memory[43706] <=  8'h00;      memory[43707] <=  8'h00;      memory[43708] <=  8'h00;      memory[43709] <=  8'h00;      memory[43710] <=  8'h00;      memory[43711] <=  8'h00;      memory[43712] <=  8'h00;      memory[43713] <=  8'h00;      memory[43714] <=  8'h00;      memory[43715] <=  8'h00;      memory[43716] <=  8'h00;      memory[43717] <=  8'h00;      memory[43718] <=  8'h00;      memory[43719] <=  8'h00;      memory[43720] <=  8'h00;      memory[43721] <=  8'h00;      memory[43722] <=  8'h00;      memory[43723] <=  8'h00;      memory[43724] <=  8'h00;      memory[43725] <=  8'h00;      memory[43726] <=  8'h00;      memory[43727] <=  8'h00;      memory[43728] <=  8'h00;      memory[43729] <=  8'h00;      memory[43730] <=  8'h00;      memory[43731] <=  8'h00;      memory[43732] <=  8'h00;      memory[43733] <=  8'h00;      memory[43734] <=  8'h00;      memory[43735] <=  8'h00;      memory[43736] <=  8'h00;      memory[43737] <=  8'h00;      memory[43738] <=  8'h00;      memory[43739] <=  8'h00;      memory[43740] <=  8'h00;      memory[43741] <=  8'h00;      memory[43742] <=  8'h00;      memory[43743] <=  8'h00;      memory[43744] <=  8'h00;      memory[43745] <=  8'h00;      memory[43746] <=  8'h00;      memory[43747] <=  8'h00;      memory[43748] <=  8'h00;      memory[43749] <=  8'h00;      memory[43750] <=  8'h00;      memory[43751] <=  8'h00;      memory[43752] <=  8'h00;      memory[43753] <=  8'h00;      memory[43754] <=  8'h00;      memory[43755] <=  8'h00;      memory[43756] <=  8'h00;      memory[43757] <=  8'h00;      memory[43758] <=  8'h00;      memory[43759] <=  8'h00;      memory[43760] <=  8'h00;      memory[43761] <=  8'h00;      memory[43762] <=  8'h00;      memory[43763] <=  8'h00;      memory[43764] <=  8'h00;      memory[43765] <=  8'h00;      memory[43766] <=  8'h00;      memory[43767] <=  8'h00;      memory[43768] <=  8'h00;      memory[43769] <=  8'h00;      memory[43770] <=  8'h00;      memory[43771] <=  8'h00;      memory[43772] <=  8'h00;      memory[43773] <=  8'h00;      memory[43774] <=  8'h00;      memory[43775] <=  8'h00;      memory[43776] <=  8'h00;      memory[43777] <=  8'h00;      memory[43778] <=  8'h00;      memory[43779] <=  8'h00;      memory[43780] <=  8'h00;      memory[43781] <=  8'h00;      memory[43782] <=  8'h00;      memory[43783] <=  8'h00;      memory[43784] <=  8'h00;      memory[43785] <=  8'h00;      memory[43786] <=  8'h00;      memory[43787] <=  8'h00;      memory[43788] <=  8'h00;      memory[43789] <=  8'h00;      memory[43790] <=  8'h00;      memory[43791] <=  8'h00;      memory[43792] <=  8'h00;      memory[43793] <=  8'h00;      memory[43794] <=  8'h00;      memory[43795] <=  8'h00;      memory[43796] <=  8'h00;      memory[43797] <=  8'h00;      memory[43798] <=  8'h00;      memory[43799] <=  8'h00;      memory[43800] <=  8'h00;      memory[43801] <=  8'h00;      memory[43802] <=  8'h00;      memory[43803] <=  8'h00;      memory[43804] <=  8'h00;      memory[43805] <=  8'h00;      memory[43806] <=  8'h00;      memory[43807] <=  8'h00;      memory[43808] <=  8'h00;      memory[43809] <=  8'h00;      memory[43810] <=  8'h00;      memory[43811] <=  8'h00;      memory[43812] <=  8'h00;      memory[43813] <=  8'h00;      memory[43814] <=  8'h00;      memory[43815] <=  8'h00;      memory[43816] <=  8'h00;      memory[43817] <=  8'h00;      memory[43818] <=  8'h00;      memory[43819] <=  8'h00;      memory[43820] <=  8'h00;      memory[43821] <=  8'h00;      memory[43822] <=  8'h00;      memory[43823] <=  8'h00;      memory[43824] <=  8'h00;      memory[43825] <=  8'h00;      memory[43826] <=  8'h00;      memory[43827] <=  8'h00;      memory[43828] <=  8'h00;      memory[43829] <=  8'h00;      memory[43830] <=  8'h00;      memory[43831] <=  8'h00;      memory[43832] <=  8'h00;      memory[43833] <=  8'h00;      memory[43834] <=  8'h00;      memory[43835] <=  8'h00;      memory[43836] <=  8'h00;      memory[43837] <=  8'h00;      memory[43838] <=  8'h00;      memory[43839] <=  8'h00;      memory[43840] <=  8'h00;      memory[43841] <=  8'h00;      memory[43842] <=  8'h00;      memory[43843] <=  8'h00;      memory[43844] <=  8'h00;      memory[43845] <=  8'h00;      memory[43846] <=  8'h00;      memory[43847] <=  8'h00;      memory[43848] <=  8'h00;      memory[43849] <=  8'h00;      memory[43850] <=  8'h00;      memory[43851] <=  8'h00;      memory[43852] <=  8'h00;      memory[43853] <=  8'h00;      memory[43854] <=  8'h00;      memory[43855] <=  8'h00;      memory[43856] <=  8'h00;      memory[43857] <=  8'h00;      memory[43858] <=  8'h00;      memory[43859] <=  8'h00;      memory[43860] <=  8'h00;      memory[43861] <=  8'h00;      memory[43862] <=  8'h00;      memory[43863] <=  8'h00;      memory[43864] <=  8'h00;      memory[43865] <=  8'h00;      memory[43866] <=  8'h00;      memory[43867] <=  8'h00;      memory[43868] <=  8'h00;      memory[43869] <=  8'h00;      memory[43870] <=  8'h00;      memory[43871] <=  8'h00;      memory[43872] <=  8'h00;      memory[43873] <=  8'h00;      memory[43874] <=  8'h00;      memory[43875] <=  8'h00;      memory[43876] <=  8'h00;      memory[43877] <=  8'h00;      memory[43878] <=  8'h00;      memory[43879] <=  8'h00;      memory[43880] <=  8'h00;      memory[43881] <=  8'h00;      memory[43882] <=  8'h00;      memory[43883] <=  8'h00;      memory[43884] <=  8'h00;      memory[43885] <=  8'h00;      memory[43886] <=  8'h00;      memory[43887] <=  8'h00;      memory[43888] <=  8'h00;      memory[43889] <=  8'h00;      memory[43890] <=  8'h00;      memory[43891] <=  8'h00;      memory[43892] <=  8'h00;      memory[43893] <=  8'h00;      memory[43894] <=  8'h00;      memory[43895] <=  8'h00;      memory[43896] <=  8'h00;      memory[43897] <=  8'h00;      memory[43898] <=  8'h00;      memory[43899] <=  8'h00;      memory[43900] <=  8'h00;      memory[43901] <=  8'h00;      memory[43902] <=  8'h00;      memory[43903] <=  8'h00;      memory[43904] <=  8'h00;      memory[43905] <=  8'h00;      memory[43906] <=  8'h00;      memory[43907] <=  8'h00;      memory[43908] <=  8'h00;      memory[43909] <=  8'h00;      memory[43910] <=  8'h00;      memory[43911] <=  8'h00;      memory[43912] <=  8'h00;      memory[43913] <=  8'h00;      memory[43914] <=  8'h00;      memory[43915] <=  8'h00;      memory[43916] <=  8'h00;      memory[43917] <=  8'h00;      memory[43918] <=  8'h00;      memory[43919] <=  8'h00;      memory[43920] <=  8'h00;      memory[43921] <=  8'h00;      memory[43922] <=  8'h00;      memory[43923] <=  8'h00;      memory[43924] <=  8'h00;      memory[43925] <=  8'h00;      memory[43926] <=  8'h00;      memory[43927] <=  8'h00;      memory[43928] <=  8'h00;      memory[43929] <=  8'h00;      memory[43930] <=  8'h00;      memory[43931] <=  8'h00;      memory[43932] <=  8'h00;      memory[43933] <=  8'h00;      memory[43934] <=  8'h00;      memory[43935] <=  8'h00;      memory[43936] <=  8'h00;      memory[43937] <=  8'h00;      memory[43938] <=  8'h00;      memory[43939] <=  8'h00;      memory[43940] <=  8'h00;      memory[43941] <=  8'h00;      memory[43942] <=  8'h00;      memory[43943] <=  8'h00;      memory[43944] <=  8'h00;      memory[43945] <=  8'h00;      memory[43946] <=  8'h00;      memory[43947] <=  8'h00;      memory[43948] <=  8'h00;      memory[43949] <=  8'h00;      memory[43950] <=  8'h00;      memory[43951] <=  8'h00;      memory[43952] <=  8'h00;      memory[43953] <=  8'h00;      memory[43954] <=  8'h00;      memory[43955] <=  8'h00;      memory[43956] <=  8'h00;      memory[43957] <=  8'h00;      memory[43958] <=  8'h00;      memory[43959] <=  8'h00;      memory[43960] <=  8'h00;      memory[43961] <=  8'h00;      memory[43962] <=  8'h00;      memory[43963] <=  8'h00;      memory[43964] <=  8'h00;      memory[43965] <=  8'h00;      memory[43966] <=  8'h00;      memory[43967] <=  8'h00;      memory[43968] <=  8'h00;      memory[43969] <=  8'h00;      memory[43970] <=  8'h00;      memory[43971] <=  8'h00;      memory[43972] <=  8'h00;      memory[43973] <=  8'h00;      memory[43974] <=  8'h00;      memory[43975] <=  8'h00;      memory[43976] <=  8'h00;      memory[43977] <=  8'h00;      memory[43978] <=  8'h00;      memory[43979] <=  8'h00;      memory[43980] <=  8'h00;      memory[43981] <=  8'h00;      memory[43982] <=  8'h00;      memory[43983] <=  8'h00;      memory[43984] <=  8'h00;      memory[43985] <=  8'h00;      memory[43986] <=  8'h00;      memory[43987] <=  8'h00;      memory[43988] <=  8'h00;      memory[43989] <=  8'h00;      memory[43990] <=  8'h00;      memory[43991] <=  8'h00;      memory[43992] <=  8'h00;      memory[43993] <=  8'h00;      memory[43994] <=  8'h00;      memory[43995] <=  8'h00;      memory[43996] <=  8'h00;      memory[43997] <=  8'h00;      memory[43998] <=  8'h00;      memory[43999] <=  8'h00;      memory[44000] <=  8'h00;      memory[44001] <=  8'h00;      memory[44002] <=  8'h00;      memory[44003] <=  8'h00;      memory[44004] <=  8'h00;      memory[44005] <=  8'h00;      memory[44006] <=  8'h00;      memory[44007] <=  8'h00;      memory[44008] <=  8'h00;      memory[44009] <=  8'h00;      memory[44010] <=  8'h00;      memory[44011] <=  8'h00;      memory[44012] <=  8'h00;      memory[44013] <=  8'h00;      memory[44014] <=  8'h00;      memory[44015] <=  8'h00;      memory[44016] <=  8'h00;      memory[44017] <=  8'h00;      memory[44018] <=  8'h00;      memory[44019] <=  8'h00;      memory[44020] <=  8'h00;      memory[44021] <=  8'h00;      memory[44022] <=  8'h00;      memory[44023] <=  8'h00;      memory[44024] <=  8'h00;      memory[44025] <=  8'h00;      memory[44026] <=  8'h00;      memory[44027] <=  8'h00;      memory[44028] <=  8'h00;      memory[44029] <=  8'h00;      memory[44030] <=  8'h00;      memory[44031] <=  8'h00;      memory[44032] <=  8'h00;      memory[44033] <=  8'h00;      memory[44034] <=  8'h00;      memory[44035] <=  8'h00;      memory[44036] <=  8'h00;      memory[44037] <=  8'h00;      memory[44038] <=  8'h00;      memory[44039] <=  8'h00;      memory[44040] <=  8'h00;      memory[44041] <=  8'h00;      memory[44042] <=  8'h00;      memory[44043] <=  8'h00;      memory[44044] <=  8'h00;      memory[44045] <=  8'h00;      memory[44046] <=  8'h00;      memory[44047] <=  8'h00;      memory[44048] <=  8'h00;      memory[44049] <=  8'h00;      memory[44050] <=  8'h00;      memory[44051] <=  8'h00;      memory[44052] <=  8'h00;      memory[44053] <=  8'h00;      memory[44054] <=  8'h00;      memory[44055] <=  8'h00;      memory[44056] <=  8'h00;      memory[44057] <=  8'h00;      memory[44058] <=  8'h00;      memory[44059] <=  8'h00;      memory[44060] <=  8'h00;      memory[44061] <=  8'h00;      memory[44062] <=  8'h00;      memory[44063] <=  8'h00;      memory[44064] <=  8'h00;      memory[44065] <=  8'h00;      memory[44066] <=  8'h00;      memory[44067] <=  8'h00;      memory[44068] <=  8'h00;      memory[44069] <=  8'h00;      memory[44070] <=  8'h00;      memory[44071] <=  8'h00;      memory[44072] <=  8'h00;      memory[44073] <=  8'h00;      memory[44074] <=  8'h00;      memory[44075] <=  8'h00;      memory[44076] <=  8'h00;      memory[44077] <=  8'h00;      memory[44078] <=  8'h00;      memory[44079] <=  8'h00;      memory[44080] <=  8'h00;      memory[44081] <=  8'h00;      memory[44082] <=  8'h00;      memory[44083] <=  8'h00;      memory[44084] <=  8'h00;      memory[44085] <=  8'h00;      memory[44086] <=  8'h00;      memory[44087] <=  8'h00;      memory[44088] <=  8'h00;      memory[44089] <=  8'h00;      memory[44090] <=  8'h00;      memory[44091] <=  8'h00;      memory[44092] <=  8'h00;      memory[44093] <=  8'h00;      memory[44094] <=  8'h00;      memory[44095] <=  8'h00;      memory[44096] <=  8'h00;      memory[44097] <=  8'h00;      memory[44098] <=  8'h00;      memory[44099] <=  8'h00;      memory[44100] <=  8'h00;      memory[44101] <=  8'h00;      memory[44102] <=  8'h00;      memory[44103] <=  8'h00;      memory[44104] <=  8'h00;      memory[44105] <=  8'h00;      memory[44106] <=  8'h00;      memory[44107] <=  8'h00;      memory[44108] <=  8'h00;      memory[44109] <=  8'h00;      memory[44110] <=  8'h00;      memory[44111] <=  8'h00;      memory[44112] <=  8'h00;      memory[44113] <=  8'h00;      memory[44114] <=  8'h00;      memory[44115] <=  8'h00;      memory[44116] <=  8'h00;      memory[44117] <=  8'h00;      memory[44118] <=  8'h00;      memory[44119] <=  8'h00;      memory[44120] <=  8'h00;      memory[44121] <=  8'h00;      memory[44122] <=  8'h00;      memory[44123] <=  8'h00;      memory[44124] <=  8'h00;      memory[44125] <=  8'h00;      memory[44126] <=  8'h00;      memory[44127] <=  8'h00;      memory[44128] <=  8'h00;      memory[44129] <=  8'h00;      memory[44130] <=  8'h00;      memory[44131] <=  8'h00;      memory[44132] <=  8'h00;      memory[44133] <=  8'h00;      memory[44134] <=  8'h00;      memory[44135] <=  8'h00;      memory[44136] <=  8'h00;      memory[44137] <=  8'h00;      memory[44138] <=  8'h00;      memory[44139] <=  8'h00;      memory[44140] <=  8'h00;      memory[44141] <=  8'h00;      memory[44142] <=  8'h00;      memory[44143] <=  8'h00;      memory[44144] <=  8'h00;      memory[44145] <=  8'h00;      memory[44146] <=  8'h00;      memory[44147] <=  8'h00;      memory[44148] <=  8'h00;      memory[44149] <=  8'h00;      memory[44150] <=  8'h00;      memory[44151] <=  8'h00;      memory[44152] <=  8'h00;      memory[44153] <=  8'h00;      memory[44154] <=  8'h00;      memory[44155] <=  8'h00;      memory[44156] <=  8'h00;      memory[44157] <=  8'h00;      memory[44158] <=  8'h00;      memory[44159] <=  8'h00;      memory[44160] <=  8'h00;      memory[44161] <=  8'h00;      memory[44162] <=  8'h00;      memory[44163] <=  8'h00;      memory[44164] <=  8'h00;      memory[44165] <=  8'h00;      memory[44166] <=  8'h00;      memory[44167] <=  8'h00;      memory[44168] <=  8'h00;      memory[44169] <=  8'h00;      memory[44170] <=  8'h00;      memory[44171] <=  8'h00;      memory[44172] <=  8'h00;      memory[44173] <=  8'h00;      memory[44174] <=  8'h00;      memory[44175] <=  8'h00;      memory[44176] <=  8'h00;      memory[44177] <=  8'h00;      memory[44178] <=  8'h00;      memory[44179] <=  8'h00;      memory[44180] <=  8'h00;      memory[44181] <=  8'h00;      memory[44182] <=  8'h00;      memory[44183] <=  8'h00;      memory[44184] <=  8'h00;      memory[44185] <=  8'h00;      memory[44186] <=  8'h00;      memory[44187] <=  8'h00;      memory[44188] <=  8'h00;      memory[44189] <=  8'h00;      memory[44190] <=  8'h00;      memory[44191] <=  8'h00;      memory[44192] <=  8'h00;      memory[44193] <=  8'h00;      memory[44194] <=  8'h00;      memory[44195] <=  8'h00;      memory[44196] <=  8'h00;      memory[44197] <=  8'h00;      memory[44198] <=  8'h00;      memory[44199] <=  8'h00;      memory[44200] <=  8'h00;      memory[44201] <=  8'h00;      memory[44202] <=  8'h00;      memory[44203] <=  8'h00;      memory[44204] <=  8'h00;      memory[44205] <=  8'h00;      memory[44206] <=  8'h00;      memory[44207] <=  8'h00;      memory[44208] <=  8'h00;      memory[44209] <=  8'h00;      memory[44210] <=  8'h00;      memory[44211] <=  8'h00;      memory[44212] <=  8'h00;      memory[44213] <=  8'h00;      memory[44214] <=  8'h00;      memory[44215] <=  8'h00;      memory[44216] <=  8'h00;      memory[44217] <=  8'h00;      memory[44218] <=  8'h00;      memory[44219] <=  8'h00;      memory[44220] <=  8'h00;      memory[44221] <=  8'h00;      memory[44222] <=  8'h00;      memory[44223] <=  8'h00;      memory[44224] <=  8'h00;      memory[44225] <=  8'h00;      memory[44226] <=  8'h00;      memory[44227] <=  8'h00;      memory[44228] <=  8'h00;      memory[44229] <=  8'h00;      memory[44230] <=  8'h00;      memory[44231] <=  8'h00;      memory[44232] <=  8'h00;      memory[44233] <=  8'h00;      memory[44234] <=  8'h00;      memory[44235] <=  8'h00;      memory[44236] <=  8'h00;      memory[44237] <=  8'h00;      memory[44238] <=  8'h00;      memory[44239] <=  8'h00;      memory[44240] <=  8'h00;      memory[44241] <=  8'h00;      memory[44242] <=  8'h00;      memory[44243] <=  8'h00;      memory[44244] <=  8'h00;      memory[44245] <=  8'h00;      memory[44246] <=  8'h00;      memory[44247] <=  8'h00;      memory[44248] <=  8'h00;      memory[44249] <=  8'h00;      memory[44250] <=  8'h00;      memory[44251] <=  8'h00;      memory[44252] <=  8'h00;      memory[44253] <=  8'h00;      memory[44254] <=  8'h00;      memory[44255] <=  8'h00;      memory[44256] <=  8'h00;      memory[44257] <=  8'h00;      memory[44258] <=  8'h00;      memory[44259] <=  8'h00;      memory[44260] <=  8'h00;      memory[44261] <=  8'h00;      memory[44262] <=  8'h00;      memory[44263] <=  8'h00;      memory[44264] <=  8'h00;      memory[44265] <=  8'h00;      memory[44266] <=  8'h00;      memory[44267] <=  8'h00;      memory[44268] <=  8'h00;      memory[44269] <=  8'h00;      memory[44270] <=  8'h00;      memory[44271] <=  8'h00;      memory[44272] <=  8'h00;      memory[44273] <=  8'h00;      memory[44274] <=  8'h00;      memory[44275] <=  8'h00;      memory[44276] <=  8'h00;      memory[44277] <=  8'h00;      memory[44278] <=  8'h00;      memory[44279] <=  8'h00;      memory[44280] <=  8'h00;      memory[44281] <=  8'h00;      memory[44282] <=  8'h00;      memory[44283] <=  8'h00;      memory[44284] <=  8'h00;      memory[44285] <=  8'h00;      memory[44286] <=  8'h00;      memory[44287] <=  8'h00;      memory[44288] <=  8'h00;      memory[44289] <=  8'h00;      memory[44290] <=  8'h00;      memory[44291] <=  8'h00;      memory[44292] <=  8'h00;      memory[44293] <=  8'h00;      memory[44294] <=  8'h00;      memory[44295] <=  8'h00;      memory[44296] <=  8'h00;      memory[44297] <=  8'h00;      memory[44298] <=  8'h00;      memory[44299] <=  8'h00;      memory[44300] <=  8'h00;      memory[44301] <=  8'h00;      memory[44302] <=  8'h00;      memory[44303] <=  8'h00;      memory[44304] <=  8'h00;      memory[44305] <=  8'h00;      memory[44306] <=  8'h00;      memory[44307] <=  8'h00;      memory[44308] <=  8'h00;      memory[44309] <=  8'h00;      memory[44310] <=  8'h00;      memory[44311] <=  8'h00;      memory[44312] <=  8'h00;      memory[44313] <=  8'h00;      memory[44314] <=  8'h00;      memory[44315] <=  8'h00;      memory[44316] <=  8'h00;      memory[44317] <=  8'h00;      memory[44318] <=  8'h00;      memory[44319] <=  8'h00;      memory[44320] <=  8'h00;      memory[44321] <=  8'h00;      memory[44322] <=  8'h00;      memory[44323] <=  8'h00;      memory[44324] <=  8'h00;      memory[44325] <=  8'h00;      memory[44326] <=  8'h00;      memory[44327] <=  8'h00;      memory[44328] <=  8'h00;      memory[44329] <=  8'h00;      memory[44330] <=  8'h00;      memory[44331] <=  8'h00;      memory[44332] <=  8'h00;      memory[44333] <=  8'h00;      memory[44334] <=  8'h00;      memory[44335] <=  8'h00;      memory[44336] <=  8'h00;      memory[44337] <=  8'h00;      memory[44338] <=  8'h00;      memory[44339] <=  8'h00;      memory[44340] <=  8'h00;      memory[44341] <=  8'h00;      memory[44342] <=  8'h00;      memory[44343] <=  8'h00;      memory[44344] <=  8'h00;      memory[44345] <=  8'h00;      memory[44346] <=  8'h00;      memory[44347] <=  8'h00;      memory[44348] <=  8'h00;      memory[44349] <=  8'h00;      memory[44350] <=  8'h00;      memory[44351] <=  8'h00;      memory[44352] <=  8'h00;      memory[44353] <=  8'h00;      memory[44354] <=  8'h00;      memory[44355] <=  8'h00;      memory[44356] <=  8'h00;      memory[44357] <=  8'h00;      memory[44358] <=  8'h00;      memory[44359] <=  8'h00;      memory[44360] <=  8'h00;      memory[44361] <=  8'h00;      memory[44362] <=  8'h00;      memory[44363] <=  8'h00;      memory[44364] <=  8'h00;      memory[44365] <=  8'h00;      memory[44366] <=  8'h00;      memory[44367] <=  8'h00;      memory[44368] <=  8'h00;      memory[44369] <=  8'h00;      memory[44370] <=  8'h00;      memory[44371] <=  8'h00;      memory[44372] <=  8'h00;      memory[44373] <=  8'h00;      memory[44374] <=  8'h00;      memory[44375] <=  8'h00;      memory[44376] <=  8'h00;      memory[44377] <=  8'h00;      memory[44378] <=  8'h00;      memory[44379] <=  8'h00;      memory[44380] <=  8'h00;      memory[44381] <=  8'h00;      memory[44382] <=  8'h00;      memory[44383] <=  8'h00;      memory[44384] <=  8'h00;      memory[44385] <=  8'h00;      memory[44386] <=  8'h00;      memory[44387] <=  8'h00;      memory[44388] <=  8'h00;      memory[44389] <=  8'h00;      memory[44390] <=  8'h00;      memory[44391] <=  8'h00;      memory[44392] <=  8'h00;      memory[44393] <=  8'h00;      memory[44394] <=  8'h00;      memory[44395] <=  8'h00;      memory[44396] <=  8'h00;      memory[44397] <=  8'h00;      memory[44398] <=  8'h00;      memory[44399] <=  8'h00;      memory[44400] <=  8'h00;      memory[44401] <=  8'h00;      memory[44402] <=  8'h00;      memory[44403] <=  8'h00;      memory[44404] <=  8'h00;      memory[44405] <=  8'h00;      memory[44406] <=  8'h00;      memory[44407] <=  8'h00;      memory[44408] <=  8'h00;      memory[44409] <=  8'h00;      memory[44410] <=  8'h00;      memory[44411] <=  8'h00;      memory[44412] <=  8'h00;      memory[44413] <=  8'h00;      memory[44414] <=  8'h00;      memory[44415] <=  8'h00;      memory[44416] <=  8'h00;      memory[44417] <=  8'h00;      memory[44418] <=  8'h00;      memory[44419] <=  8'h00;      memory[44420] <=  8'h00;      memory[44421] <=  8'h00;      memory[44422] <=  8'h00;      memory[44423] <=  8'h00;      memory[44424] <=  8'h00;      memory[44425] <=  8'h00;      memory[44426] <=  8'h00;      memory[44427] <=  8'h00;      memory[44428] <=  8'h00;      memory[44429] <=  8'h00;      memory[44430] <=  8'h00;      memory[44431] <=  8'h00;      memory[44432] <=  8'h00;      memory[44433] <=  8'h00;      memory[44434] <=  8'h00;      memory[44435] <=  8'h00;      memory[44436] <=  8'h00;      memory[44437] <=  8'h00;      memory[44438] <=  8'h00;      memory[44439] <=  8'h00;      memory[44440] <=  8'h00;      memory[44441] <=  8'h00;      memory[44442] <=  8'h00;      memory[44443] <=  8'h00;      memory[44444] <=  8'h00;      memory[44445] <=  8'h00;      memory[44446] <=  8'h00;      memory[44447] <=  8'h00;      memory[44448] <=  8'h00;      memory[44449] <=  8'h00;      memory[44450] <=  8'h00;      memory[44451] <=  8'h00;      memory[44452] <=  8'h00;      memory[44453] <=  8'h00;      memory[44454] <=  8'h00;      memory[44455] <=  8'h00;      memory[44456] <=  8'h00;      memory[44457] <=  8'h00;      memory[44458] <=  8'h00;      memory[44459] <=  8'h00;      memory[44460] <=  8'h00;      memory[44461] <=  8'h00;      memory[44462] <=  8'h00;      memory[44463] <=  8'h00;      memory[44464] <=  8'h00;      memory[44465] <=  8'h00;      memory[44466] <=  8'h00;      memory[44467] <=  8'h00;      memory[44468] <=  8'h00;      memory[44469] <=  8'h00;      memory[44470] <=  8'h00;      memory[44471] <=  8'h00;      memory[44472] <=  8'h00;      memory[44473] <=  8'h00;      memory[44474] <=  8'h00;      memory[44475] <=  8'h00;      memory[44476] <=  8'h00;      memory[44477] <=  8'h00;      memory[44478] <=  8'h00;      memory[44479] <=  8'h00;      memory[44480] <=  8'h00;      memory[44481] <=  8'h00;      memory[44482] <=  8'h00;      memory[44483] <=  8'h00;      memory[44484] <=  8'h00;      memory[44485] <=  8'h00;      memory[44486] <=  8'h00;      memory[44487] <=  8'h00;      memory[44488] <=  8'h00;      memory[44489] <=  8'h00;      memory[44490] <=  8'h00;      memory[44491] <=  8'h00;      memory[44492] <=  8'h00;      memory[44493] <=  8'h00;      memory[44494] <=  8'h00;      memory[44495] <=  8'h00;      memory[44496] <=  8'h00;      memory[44497] <=  8'h00;      memory[44498] <=  8'h00;      memory[44499] <=  8'h00;      memory[44500] <=  8'h00;      memory[44501] <=  8'h00;      memory[44502] <=  8'h00;      memory[44503] <=  8'h00;      memory[44504] <=  8'h00;      memory[44505] <=  8'h00;      memory[44506] <=  8'h00;      memory[44507] <=  8'h00;      memory[44508] <=  8'h00;      memory[44509] <=  8'h00;      memory[44510] <=  8'h00;      memory[44511] <=  8'h00;      memory[44512] <=  8'h00;      memory[44513] <=  8'h00;      memory[44514] <=  8'h00;      memory[44515] <=  8'h00;      memory[44516] <=  8'h00;      memory[44517] <=  8'h00;      memory[44518] <=  8'h00;      memory[44519] <=  8'h00;      memory[44520] <=  8'h00;      memory[44521] <=  8'h00;      memory[44522] <=  8'h00;      memory[44523] <=  8'h00;      memory[44524] <=  8'h00;      memory[44525] <=  8'h00;      memory[44526] <=  8'h00;      memory[44527] <=  8'h00;      memory[44528] <=  8'h00;      memory[44529] <=  8'h00;      memory[44530] <=  8'h00;      memory[44531] <=  8'h00;      memory[44532] <=  8'h00;      memory[44533] <=  8'h00;      memory[44534] <=  8'h00;      memory[44535] <=  8'h00;      memory[44536] <=  8'h00;      memory[44537] <=  8'h00;      memory[44538] <=  8'h00;      memory[44539] <=  8'h00;      memory[44540] <=  8'h00;      memory[44541] <=  8'h00;      memory[44542] <=  8'h00;      memory[44543] <=  8'h00;      memory[44544] <=  8'h00;      memory[44545] <=  8'h00;      memory[44546] <=  8'h00;      memory[44547] <=  8'h00;      memory[44548] <=  8'h00;      memory[44549] <=  8'h00;      memory[44550] <=  8'h00;      memory[44551] <=  8'h00;      memory[44552] <=  8'h00;      memory[44553] <=  8'h00;      memory[44554] <=  8'h00;      memory[44555] <=  8'h00;      memory[44556] <=  8'h00;      memory[44557] <=  8'h00;      memory[44558] <=  8'h00;      memory[44559] <=  8'h00;      memory[44560] <=  8'h00;      memory[44561] <=  8'h00;      memory[44562] <=  8'h00;      memory[44563] <=  8'h00;      memory[44564] <=  8'h00;      memory[44565] <=  8'h00;      memory[44566] <=  8'h00;      memory[44567] <=  8'h00;      memory[44568] <=  8'h00;      memory[44569] <=  8'h00;      memory[44570] <=  8'h00;      memory[44571] <=  8'h00;      memory[44572] <=  8'h00;      memory[44573] <=  8'h00;      memory[44574] <=  8'h00;      memory[44575] <=  8'h00;      memory[44576] <=  8'h00;      memory[44577] <=  8'h00;      memory[44578] <=  8'h00;      memory[44579] <=  8'h00;      memory[44580] <=  8'h00;      memory[44581] <=  8'h00;      memory[44582] <=  8'h00;      memory[44583] <=  8'h00;      memory[44584] <=  8'h00;      memory[44585] <=  8'h00;      memory[44586] <=  8'h00;      memory[44587] <=  8'h00;      memory[44588] <=  8'h00;      memory[44589] <=  8'h00;      memory[44590] <=  8'h00;      memory[44591] <=  8'h00;      memory[44592] <=  8'h00;      memory[44593] <=  8'h00;      memory[44594] <=  8'h00;      memory[44595] <=  8'h00;      memory[44596] <=  8'h00;      memory[44597] <=  8'h00;      memory[44598] <=  8'h00;      memory[44599] <=  8'h00;      memory[44600] <=  8'h00;      memory[44601] <=  8'h00;      memory[44602] <=  8'h00;      memory[44603] <=  8'h00;      memory[44604] <=  8'h00;      memory[44605] <=  8'h00;      memory[44606] <=  8'h00;      memory[44607] <=  8'h00;      memory[44608] <=  8'h00;      memory[44609] <=  8'h00;      memory[44610] <=  8'h00;      memory[44611] <=  8'h00;      memory[44612] <=  8'h00;      memory[44613] <=  8'h00;      memory[44614] <=  8'h00;      memory[44615] <=  8'h00;      memory[44616] <=  8'h00;      memory[44617] <=  8'h00;      memory[44618] <=  8'h00;      memory[44619] <=  8'h00;      memory[44620] <=  8'h00;      memory[44621] <=  8'h00;      memory[44622] <=  8'h00;      memory[44623] <=  8'h00;      memory[44624] <=  8'h00;      memory[44625] <=  8'h00;      memory[44626] <=  8'h00;      memory[44627] <=  8'h00;      memory[44628] <=  8'h00;      memory[44629] <=  8'h00;      memory[44630] <=  8'h00;      memory[44631] <=  8'h00;      memory[44632] <=  8'h00;      memory[44633] <=  8'h00;      memory[44634] <=  8'h00;      memory[44635] <=  8'h00;      memory[44636] <=  8'h00;      memory[44637] <=  8'h00;      memory[44638] <=  8'h00;      memory[44639] <=  8'h00;      memory[44640] <=  8'h00;      memory[44641] <=  8'h00;      memory[44642] <=  8'h00;      memory[44643] <=  8'h00;      memory[44644] <=  8'h00;      memory[44645] <=  8'h00;      memory[44646] <=  8'h00;      memory[44647] <=  8'h00;      memory[44648] <=  8'h00;      memory[44649] <=  8'h00;      memory[44650] <=  8'h00;      memory[44651] <=  8'h00;      memory[44652] <=  8'h00;      memory[44653] <=  8'h00;      memory[44654] <=  8'h00;      memory[44655] <=  8'h00;      memory[44656] <=  8'h00;      memory[44657] <=  8'h00;      memory[44658] <=  8'h00;      memory[44659] <=  8'h00;      memory[44660] <=  8'h00;      memory[44661] <=  8'h00;      memory[44662] <=  8'h00;      memory[44663] <=  8'h00;      memory[44664] <=  8'h00;      memory[44665] <=  8'h00;      memory[44666] <=  8'h00;      memory[44667] <=  8'h00;      memory[44668] <=  8'h00;      memory[44669] <=  8'h00;      memory[44670] <=  8'h00;      memory[44671] <=  8'h00;      memory[44672] <=  8'h00;      memory[44673] <=  8'h00;      memory[44674] <=  8'h00;      memory[44675] <=  8'h00;      memory[44676] <=  8'h00;      memory[44677] <=  8'h00;      memory[44678] <=  8'h00;      memory[44679] <=  8'h00;      memory[44680] <=  8'h00;      memory[44681] <=  8'h00;      memory[44682] <=  8'h00;      memory[44683] <=  8'h00;      memory[44684] <=  8'h00;      memory[44685] <=  8'h00;      memory[44686] <=  8'h00;      memory[44687] <=  8'h00;      memory[44688] <=  8'h00;      memory[44689] <=  8'h00;      memory[44690] <=  8'h00;      memory[44691] <=  8'h00;      memory[44692] <=  8'h00;      memory[44693] <=  8'h00;      memory[44694] <=  8'h00;      memory[44695] <=  8'h00;      memory[44696] <=  8'h00;      memory[44697] <=  8'h00;      memory[44698] <=  8'h00;      memory[44699] <=  8'h00;      memory[44700] <=  8'h00;      memory[44701] <=  8'h00;      memory[44702] <=  8'h00;      memory[44703] <=  8'h00;      memory[44704] <=  8'h00;      memory[44705] <=  8'h00;      memory[44706] <=  8'h00;      memory[44707] <=  8'h00;      memory[44708] <=  8'h00;      memory[44709] <=  8'h00;      memory[44710] <=  8'h00;      memory[44711] <=  8'h00;      memory[44712] <=  8'h00;      memory[44713] <=  8'h00;      memory[44714] <=  8'h00;      memory[44715] <=  8'h00;      memory[44716] <=  8'h00;      memory[44717] <=  8'h00;      memory[44718] <=  8'h00;      memory[44719] <=  8'h00;      memory[44720] <=  8'h00;      memory[44721] <=  8'h00;      memory[44722] <=  8'h00;      memory[44723] <=  8'h00;      memory[44724] <=  8'h00;      memory[44725] <=  8'h00;      memory[44726] <=  8'h00;      memory[44727] <=  8'h00;      memory[44728] <=  8'h00;      memory[44729] <=  8'h00;      memory[44730] <=  8'h00;      memory[44731] <=  8'h00;      memory[44732] <=  8'h00;      memory[44733] <=  8'h00;      memory[44734] <=  8'h00;      memory[44735] <=  8'h00;      memory[44736] <=  8'h00;      memory[44737] <=  8'h00;      memory[44738] <=  8'h00;      memory[44739] <=  8'h00;      memory[44740] <=  8'h00;      memory[44741] <=  8'h00;      memory[44742] <=  8'h00;      memory[44743] <=  8'h00;      memory[44744] <=  8'h00;      memory[44745] <=  8'h00;      memory[44746] <=  8'h00;      memory[44747] <=  8'h00;      memory[44748] <=  8'h00;      memory[44749] <=  8'h00;      memory[44750] <=  8'h00;      memory[44751] <=  8'h00;      memory[44752] <=  8'h00;      memory[44753] <=  8'h00;      memory[44754] <=  8'h00;      memory[44755] <=  8'h00;      memory[44756] <=  8'h00;      memory[44757] <=  8'h00;      memory[44758] <=  8'h00;      memory[44759] <=  8'h00;      memory[44760] <=  8'h00;      memory[44761] <=  8'h00;      memory[44762] <=  8'h00;      memory[44763] <=  8'h00;      memory[44764] <=  8'h00;      memory[44765] <=  8'h00;      memory[44766] <=  8'h00;      memory[44767] <=  8'h00;      memory[44768] <=  8'h00;      memory[44769] <=  8'h00;      memory[44770] <=  8'h00;      memory[44771] <=  8'h00;      memory[44772] <=  8'h00;      memory[44773] <=  8'h00;      memory[44774] <=  8'h00;      memory[44775] <=  8'h00;      memory[44776] <=  8'h00;      memory[44777] <=  8'h00;      memory[44778] <=  8'h00;      memory[44779] <=  8'h00;      memory[44780] <=  8'h00;      memory[44781] <=  8'h00;      memory[44782] <=  8'h00;      memory[44783] <=  8'h00;      memory[44784] <=  8'h00;      memory[44785] <=  8'h00;      memory[44786] <=  8'h00;      memory[44787] <=  8'h00;      memory[44788] <=  8'h00;      memory[44789] <=  8'h00;      memory[44790] <=  8'h00;      memory[44791] <=  8'h00;      memory[44792] <=  8'h00;      memory[44793] <=  8'h00;      memory[44794] <=  8'h00;      memory[44795] <=  8'h00;      memory[44796] <=  8'h00;      memory[44797] <=  8'h00;      memory[44798] <=  8'h00;      memory[44799] <=  8'h00;      memory[44800] <=  8'h00;      memory[44801] <=  8'h00;      memory[44802] <=  8'h00;      memory[44803] <=  8'h00;      memory[44804] <=  8'h00;      memory[44805] <=  8'h00;      memory[44806] <=  8'h00;      memory[44807] <=  8'h00;      memory[44808] <=  8'h00;      memory[44809] <=  8'h00;      memory[44810] <=  8'h00;      memory[44811] <=  8'h00;      memory[44812] <=  8'h00;      memory[44813] <=  8'h00;      memory[44814] <=  8'h00;      memory[44815] <=  8'h00;      memory[44816] <=  8'h00;      memory[44817] <=  8'h00;      memory[44818] <=  8'h00;      memory[44819] <=  8'h00;      memory[44820] <=  8'h00;      memory[44821] <=  8'h00;      memory[44822] <=  8'h00;      memory[44823] <=  8'h00;      memory[44824] <=  8'h00;      memory[44825] <=  8'h00;      memory[44826] <=  8'h00;      memory[44827] <=  8'h00;      memory[44828] <=  8'h00;      memory[44829] <=  8'h00;      memory[44830] <=  8'h00;      memory[44831] <=  8'h00;      memory[44832] <=  8'h00;      memory[44833] <=  8'h00;      memory[44834] <=  8'h00;      memory[44835] <=  8'h00;      memory[44836] <=  8'h00;      memory[44837] <=  8'h00;      memory[44838] <=  8'h00;      memory[44839] <=  8'h00;      memory[44840] <=  8'h00;      memory[44841] <=  8'h00;      memory[44842] <=  8'h00;      memory[44843] <=  8'h00;      memory[44844] <=  8'h00;      memory[44845] <=  8'h00;      memory[44846] <=  8'h00;      memory[44847] <=  8'h00;      memory[44848] <=  8'h00;      memory[44849] <=  8'h00;      memory[44850] <=  8'h00;      memory[44851] <=  8'h00;      memory[44852] <=  8'h00;      memory[44853] <=  8'h00;      memory[44854] <=  8'h00;      memory[44855] <=  8'h00;      memory[44856] <=  8'h00;      memory[44857] <=  8'h00;      memory[44858] <=  8'h00;      memory[44859] <=  8'h00;      memory[44860] <=  8'h00;      memory[44861] <=  8'h00;      memory[44862] <=  8'h00;      memory[44863] <=  8'h00;      memory[44864] <=  8'h00;      memory[44865] <=  8'h00;      memory[44866] <=  8'h00;      memory[44867] <=  8'h00;      memory[44868] <=  8'h00;      memory[44869] <=  8'h00;      memory[44870] <=  8'h00;      memory[44871] <=  8'h00;      memory[44872] <=  8'h00;      memory[44873] <=  8'h00;      memory[44874] <=  8'h00;      memory[44875] <=  8'h00;      memory[44876] <=  8'h00;      memory[44877] <=  8'h00;      memory[44878] <=  8'h00;      memory[44879] <=  8'h00;      memory[44880] <=  8'h00;      memory[44881] <=  8'h00;      memory[44882] <=  8'h00;      memory[44883] <=  8'h00;      memory[44884] <=  8'h00;      memory[44885] <=  8'h00;      memory[44886] <=  8'h00;      memory[44887] <=  8'h00;      memory[44888] <=  8'h00;      memory[44889] <=  8'h00;      memory[44890] <=  8'h00;      memory[44891] <=  8'h00;      memory[44892] <=  8'h00;      memory[44893] <=  8'h00;      memory[44894] <=  8'h00;      memory[44895] <=  8'h00;      memory[44896] <=  8'h00;      memory[44897] <=  8'h00;      memory[44898] <=  8'h00;      memory[44899] <=  8'h00;      memory[44900] <=  8'h00;      memory[44901] <=  8'h00;      memory[44902] <=  8'h00;      memory[44903] <=  8'h00;      memory[44904] <=  8'h00;      memory[44905] <=  8'h00;      memory[44906] <=  8'h00;      memory[44907] <=  8'h00;      memory[44908] <=  8'h00;      memory[44909] <=  8'h00;      memory[44910] <=  8'h00;      memory[44911] <=  8'h00;      memory[44912] <=  8'h00;      memory[44913] <=  8'h00;      memory[44914] <=  8'h00;      memory[44915] <=  8'h00;      memory[44916] <=  8'h00;      memory[44917] <=  8'h00;      memory[44918] <=  8'h00;      memory[44919] <=  8'h00;      memory[44920] <=  8'h00;      memory[44921] <=  8'h00;      memory[44922] <=  8'h00;      memory[44923] <=  8'h00;      memory[44924] <=  8'h00;      memory[44925] <=  8'h00;      memory[44926] <=  8'h00;      memory[44927] <=  8'h00;      memory[44928] <=  8'h00;      memory[44929] <=  8'h00;      memory[44930] <=  8'h00;      memory[44931] <=  8'h00;      memory[44932] <=  8'h00;      memory[44933] <=  8'h00;      memory[44934] <=  8'h00;      memory[44935] <=  8'h00;      memory[44936] <=  8'h00;      memory[44937] <=  8'h00;      memory[44938] <=  8'h00;      memory[44939] <=  8'h00;      memory[44940] <=  8'h00;      memory[44941] <=  8'h00;      memory[44942] <=  8'h00;      memory[44943] <=  8'h00;      memory[44944] <=  8'h00;      memory[44945] <=  8'h00;      memory[44946] <=  8'h00;      memory[44947] <=  8'h00;      memory[44948] <=  8'h00;      memory[44949] <=  8'h00;      memory[44950] <=  8'h00;      memory[44951] <=  8'h00;      memory[44952] <=  8'h00;      memory[44953] <=  8'h00;      memory[44954] <=  8'h00;      memory[44955] <=  8'h00;      memory[44956] <=  8'h00;      memory[44957] <=  8'h00;      memory[44958] <=  8'h00;      memory[44959] <=  8'h00;      memory[44960] <=  8'h00;      memory[44961] <=  8'h00;      memory[44962] <=  8'h00;      memory[44963] <=  8'h00;      memory[44964] <=  8'h00;      memory[44965] <=  8'h00;      memory[44966] <=  8'h00;      memory[44967] <=  8'h00;      memory[44968] <=  8'h00;      memory[44969] <=  8'h00;      memory[44970] <=  8'h00;      memory[44971] <=  8'h00;      memory[44972] <=  8'h00;      memory[44973] <=  8'h00;      memory[44974] <=  8'h00;      memory[44975] <=  8'h00;      memory[44976] <=  8'h00;      memory[44977] <=  8'h00;      memory[44978] <=  8'h00;      memory[44979] <=  8'h00;      memory[44980] <=  8'h00;      memory[44981] <=  8'h00;      memory[44982] <=  8'h00;      memory[44983] <=  8'h00;      memory[44984] <=  8'h00;      memory[44985] <=  8'h00;      memory[44986] <=  8'h00;      memory[44987] <=  8'h00;      memory[44988] <=  8'h00;      memory[44989] <=  8'h00;      memory[44990] <=  8'h00;      memory[44991] <=  8'h00;      memory[44992] <=  8'h00;      memory[44993] <=  8'h00;      memory[44994] <=  8'h00;      memory[44995] <=  8'h00;      memory[44996] <=  8'h00;      memory[44997] <=  8'h00;      memory[44998] <=  8'h00;      memory[44999] <=  8'h00;      memory[45000] <=  8'h00;      memory[45001] <=  8'h00;      memory[45002] <=  8'h00;      memory[45003] <=  8'h00;      memory[45004] <=  8'h00;      memory[45005] <=  8'h00;      memory[45006] <=  8'h00;      memory[45007] <=  8'h00;      memory[45008] <=  8'h00;      memory[45009] <=  8'h00;      memory[45010] <=  8'h00;      memory[45011] <=  8'h00;      memory[45012] <=  8'h00;      memory[45013] <=  8'h00;      memory[45014] <=  8'h00;      memory[45015] <=  8'h00;      memory[45016] <=  8'h00;      memory[45017] <=  8'h00;      memory[45018] <=  8'h00;      memory[45019] <=  8'h00;      memory[45020] <=  8'h00;      memory[45021] <=  8'h00;      memory[45022] <=  8'h00;      memory[45023] <=  8'h00;      memory[45024] <=  8'h00;      memory[45025] <=  8'h00;      memory[45026] <=  8'h00;      memory[45027] <=  8'h00;      memory[45028] <=  8'h00;      memory[45029] <=  8'h00;      memory[45030] <=  8'h00;      memory[45031] <=  8'h00;      memory[45032] <=  8'h00;      memory[45033] <=  8'h00;      memory[45034] <=  8'h00;      memory[45035] <=  8'h00;      memory[45036] <=  8'h00;      memory[45037] <=  8'h00;      memory[45038] <=  8'h00;      memory[45039] <=  8'h00;      memory[45040] <=  8'h00;      memory[45041] <=  8'h00;      memory[45042] <=  8'h00;      memory[45043] <=  8'h00;      memory[45044] <=  8'h00;      memory[45045] <=  8'h00;      memory[45046] <=  8'h00;      memory[45047] <=  8'h00;      memory[45048] <=  8'h00;      memory[45049] <=  8'h00;      memory[45050] <=  8'h00;      memory[45051] <=  8'h00;      memory[45052] <=  8'h00;      memory[45053] <=  8'h00;      memory[45054] <=  8'h00;      memory[45055] <=  8'h00;      memory[45056] <=  8'h00;      memory[45057] <=  8'h00;      memory[45058] <=  8'h00;      memory[45059] <=  8'h00;      memory[45060] <=  8'h00;      memory[45061] <=  8'h00;      memory[45062] <=  8'h00;      memory[45063] <=  8'h00;      memory[45064] <=  8'h00;      memory[45065] <=  8'h00;      memory[45066] <=  8'h00;      memory[45067] <=  8'h00;      memory[45068] <=  8'h00;      memory[45069] <=  8'h00;      memory[45070] <=  8'h00;      memory[45071] <=  8'h00;      memory[45072] <=  8'h00;      memory[45073] <=  8'h00;      memory[45074] <=  8'h00;      memory[45075] <=  8'h00;      memory[45076] <=  8'h00;      memory[45077] <=  8'h00;      memory[45078] <=  8'h00;      memory[45079] <=  8'h00;      memory[45080] <=  8'h00;      memory[45081] <=  8'h00;      memory[45082] <=  8'h00;      memory[45083] <=  8'h00;      memory[45084] <=  8'h00;      memory[45085] <=  8'h00;      memory[45086] <=  8'h00;      memory[45087] <=  8'h00;      memory[45088] <=  8'h00;      memory[45089] <=  8'h00;      memory[45090] <=  8'h00;      memory[45091] <=  8'h00;      memory[45092] <=  8'h00;      memory[45093] <=  8'h00;      memory[45094] <=  8'h00;      memory[45095] <=  8'h00;      memory[45096] <=  8'h00;      memory[45097] <=  8'h00;      memory[45098] <=  8'h00;      memory[45099] <=  8'h00;      memory[45100] <=  8'h00;      memory[45101] <=  8'h00;      memory[45102] <=  8'h00;      memory[45103] <=  8'h00;      memory[45104] <=  8'h00;      memory[45105] <=  8'h00;      memory[45106] <=  8'h00;      memory[45107] <=  8'h00;      memory[45108] <=  8'h00;      memory[45109] <=  8'h00;      memory[45110] <=  8'h00;      memory[45111] <=  8'h00;      memory[45112] <=  8'h00;      memory[45113] <=  8'h00;      memory[45114] <=  8'h00;      memory[45115] <=  8'h00;      memory[45116] <=  8'h00;      memory[45117] <=  8'h00;      memory[45118] <=  8'h00;      memory[45119] <=  8'h00;      memory[45120] <=  8'h00;      memory[45121] <=  8'h00;      memory[45122] <=  8'h00;      memory[45123] <=  8'h00;      memory[45124] <=  8'h00;      memory[45125] <=  8'h00;      memory[45126] <=  8'h00;      memory[45127] <=  8'h00;      memory[45128] <=  8'h00;      memory[45129] <=  8'h00;      memory[45130] <=  8'h00;      memory[45131] <=  8'h00;      memory[45132] <=  8'h00;      memory[45133] <=  8'h00;      memory[45134] <=  8'h00;      memory[45135] <=  8'h00;      memory[45136] <=  8'h00;      memory[45137] <=  8'h00;      memory[45138] <=  8'h00;      memory[45139] <=  8'h00;      memory[45140] <=  8'h00;      memory[45141] <=  8'h00;      memory[45142] <=  8'h00;      memory[45143] <=  8'h00;      memory[45144] <=  8'h00;      memory[45145] <=  8'h00;      memory[45146] <=  8'h00;      memory[45147] <=  8'h00;      memory[45148] <=  8'h00;      memory[45149] <=  8'h00;      memory[45150] <=  8'h00;      memory[45151] <=  8'h00;      memory[45152] <=  8'h00;      memory[45153] <=  8'h00;      memory[45154] <=  8'h00;      memory[45155] <=  8'h00;      memory[45156] <=  8'h00;      memory[45157] <=  8'h00;      memory[45158] <=  8'h00;      memory[45159] <=  8'h00;      memory[45160] <=  8'h00;      memory[45161] <=  8'h00;      memory[45162] <=  8'h00;      memory[45163] <=  8'h00;      memory[45164] <=  8'h00;      memory[45165] <=  8'h00;      memory[45166] <=  8'h00;      memory[45167] <=  8'h00;      memory[45168] <=  8'h00;      memory[45169] <=  8'h00;      memory[45170] <=  8'h00;      memory[45171] <=  8'h00;      memory[45172] <=  8'h00;      memory[45173] <=  8'h00;      memory[45174] <=  8'h00;      memory[45175] <=  8'h00;      memory[45176] <=  8'h00;      memory[45177] <=  8'h00;      memory[45178] <=  8'h00;      memory[45179] <=  8'h00;      memory[45180] <=  8'h00;      memory[45181] <=  8'h00;      memory[45182] <=  8'h00;      memory[45183] <=  8'h00;      memory[45184] <=  8'h00;      memory[45185] <=  8'h00;      memory[45186] <=  8'h00;      memory[45187] <=  8'h00;      memory[45188] <=  8'h00;      memory[45189] <=  8'h00;      memory[45190] <=  8'h00;      memory[45191] <=  8'h00;      memory[45192] <=  8'h00;      memory[45193] <=  8'h00;      memory[45194] <=  8'h00;      memory[45195] <=  8'h00;      memory[45196] <=  8'h00;      memory[45197] <=  8'h00;      memory[45198] <=  8'h00;      memory[45199] <=  8'h00;      memory[45200] <=  8'h00;      memory[45201] <=  8'h00;      memory[45202] <=  8'h00;      memory[45203] <=  8'h00;      memory[45204] <=  8'h00;      memory[45205] <=  8'h00;      memory[45206] <=  8'h00;      memory[45207] <=  8'h00;      memory[45208] <=  8'h00;      memory[45209] <=  8'h00;      memory[45210] <=  8'h00;      memory[45211] <=  8'h00;      memory[45212] <=  8'h00;      memory[45213] <=  8'h00;      memory[45214] <=  8'h00;      memory[45215] <=  8'h00;      memory[45216] <=  8'h00;      memory[45217] <=  8'h00;      memory[45218] <=  8'h00;      memory[45219] <=  8'h00;      memory[45220] <=  8'h00;      memory[45221] <=  8'h00;      memory[45222] <=  8'h00;      memory[45223] <=  8'h00;      memory[45224] <=  8'h00;      memory[45225] <=  8'h00;      memory[45226] <=  8'h00;      memory[45227] <=  8'h00;      memory[45228] <=  8'h00;      memory[45229] <=  8'h00;      memory[45230] <=  8'h00;      memory[45231] <=  8'h00;      memory[45232] <=  8'h00;      memory[45233] <=  8'h00;      memory[45234] <=  8'h00;      memory[45235] <=  8'h00;      memory[45236] <=  8'h00;      memory[45237] <=  8'h00;      memory[45238] <=  8'h00;      memory[45239] <=  8'h00;      memory[45240] <=  8'h00;      memory[45241] <=  8'h00;      memory[45242] <=  8'h00;      memory[45243] <=  8'h00;      memory[45244] <=  8'h00;      memory[45245] <=  8'h00;      memory[45246] <=  8'h00;      memory[45247] <=  8'h00;      memory[45248] <=  8'h00;      memory[45249] <=  8'h00;      memory[45250] <=  8'h00;      memory[45251] <=  8'h00;      memory[45252] <=  8'h00;      memory[45253] <=  8'h00;      memory[45254] <=  8'h00;      memory[45255] <=  8'h00;      memory[45256] <=  8'h00;      memory[45257] <=  8'h00;      memory[45258] <=  8'h00;      memory[45259] <=  8'h00;      memory[45260] <=  8'h00;      memory[45261] <=  8'h00;      memory[45262] <=  8'h00;      memory[45263] <=  8'h00;      memory[45264] <=  8'h00;      memory[45265] <=  8'h00;      memory[45266] <=  8'h00;      memory[45267] <=  8'h00;      memory[45268] <=  8'h00;      memory[45269] <=  8'h00;      memory[45270] <=  8'h00;      memory[45271] <=  8'h00;      memory[45272] <=  8'h00;      memory[45273] <=  8'h00;      memory[45274] <=  8'h00;      memory[45275] <=  8'h00;      memory[45276] <=  8'h00;      memory[45277] <=  8'h00;      memory[45278] <=  8'h00;      memory[45279] <=  8'h00;      memory[45280] <=  8'h00;      memory[45281] <=  8'h00;      memory[45282] <=  8'h00;      memory[45283] <=  8'h00;      memory[45284] <=  8'h00;      memory[45285] <=  8'h00;      memory[45286] <=  8'h00;      memory[45287] <=  8'h00;      memory[45288] <=  8'h00;      memory[45289] <=  8'h00;      memory[45290] <=  8'h00;      memory[45291] <=  8'h00;      memory[45292] <=  8'h00;      memory[45293] <=  8'h00;      memory[45294] <=  8'h00;      memory[45295] <=  8'h00;      memory[45296] <=  8'h00;      memory[45297] <=  8'h00;      memory[45298] <=  8'h00;      memory[45299] <=  8'h00;      memory[45300] <=  8'h00;      memory[45301] <=  8'h00;      memory[45302] <=  8'h00;      memory[45303] <=  8'h00;      memory[45304] <=  8'h00;      memory[45305] <=  8'h00;      memory[45306] <=  8'h00;      memory[45307] <=  8'h00;      memory[45308] <=  8'h00;      memory[45309] <=  8'h00;      memory[45310] <=  8'h00;      memory[45311] <=  8'h00;      memory[45312] <=  8'h00;      memory[45313] <=  8'h00;      memory[45314] <=  8'h00;      memory[45315] <=  8'h00;      memory[45316] <=  8'h00;      memory[45317] <=  8'h00;      memory[45318] <=  8'h00;      memory[45319] <=  8'h00;      memory[45320] <=  8'h00;      memory[45321] <=  8'h00;      memory[45322] <=  8'h00;      memory[45323] <=  8'h00;      memory[45324] <=  8'h00;      memory[45325] <=  8'h00;      memory[45326] <=  8'h00;      memory[45327] <=  8'h00;      memory[45328] <=  8'h00;      memory[45329] <=  8'h00;      memory[45330] <=  8'h00;      memory[45331] <=  8'h00;      memory[45332] <=  8'h00;      memory[45333] <=  8'h00;      memory[45334] <=  8'h00;      memory[45335] <=  8'h00;      memory[45336] <=  8'h00;      memory[45337] <=  8'h00;      memory[45338] <=  8'h00;      memory[45339] <=  8'h00;      memory[45340] <=  8'h00;      memory[45341] <=  8'h00;      memory[45342] <=  8'h00;      memory[45343] <=  8'h00;      memory[45344] <=  8'h00;      memory[45345] <=  8'h00;      memory[45346] <=  8'h00;      memory[45347] <=  8'h00;      memory[45348] <=  8'h00;      memory[45349] <=  8'h00;      memory[45350] <=  8'h00;      memory[45351] <=  8'h00;      memory[45352] <=  8'h00;      memory[45353] <=  8'h00;      memory[45354] <=  8'h00;      memory[45355] <=  8'h00;      memory[45356] <=  8'h00;      memory[45357] <=  8'h00;      memory[45358] <=  8'h00;      memory[45359] <=  8'h00;      memory[45360] <=  8'h00;      memory[45361] <=  8'h00;      memory[45362] <=  8'h00;      memory[45363] <=  8'h00;      memory[45364] <=  8'h00;      memory[45365] <=  8'h00;      memory[45366] <=  8'h00;      memory[45367] <=  8'h00;      memory[45368] <=  8'h00;      memory[45369] <=  8'h00;      memory[45370] <=  8'h00;      memory[45371] <=  8'h00;      memory[45372] <=  8'h00;      memory[45373] <=  8'h00;      memory[45374] <=  8'h00;      memory[45375] <=  8'h00;      memory[45376] <=  8'h00;      memory[45377] <=  8'h00;      memory[45378] <=  8'h00;      memory[45379] <=  8'h00;      memory[45380] <=  8'h00;      memory[45381] <=  8'h00;      memory[45382] <=  8'h00;      memory[45383] <=  8'h00;      memory[45384] <=  8'h00;      memory[45385] <=  8'h00;      memory[45386] <=  8'h00;      memory[45387] <=  8'h00;      memory[45388] <=  8'h00;      memory[45389] <=  8'h00;      memory[45390] <=  8'h00;      memory[45391] <=  8'h00;      memory[45392] <=  8'h00;      memory[45393] <=  8'h00;      memory[45394] <=  8'h00;      memory[45395] <=  8'h00;      memory[45396] <=  8'h00;      memory[45397] <=  8'h00;      memory[45398] <=  8'h00;      memory[45399] <=  8'h00;      memory[45400] <=  8'h00;      memory[45401] <=  8'h00;      memory[45402] <=  8'h00;      memory[45403] <=  8'h00;      memory[45404] <=  8'h00;      memory[45405] <=  8'h00;      memory[45406] <=  8'h00;      memory[45407] <=  8'h00;      memory[45408] <=  8'h00;      memory[45409] <=  8'h00;      memory[45410] <=  8'h00;      memory[45411] <=  8'h00;      memory[45412] <=  8'h00;      memory[45413] <=  8'h00;      memory[45414] <=  8'h00;      memory[45415] <=  8'h00;      memory[45416] <=  8'h00;      memory[45417] <=  8'h00;      memory[45418] <=  8'h00;      memory[45419] <=  8'h00;      memory[45420] <=  8'h00;      memory[45421] <=  8'h00;      memory[45422] <=  8'h00;      memory[45423] <=  8'h00;      memory[45424] <=  8'h00;      memory[45425] <=  8'h00;      memory[45426] <=  8'h00;      memory[45427] <=  8'h00;      memory[45428] <=  8'h00;      memory[45429] <=  8'h00;      memory[45430] <=  8'h00;      memory[45431] <=  8'h00;      memory[45432] <=  8'h00;      memory[45433] <=  8'h00;      memory[45434] <=  8'h00;      memory[45435] <=  8'h00;      memory[45436] <=  8'h00;      memory[45437] <=  8'h00;      memory[45438] <=  8'h00;      memory[45439] <=  8'h00;      memory[45440] <=  8'h00;      memory[45441] <=  8'h00;      memory[45442] <=  8'h00;      memory[45443] <=  8'h00;      memory[45444] <=  8'h00;      memory[45445] <=  8'h00;      memory[45446] <=  8'h00;      memory[45447] <=  8'h00;      memory[45448] <=  8'h00;      memory[45449] <=  8'h00;      memory[45450] <=  8'h00;      memory[45451] <=  8'h00;      memory[45452] <=  8'h00;      memory[45453] <=  8'h00;      memory[45454] <=  8'h00;      memory[45455] <=  8'h00;      memory[45456] <=  8'h00;      memory[45457] <=  8'h00;      memory[45458] <=  8'h00;      memory[45459] <=  8'h00;      memory[45460] <=  8'h00;      memory[45461] <=  8'h00;      memory[45462] <=  8'h00;      memory[45463] <=  8'h00;      memory[45464] <=  8'h00;      memory[45465] <=  8'h00;      memory[45466] <=  8'h00;      memory[45467] <=  8'h00;      memory[45468] <=  8'h00;      memory[45469] <=  8'h00;      memory[45470] <=  8'h00;      memory[45471] <=  8'h00;      memory[45472] <=  8'h00;      memory[45473] <=  8'h00;      memory[45474] <=  8'h00;      memory[45475] <=  8'h00;      memory[45476] <=  8'h00;      memory[45477] <=  8'h00;      memory[45478] <=  8'h00;      memory[45479] <=  8'h00;      memory[45480] <=  8'h00;      memory[45481] <=  8'h00;      memory[45482] <=  8'h00;      memory[45483] <=  8'h00;      memory[45484] <=  8'h00;      memory[45485] <=  8'h00;      memory[45486] <=  8'h00;      memory[45487] <=  8'h00;      memory[45488] <=  8'h00;      memory[45489] <=  8'h00;      memory[45490] <=  8'h00;      memory[45491] <=  8'h00;      memory[45492] <=  8'h00;      memory[45493] <=  8'h00;      memory[45494] <=  8'h00;      memory[45495] <=  8'h00;      memory[45496] <=  8'h00;      memory[45497] <=  8'h00;      memory[45498] <=  8'h00;      memory[45499] <=  8'h00;      memory[45500] <=  8'h00;      memory[45501] <=  8'h00;      memory[45502] <=  8'h00;      memory[45503] <=  8'h00;      memory[45504] <=  8'h00;      memory[45505] <=  8'h00;      memory[45506] <=  8'h00;      memory[45507] <=  8'h00;      memory[45508] <=  8'h00;      memory[45509] <=  8'h00;      memory[45510] <=  8'h00;      memory[45511] <=  8'h00;      memory[45512] <=  8'h00;      memory[45513] <=  8'h00;      memory[45514] <=  8'h00;      memory[45515] <=  8'h00;      memory[45516] <=  8'h00;      memory[45517] <=  8'h00;      memory[45518] <=  8'h00;      memory[45519] <=  8'h00;      memory[45520] <=  8'h00;      memory[45521] <=  8'h00;      memory[45522] <=  8'h00;      memory[45523] <=  8'h00;      memory[45524] <=  8'h00;      memory[45525] <=  8'h00;      memory[45526] <=  8'h00;      memory[45527] <=  8'h00;      memory[45528] <=  8'h00;      memory[45529] <=  8'h00;      memory[45530] <=  8'h00;      memory[45531] <=  8'h00;      memory[45532] <=  8'h00;      memory[45533] <=  8'h00;      memory[45534] <=  8'h00;      memory[45535] <=  8'h00;      memory[45536] <=  8'h00;      memory[45537] <=  8'h00;      memory[45538] <=  8'h00;      memory[45539] <=  8'h00;      memory[45540] <=  8'h00;      memory[45541] <=  8'h00;      memory[45542] <=  8'h00;      memory[45543] <=  8'h00;      memory[45544] <=  8'h00;      memory[45545] <=  8'h00;      memory[45546] <=  8'h00;      memory[45547] <=  8'h00;      memory[45548] <=  8'h00;      memory[45549] <=  8'h00;      memory[45550] <=  8'h00;      memory[45551] <=  8'h00;      memory[45552] <=  8'h00;      memory[45553] <=  8'h00;      memory[45554] <=  8'h00;      memory[45555] <=  8'h00;      memory[45556] <=  8'h00;      memory[45557] <=  8'h00;      memory[45558] <=  8'h00;      memory[45559] <=  8'h00;      memory[45560] <=  8'h00;      memory[45561] <=  8'h00;      memory[45562] <=  8'h00;      memory[45563] <=  8'h00;      memory[45564] <=  8'h00;      memory[45565] <=  8'h00;      memory[45566] <=  8'h00;      memory[45567] <=  8'h00;      memory[45568] <=  8'h00;      memory[45569] <=  8'h00;      memory[45570] <=  8'h00;      memory[45571] <=  8'h00;      memory[45572] <=  8'h00;      memory[45573] <=  8'h00;      memory[45574] <=  8'h00;      memory[45575] <=  8'h00;      memory[45576] <=  8'h00;      memory[45577] <=  8'h00;      memory[45578] <=  8'h00;      memory[45579] <=  8'h00;      memory[45580] <=  8'h00;      memory[45581] <=  8'h00;      memory[45582] <=  8'h00;      memory[45583] <=  8'h00;      memory[45584] <=  8'h00;      memory[45585] <=  8'h00;      memory[45586] <=  8'h00;      memory[45587] <=  8'h00;      memory[45588] <=  8'h00;      memory[45589] <=  8'h00;      memory[45590] <=  8'h00;      memory[45591] <=  8'h00;      memory[45592] <=  8'h00;      memory[45593] <=  8'h00;      memory[45594] <=  8'h00;      memory[45595] <=  8'h00;      memory[45596] <=  8'h00;      memory[45597] <=  8'h00;      memory[45598] <=  8'h00;      memory[45599] <=  8'h00;      memory[45600] <=  8'h00;      memory[45601] <=  8'h00;      memory[45602] <=  8'h00;      memory[45603] <=  8'h00;      memory[45604] <=  8'h00;      memory[45605] <=  8'h00;      memory[45606] <=  8'h00;      memory[45607] <=  8'h00;      memory[45608] <=  8'h00;      memory[45609] <=  8'h00;      memory[45610] <=  8'h00;      memory[45611] <=  8'h00;      memory[45612] <=  8'h00;      memory[45613] <=  8'h00;      memory[45614] <=  8'h00;      memory[45615] <=  8'h00;      memory[45616] <=  8'h00;      memory[45617] <=  8'h00;      memory[45618] <=  8'h00;      memory[45619] <=  8'h00;      memory[45620] <=  8'h00;      memory[45621] <=  8'h00;      memory[45622] <=  8'h00;      memory[45623] <=  8'h00;      memory[45624] <=  8'h00;      memory[45625] <=  8'h00;      memory[45626] <=  8'h00;      memory[45627] <=  8'h00;      memory[45628] <=  8'h00;      memory[45629] <=  8'h00;      memory[45630] <=  8'h00;      memory[45631] <=  8'h00;      memory[45632] <=  8'h00;      memory[45633] <=  8'h00;      memory[45634] <=  8'h00;      memory[45635] <=  8'h00;      memory[45636] <=  8'h00;      memory[45637] <=  8'h00;      memory[45638] <=  8'h00;      memory[45639] <=  8'h00;      memory[45640] <=  8'h00;      memory[45641] <=  8'h00;      memory[45642] <=  8'h00;      memory[45643] <=  8'h00;      memory[45644] <=  8'h00;      memory[45645] <=  8'h00;      memory[45646] <=  8'h00;      memory[45647] <=  8'h00;      memory[45648] <=  8'h00;      memory[45649] <=  8'h00;      memory[45650] <=  8'h00;      memory[45651] <=  8'h00;      memory[45652] <=  8'h00;      memory[45653] <=  8'h00;      memory[45654] <=  8'h00;      memory[45655] <=  8'h00;      memory[45656] <=  8'h00;      memory[45657] <=  8'h00;      memory[45658] <=  8'h00;      memory[45659] <=  8'h00;      memory[45660] <=  8'h00;      memory[45661] <=  8'h00;      memory[45662] <=  8'h00;      memory[45663] <=  8'h00;      memory[45664] <=  8'h00;      memory[45665] <=  8'h00;      memory[45666] <=  8'h00;      memory[45667] <=  8'h00;      memory[45668] <=  8'h00;      memory[45669] <=  8'h00;      memory[45670] <=  8'h00;      memory[45671] <=  8'h00;      memory[45672] <=  8'h00;      memory[45673] <=  8'h00;      memory[45674] <=  8'h00;      memory[45675] <=  8'h00;      memory[45676] <=  8'h00;      memory[45677] <=  8'h00;      memory[45678] <=  8'h00;      memory[45679] <=  8'h00;      memory[45680] <=  8'h00;      memory[45681] <=  8'h00;      memory[45682] <=  8'h00;      memory[45683] <=  8'h00;      memory[45684] <=  8'h00;      memory[45685] <=  8'h00;      memory[45686] <=  8'h00;      memory[45687] <=  8'h00;      memory[45688] <=  8'h00;      memory[45689] <=  8'h00;      memory[45690] <=  8'h00;      memory[45691] <=  8'h00;      memory[45692] <=  8'h00;      memory[45693] <=  8'h00;      memory[45694] <=  8'h00;      memory[45695] <=  8'h00;      memory[45696] <=  8'h00;      memory[45697] <=  8'h00;      memory[45698] <=  8'h00;      memory[45699] <=  8'h00;      memory[45700] <=  8'h00;      memory[45701] <=  8'h00;      memory[45702] <=  8'h00;      memory[45703] <=  8'h00;      memory[45704] <=  8'h00;      memory[45705] <=  8'h00;      memory[45706] <=  8'h00;      memory[45707] <=  8'h00;      memory[45708] <=  8'h00;      memory[45709] <=  8'h00;      memory[45710] <=  8'h00;      memory[45711] <=  8'h00;      memory[45712] <=  8'h00;      memory[45713] <=  8'h00;      memory[45714] <=  8'h00;      memory[45715] <=  8'h00;      memory[45716] <=  8'h00;      memory[45717] <=  8'h00;      memory[45718] <=  8'h00;      memory[45719] <=  8'h00;      memory[45720] <=  8'h00;      memory[45721] <=  8'h00;      memory[45722] <=  8'h00;      memory[45723] <=  8'h00;      memory[45724] <=  8'h00;      memory[45725] <=  8'h00;      memory[45726] <=  8'h00;      memory[45727] <=  8'h00;      memory[45728] <=  8'h00;      memory[45729] <=  8'h00;      memory[45730] <=  8'h00;      memory[45731] <=  8'h00;      memory[45732] <=  8'h00;      memory[45733] <=  8'h00;      memory[45734] <=  8'h00;      memory[45735] <=  8'h00;      memory[45736] <=  8'h00;      memory[45737] <=  8'h00;      memory[45738] <=  8'h00;      memory[45739] <=  8'h00;      memory[45740] <=  8'h00;      memory[45741] <=  8'h00;      memory[45742] <=  8'h00;      memory[45743] <=  8'h00;      memory[45744] <=  8'h00;      memory[45745] <=  8'h00;      memory[45746] <=  8'h00;      memory[45747] <=  8'h00;      memory[45748] <=  8'h00;      memory[45749] <=  8'h00;      memory[45750] <=  8'h00;      memory[45751] <=  8'h00;      memory[45752] <=  8'h00;      memory[45753] <=  8'h00;      memory[45754] <=  8'h00;      memory[45755] <=  8'h00;      memory[45756] <=  8'h00;      memory[45757] <=  8'h00;      memory[45758] <=  8'h00;      memory[45759] <=  8'h00;      memory[45760] <=  8'h00;      memory[45761] <=  8'h00;      memory[45762] <=  8'h00;      memory[45763] <=  8'h00;      memory[45764] <=  8'h00;      memory[45765] <=  8'h00;      memory[45766] <=  8'h00;      memory[45767] <=  8'h00;      memory[45768] <=  8'h00;      memory[45769] <=  8'h00;      memory[45770] <=  8'h00;      memory[45771] <=  8'h00;      memory[45772] <=  8'h00;      memory[45773] <=  8'h00;      memory[45774] <=  8'h00;      memory[45775] <=  8'h00;      memory[45776] <=  8'h00;      memory[45777] <=  8'h00;      memory[45778] <=  8'h00;      memory[45779] <=  8'h00;      memory[45780] <=  8'h00;      memory[45781] <=  8'h00;      memory[45782] <=  8'h00;      memory[45783] <=  8'h00;      memory[45784] <=  8'h00;      memory[45785] <=  8'h00;      memory[45786] <=  8'h00;      memory[45787] <=  8'h00;      memory[45788] <=  8'h00;      memory[45789] <=  8'h00;      memory[45790] <=  8'h00;      memory[45791] <=  8'h00;      memory[45792] <=  8'h00;      memory[45793] <=  8'h00;      memory[45794] <=  8'h00;      memory[45795] <=  8'h00;      memory[45796] <=  8'h00;      memory[45797] <=  8'h00;      memory[45798] <=  8'h00;      memory[45799] <=  8'h00;      memory[45800] <=  8'h00;      memory[45801] <=  8'h00;      memory[45802] <=  8'h00;      memory[45803] <=  8'h00;      memory[45804] <=  8'h00;      memory[45805] <=  8'h00;      memory[45806] <=  8'h00;      memory[45807] <=  8'h00;      memory[45808] <=  8'h00;      memory[45809] <=  8'h00;      memory[45810] <=  8'h00;      memory[45811] <=  8'h00;      memory[45812] <=  8'h00;      memory[45813] <=  8'h00;      memory[45814] <=  8'h00;      memory[45815] <=  8'h00;      memory[45816] <=  8'h00;      memory[45817] <=  8'h00;      memory[45818] <=  8'h00;      memory[45819] <=  8'h00;      memory[45820] <=  8'h00;      memory[45821] <=  8'h00;      memory[45822] <=  8'h00;      memory[45823] <=  8'h00;      memory[45824] <=  8'h00;      memory[45825] <=  8'h00;      memory[45826] <=  8'h00;      memory[45827] <=  8'h00;      memory[45828] <=  8'h00;      memory[45829] <=  8'h00;      memory[45830] <=  8'h00;      memory[45831] <=  8'h00;      memory[45832] <=  8'h00;      memory[45833] <=  8'h00;      memory[45834] <=  8'h00;      memory[45835] <=  8'h00;      memory[45836] <=  8'h00;      memory[45837] <=  8'h00;      memory[45838] <=  8'h00;      memory[45839] <=  8'h00;      memory[45840] <=  8'h00;      memory[45841] <=  8'h00;      memory[45842] <=  8'h00;      memory[45843] <=  8'h00;      memory[45844] <=  8'h00;      memory[45845] <=  8'h00;      memory[45846] <=  8'h00;      memory[45847] <=  8'h00;      memory[45848] <=  8'h00;      memory[45849] <=  8'h00;      memory[45850] <=  8'h00;      memory[45851] <=  8'h00;      memory[45852] <=  8'h00;      memory[45853] <=  8'h00;      memory[45854] <=  8'h00;      memory[45855] <=  8'h00;      memory[45856] <=  8'h00;      memory[45857] <=  8'h00;      memory[45858] <=  8'h00;      memory[45859] <=  8'h00;      memory[45860] <=  8'h00;      memory[45861] <=  8'h00;      memory[45862] <=  8'h00;      memory[45863] <=  8'h00;      memory[45864] <=  8'h00;      memory[45865] <=  8'h00;      memory[45866] <=  8'h00;      memory[45867] <=  8'h00;      memory[45868] <=  8'h00;      memory[45869] <=  8'h00;      memory[45870] <=  8'h00;      memory[45871] <=  8'h00;      memory[45872] <=  8'h00;      memory[45873] <=  8'h00;      memory[45874] <=  8'h00;      memory[45875] <=  8'h00;      memory[45876] <=  8'h00;      memory[45877] <=  8'h00;      memory[45878] <=  8'h00;      memory[45879] <=  8'h00;      memory[45880] <=  8'h00;      memory[45881] <=  8'h00;      memory[45882] <=  8'h00;      memory[45883] <=  8'h00;      memory[45884] <=  8'h00;      memory[45885] <=  8'h00;      memory[45886] <=  8'h00;      memory[45887] <=  8'h00;      memory[45888] <=  8'h00;      memory[45889] <=  8'h00;      memory[45890] <=  8'h00;      memory[45891] <=  8'h00;      memory[45892] <=  8'h00;      memory[45893] <=  8'h00;      memory[45894] <=  8'h00;      memory[45895] <=  8'h00;      memory[45896] <=  8'h00;      memory[45897] <=  8'h00;      memory[45898] <=  8'h00;      memory[45899] <=  8'h00;      memory[45900] <=  8'h00;      memory[45901] <=  8'h00;      memory[45902] <=  8'h00;      memory[45903] <=  8'h00;      memory[45904] <=  8'h00;      memory[45905] <=  8'h00;      memory[45906] <=  8'h00;      memory[45907] <=  8'h00;      memory[45908] <=  8'h00;      memory[45909] <=  8'h00;      memory[45910] <=  8'h00;      memory[45911] <=  8'h00;      memory[45912] <=  8'h00;      memory[45913] <=  8'h00;      memory[45914] <=  8'h00;      memory[45915] <=  8'h00;      memory[45916] <=  8'h00;      memory[45917] <=  8'h00;      memory[45918] <=  8'h00;      memory[45919] <=  8'h00;      memory[45920] <=  8'h00;      memory[45921] <=  8'h00;      memory[45922] <=  8'h00;      memory[45923] <=  8'h00;      memory[45924] <=  8'h00;      memory[45925] <=  8'h00;      memory[45926] <=  8'h00;      memory[45927] <=  8'h00;      memory[45928] <=  8'h00;      memory[45929] <=  8'h00;      memory[45930] <=  8'h00;      memory[45931] <=  8'h00;      memory[45932] <=  8'h00;      memory[45933] <=  8'h00;      memory[45934] <=  8'h00;      memory[45935] <=  8'h00;      memory[45936] <=  8'h00;      memory[45937] <=  8'h00;      memory[45938] <=  8'h00;      memory[45939] <=  8'h00;      memory[45940] <=  8'h00;      memory[45941] <=  8'h00;      memory[45942] <=  8'h00;      memory[45943] <=  8'h00;      memory[45944] <=  8'h00;      memory[45945] <=  8'h00;      memory[45946] <=  8'h00;      memory[45947] <=  8'h00;      memory[45948] <=  8'h00;      memory[45949] <=  8'h00;      memory[45950] <=  8'h00;      memory[45951] <=  8'h00;      memory[45952] <=  8'h00;      memory[45953] <=  8'h00;      memory[45954] <=  8'h00;      memory[45955] <=  8'h00;      memory[45956] <=  8'h00;      memory[45957] <=  8'h00;      memory[45958] <=  8'h00;      memory[45959] <=  8'h00;      memory[45960] <=  8'h00;      memory[45961] <=  8'h00;      memory[45962] <=  8'h00;      memory[45963] <=  8'h00;      memory[45964] <=  8'h00;      memory[45965] <=  8'h00;      memory[45966] <=  8'h00;      memory[45967] <=  8'h00;      memory[45968] <=  8'h00;      memory[45969] <=  8'h00;      memory[45970] <=  8'h00;      memory[45971] <=  8'h00;      memory[45972] <=  8'h00;      memory[45973] <=  8'h00;      memory[45974] <=  8'h00;      memory[45975] <=  8'h00;      memory[45976] <=  8'h00;      memory[45977] <=  8'h00;      memory[45978] <=  8'h00;      memory[45979] <=  8'h00;      memory[45980] <=  8'h00;      memory[45981] <=  8'h00;      memory[45982] <=  8'h00;      memory[45983] <=  8'h00;      memory[45984] <=  8'h00;      memory[45985] <=  8'h00;      memory[45986] <=  8'h00;      memory[45987] <=  8'h00;      memory[45988] <=  8'h00;      memory[45989] <=  8'h00;      memory[45990] <=  8'h00;      memory[45991] <=  8'h00;      memory[45992] <=  8'h00;      memory[45993] <=  8'h00;      memory[45994] <=  8'h00;      memory[45995] <=  8'h00;      memory[45996] <=  8'h00;      memory[45997] <=  8'h00;      memory[45998] <=  8'h00;      memory[45999] <=  8'h00;      memory[46000] <=  8'h00;      memory[46001] <=  8'h00;      memory[46002] <=  8'h00;      memory[46003] <=  8'h00;      memory[46004] <=  8'h00;      memory[46005] <=  8'h00;      memory[46006] <=  8'h00;      memory[46007] <=  8'h00;      memory[46008] <=  8'h00;      memory[46009] <=  8'h00;      memory[46010] <=  8'h00;      memory[46011] <=  8'h00;      memory[46012] <=  8'h00;      memory[46013] <=  8'h00;      memory[46014] <=  8'h00;      memory[46015] <=  8'h00;      memory[46016] <=  8'h00;      memory[46017] <=  8'h00;      memory[46018] <=  8'h00;      memory[46019] <=  8'h00;      memory[46020] <=  8'h00;      memory[46021] <=  8'h00;      memory[46022] <=  8'h00;      memory[46023] <=  8'h00;      memory[46024] <=  8'h00;      memory[46025] <=  8'h00;      memory[46026] <=  8'h00;      memory[46027] <=  8'h00;      memory[46028] <=  8'h00;      memory[46029] <=  8'h00;      memory[46030] <=  8'h00;      memory[46031] <=  8'h00;      memory[46032] <=  8'h00;      memory[46033] <=  8'h00;      memory[46034] <=  8'h00;      memory[46035] <=  8'h00;      memory[46036] <=  8'h00;      memory[46037] <=  8'h00;      memory[46038] <=  8'h00;      memory[46039] <=  8'h00;      memory[46040] <=  8'h00;      memory[46041] <=  8'h00;      memory[46042] <=  8'h00;      memory[46043] <=  8'h00;      memory[46044] <=  8'h00;      memory[46045] <=  8'h00;      memory[46046] <=  8'h00;      memory[46047] <=  8'h00;      memory[46048] <=  8'h00;      memory[46049] <=  8'h00;      memory[46050] <=  8'h00;      memory[46051] <=  8'h00;      memory[46052] <=  8'h00;      memory[46053] <=  8'h00;      memory[46054] <=  8'h00;      memory[46055] <=  8'h00;      memory[46056] <=  8'h00;      memory[46057] <=  8'h00;      memory[46058] <=  8'h00;      memory[46059] <=  8'h00;      memory[46060] <=  8'h00;      memory[46061] <=  8'h00;      memory[46062] <=  8'h00;      memory[46063] <=  8'h00;      memory[46064] <=  8'h00;      memory[46065] <=  8'h00;      memory[46066] <=  8'h00;      memory[46067] <=  8'h00;      memory[46068] <=  8'h00;      memory[46069] <=  8'h00;      memory[46070] <=  8'h00;      memory[46071] <=  8'h00;      memory[46072] <=  8'h00;      memory[46073] <=  8'h00;      memory[46074] <=  8'h00;      memory[46075] <=  8'h00;      memory[46076] <=  8'h00;      memory[46077] <=  8'h00;      memory[46078] <=  8'h00;      memory[46079] <=  8'h00;      memory[46080] <=  8'h00;      memory[46081] <=  8'h00;      memory[46082] <=  8'h00;      memory[46083] <=  8'h00;      memory[46084] <=  8'h00;      memory[46085] <=  8'h00;      memory[46086] <=  8'h00;      memory[46087] <=  8'h00;      memory[46088] <=  8'h00;      memory[46089] <=  8'h00;      memory[46090] <=  8'h00;      memory[46091] <=  8'h00;      memory[46092] <=  8'h00;      memory[46093] <=  8'h00;      memory[46094] <=  8'h00;      memory[46095] <=  8'h00;      memory[46096] <=  8'h00;      memory[46097] <=  8'h00;      memory[46098] <=  8'h00;      memory[46099] <=  8'h00;      memory[46100] <=  8'h00;      memory[46101] <=  8'h00;      memory[46102] <=  8'h00;      memory[46103] <=  8'h00;      memory[46104] <=  8'h00;      memory[46105] <=  8'h00;      memory[46106] <=  8'h00;      memory[46107] <=  8'h00;      memory[46108] <=  8'h00;      memory[46109] <=  8'h00;      memory[46110] <=  8'h00;      memory[46111] <=  8'h00;      memory[46112] <=  8'h00;      memory[46113] <=  8'h00;      memory[46114] <=  8'h00;      memory[46115] <=  8'h00;      memory[46116] <=  8'h00;      memory[46117] <=  8'h00;      memory[46118] <=  8'h00;      memory[46119] <=  8'h00;      memory[46120] <=  8'h00;      memory[46121] <=  8'h00;      memory[46122] <=  8'h00;      memory[46123] <=  8'h00;      memory[46124] <=  8'h00;      memory[46125] <=  8'h00;      memory[46126] <=  8'h00;      memory[46127] <=  8'h00;      memory[46128] <=  8'h00;      memory[46129] <=  8'h00;      memory[46130] <=  8'h00;      memory[46131] <=  8'h00;      memory[46132] <=  8'h00;      memory[46133] <=  8'h00;      memory[46134] <=  8'h00;      memory[46135] <=  8'h00;      memory[46136] <=  8'h00;      memory[46137] <=  8'h00;      memory[46138] <=  8'h00;      memory[46139] <=  8'h00;      memory[46140] <=  8'h00;      memory[46141] <=  8'h00;      memory[46142] <=  8'h00;      memory[46143] <=  8'h00;      memory[46144] <=  8'h00;      memory[46145] <=  8'h00;      memory[46146] <=  8'h00;      memory[46147] <=  8'h00;      memory[46148] <=  8'h00;      memory[46149] <=  8'h00;      memory[46150] <=  8'h00;      memory[46151] <=  8'h00;      memory[46152] <=  8'h00;      memory[46153] <=  8'h00;      memory[46154] <=  8'h00;      memory[46155] <=  8'h00;      memory[46156] <=  8'h00;      memory[46157] <=  8'h00;      memory[46158] <=  8'h00;      memory[46159] <=  8'h00;      memory[46160] <=  8'h00;      memory[46161] <=  8'h00;      memory[46162] <=  8'h00;      memory[46163] <=  8'h00;      memory[46164] <=  8'h00;      memory[46165] <=  8'h00;      memory[46166] <=  8'h00;      memory[46167] <=  8'h00;      memory[46168] <=  8'h00;      memory[46169] <=  8'h00;      memory[46170] <=  8'h00;      memory[46171] <=  8'h00;      memory[46172] <=  8'h00;      memory[46173] <=  8'h00;      memory[46174] <=  8'h00;      memory[46175] <=  8'h00;      memory[46176] <=  8'h00;      memory[46177] <=  8'h00;      memory[46178] <=  8'h00;      memory[46179] <=  8'h00;      memory[46180] <=  8'h00;      memory[46181] <=  8'h00;      memory[46182] <=  8'h00;      memory[46183] <=  8'h00;      memory[46184] <=  8'h00;      memory[46185] <=  8'h00;      memory[46186] <=  8'h00;      memory[46187] <=  8'h00;      memory[46188] <=  8'h00;      memory[46189] <=  8'h00;      memory[46190] <=  8'h00;      memory[46191] <=  8'h00;      memory[46192] <=  8'h00;      memory[46193] <=  8'h00;      memory[46194] <=  8'h00;      memory[46195] <=  8'h00;      memory[46196] <=  8'h00;      memory[46197] <=  8'h00;      memory[46198] <=  8'h00;      memory[46199] <=  8'h00;      memory[46200] <=  8'h00;      memory[46201] <=  8'h00;      memory[46202] <=  8'h00;      memory[46203] <=  8'h00;      memory[46204] <=  8'h00;      memory[46205] <=  8'h00;      memory[46206] <=  8'h00;      memory[46207] <=  8'h00;      memory[46208] <=  8'h00;      memory[46209] <=  8'h00;      memory[46210] <=  8'h00;      memory[46211] <=  8'h00;      memory[46212] <=  8'h00;      memory[46213] <=  8'h00;      memory[46214] <=  8'h00;      memory[46215] <=  8'h00;      memory[46216] <=  8'h00;      memory[46217] <=  8'h00;      memory[46218] <=  8'h00;      memory[46219] <=  8'h00;      memory[46220] <=  8'h00;      memory[46221] <=  8'h00;      memory[46222] <=  8'h00;      memory[46223] <=  8'h00;      memory[46224] <=  8'h00;      memory[46225] <=  8'h00;      memory[46226] <=  8'h00;      memory[46227] <=  8'h00;      memory[46228] <=  8'h00;      memory[46229] <=  8'h00;      memory[46230] <=  8'h00;      memory[46231] <=  8'h00;      memory[46232] <=  8'h00;      memory[46233] <=  8'h00;      memory[46234] <=  8'h00;      memory[46235] <=  8'h00;      memory[46236] <=  8'h00;      memory[46237] <=  8'h00;      memory[46238] <=  8'h00;      memory[46239] <=  8'h00;      memory[46240] <=  8'h00;      memory[46241] <=  8'h00;      memory[46242] <=  8'h00;      memory[46243] <=  8'h00;      memory[46244] <=  8'h00;      memory[46245] <=  8'h00;      memory[46246] <=  8'h00;      memory[46247] <=  8'h00;      memory[46248] <=  8'h00;      memory[46249] <=  8'h00;      memory[46250] <=  8'h00;      memory[46251] <=  8'h00;      memory[46252] <=  8'h00;      memory[46253] <=  8'h00;      memory[46254] <=  8'h00;      memory[46255] <=  8'h00;      memory[46256] <=  8'h00;      memory[46257] <=  8'h00;      memory[46258] <=  8'h00;      memory[46259] <=  8'h00;      memory[46260] <=  8'h00;      memory[46261] <=  8'h00;      memory[46262] <=  8'h00;      memory[46263] <=  8'h00;      memory[46264] <=  8'h00;      memory[46265] <=  8'h00;      memory[46266] <=  8'h00;      memory[46267] <=  8'h00;      memory[46268] <=  8'h00;      memory[46269] <=  8'h00;      memory[46270] <=  8'h00;      memory[46271] <=  8'h00;      memory[46272] <=  8'h00;      memory[46273] <=  8'h00;      memory[46274] <=  8'h00;      memory[46275] <=  8'h00;      memory[46276] <=  8'h00;      memory[46277] <=  8'h00;      memory[46278] <=  8'h00;      memory[46279] <=  8'h00;      memory[46280] <=  8'h00;      memory[46281] <=  8'h00;      memory[46282] <=  8'h00;      memory[46283] <=  8'h00;      memory[46284] <=  8'h00;      memory[46285] <=  8'h00;      memory[46286] <=  8'h00;      memory[46287] <=  8'h00;      memory[46288] <=  8'h00;      memory[46289] <=  8'h00;      memory[46290] <=  8'h00;      memory[46291] <=  8'h00;      memory[46292] <=  8'h00;      memory[46293] <=  8'h00;      memory[46294] <=  8'h00;      memory[46295] <=  8'h00;      memory[46296] <=  8'h00;      memory[46297] <=  8'h00;      memory[46298] <=  8'h00;      memory[46299] <=  8'h00;      memory[46300] <=  8'h00;      memory[46301] <=  8'h00;      memory[46302] <=  8'h00;      memory[46303] <=  8'h00;      memory[46304] <=  8'h00;      memory[46305] <=  8'h00;      memory[46306] <=  8'h00;      memory[46307] <=  8'h00;      memory[46308] <=  8'h00;      memory[46309] <=  8'h00;      memory[46310] <=  8'h00;      memory[46311] <=  8'h00;      memory[46312] <=  8'h00;      memory[46313] <=  8'h00;      memory[46314] <=  8'h00;      memory[46315] <=  8'h00;      memory[46316] <=  8'h00;      memory[46317] <=  8'h00;      memory[46318] <=  8'h00;      memory[46319] <=  8'h00;      memory[46320] <=  8'h00;      memory[46321] <=  8'h00;      memory[46322] <=  8'h00;      memory[46323] <=  8'h00;      memory[46324] <=  8'h00;      memory[46325] <=  8'h00;      memory[46326] <=  8'h00;      memory[46327] <=  8'h00;      memory[46328] <=  8'h00;      memory[46329] <=  8'h00;      memory[46330] <=  8'h00;      memory[46331] <=  8'h00;      memory[46332] <=  8'h00;      memory[46333] <=  8'h00;      memory[46334] <=  8'h00;      memory[46335] <=  8'h00;      memory[46336] <=  8'h00;      memory[46337] <=  8'h00;      memory[46338] <=  8'h00;      memory[46339] <=  8'h00;      memory[46340] <=  8'h00;      memory[46341] <=  8'h00;      memory[46342] <=  8'h00;      memory[46343] <=  8'h00;      memory[46344] <=  8'h00;      memory[46345] <=  8'h00;      memory[46346] <=  8'h00;      memory[46347] <=  8'h00;      memory[46348] <=  8'h00;      memory[46349] <=  8'h00;      memory[46350] <=  8'h00;      memory[46351] <=  8'h00;      memory[46352] <=  8'h00;      memory[46353] <=  8'h00;      memory[46354] <=  8'h00;      memory[46355] <=  8'h00;      memory[46356] <=  8'h00;      memory[46357] <=  8'h00;      memory[46358] <=  8'h00;      memory[46359] <=  8'h00;      memory[46360] <=  8'h00;      memory[46361] <=  8'h00;      memory[46362] <=  8'h00;      memory[46363] <=  8'h00;      memory[46364] <=  8'h00;      memory[46365] <=  8'h00;      memory[46366] <=  8'h00;      memory[46367] <=  8'h00;      memory[46368] <=  8'h00;      memory[46369] <=  8'h00;      memory[46370] <=  8'h00;      memory[46371] <=  8'h00;      memory[46372] <=  8'h00;      memory[46373] <=  8'h00;      memory[46374] <=  8'h00;      memory[46375] <=  8'h00;      memory[46376] <=  8'h00;      memory[46377] <=  8'h00;      memory[46378] <=  8'h00;      memory[46379] <=  8'h00;      memory[46380] <=  8'h00;      memory[46381] <=  8'h00;      memory[46382] <=  8'h00;      memory[46383] <=  8'h00;      memory[46384] <=  8'h00;      memory[46385] <=  8'h00;      memory[46386] <=  8'h00;      memory[46387] <=  8'h00;      memory[46388] <=  8'h00;      memory[46389] <=  8'h00;      memory[46390] <=  8'h00;      memory[46391] <=  8'h00;      memory[46392] <=  8'h00;      memory[46393] <=  8'h00;      memory[46394] <=  8'h00;      memory[46395] <=  8'h00;      memory[46396] <=  8'h00;      memory[46397] <=  8'h00;      memory[46398] <=  8'h00;      memory[46399] <=  8'h00;      memory[46400] <=  8'h00;      memory[46401] <=  8'h00;      memory[46402] <=  8'h00;      memory[46403] <=  8'h00;      memory[46404] <=  8'h00;      memory[46405] <=  8'h00;      memory[46406] <=  8'h00;      memory[46407] <=  8'h00;      memory[46408] <=  8'h00;      memory[46409] <=  8'h00;      memory[46410] <=  8'h00;      memory[46411] <=  8'h00;      memory[46412] <=  8'h00;      memory[46413] <=  8'h00;      memory[46414] <=  8'h00;      memory[46415] <=  8'h00;      memory[46416] <=  8'h00;      memory[46417] <=  8'h00;      memory[46418] <=  8'h00;      memory[46419] <=  8'h00;      memory[46420] <=  8'h00;      memory[46421] <=  8'h00;      memory[46422] <=  8'h00;      memory[46423] <=  8'h00;      memory[46424] <=  8'h00;      memory[46425] <=  8'h00;      memory[46426] <=  8'h00;      memory[46427] <=  8'h00;      memory[46428] <=  8'h00;      memory[46429] <=  8'h00;      memory[46430] <=  8'h00;      memory[46431] <=  8'h00;      memory[46432] <=  8'h00;      memory[46433] <=  8'h00;      memory[46434] <=  8'h00;      memory[46435] <=  8'h00;      memory[46436] <=  8'h00;      memory[46437] <=  8'h00;      memory[46438] <=  8'h00;      memory[46439] <=  8'h00;      memory[46440] <=  8'h00;      memory[46441] <=  8'h00;      memory[46442] <=  8'h00;      memory[46443] <=  8'h00;      memory[46444] <=  8'h00;      memory[46445] <=  8'h00;      memory[46446] <=  8'h00;      memory[46447] <=  8'h00;      memory[46448] <=  8'h00;      memory[46449] <=  8'h00;      memory[46450] <=  8'h00;      memory[46451] <=  8'h00;      memory[46452] <=  8'h00;      memory[46453] <=  8'h00;      memory[46454] <=  8'h00;      memory[46455] <=  8'h00;      memory[46456] <=  8'h00;      memory[46457] <=  8'h00;      memory[46458] <=  8'h00;      memory[46459] <=  8'h00;      memory[46460] <=  8'h00;      memory[46461] <=  8'h00;      memory[46462] <=  8'h00;      memory[46463] <=  8'h00;      memory[46464] <=  8'h00;      memory[46465] <=  8'h00;      memory[46466] <=  8'h00;      memory[46467] <=  8'h00;      memory[46468] <=  8'h00;      memory[46469] <=  8'h00;      memory[46470] <=  8'h00;      memory[46471] <=  8'h00;      memory[46472] <=  8'h00;      memory[46473] <=  8'h00;      memory[46474] <=  8'h00;      memory[46475] <=  8'h00;      memory[46476] <=  8'h00;      memory[46477] <=  8'h00;      memory[46478] <=  8'h00;      memory[46479] <=  8'h00;      memory[46480] <=  8'h00;      memory[46481] <=  8'h00;      memory[46482] <=  8'h00;      memory[46483] <=  8'h00;      memory[46484] <=  8'h00;      memory[46485] <=  8'h00;      memory[46486] <=  8'h00;      memory[46487] <=  8'h00;      memory[46488] <=  8'h00;      memory[46489] <=  8'h00;      memory[46490] <=  8'h00;      memory[46491] <=  8'h00;      memory[46492] <=  8'h00;      memory[46493] <=  8'h00;      memory[46494] <=  8'h00;      memory[46495] <=  8'h00;      memory[46496] <=  8'h00;      memory[46497] <=  8'h00;      memory[46498] <=  8'h00;      memory[46499] <=  8'h00;      memory[46500] <=  8'h00;      memory[46501] <=  8'h00;      memory[46502] <=  8'h00;      memory[46503] <=  8'h00;      memory[46504] <=  8'h00;      memory[46505] <=  8'h00;      memory[46506] <=  8'h00;      memory[46507] <=  8'h00;      memory[46508] <=  8'h00;      memory[46509] <=  8'h00;      memory[46510] <=  8'h00;      memory[46511] <=  8'h00;      memory[46512] <=  8'h00;      memory[46513] <=  8'h00;      memory[46514] <=  8'h00;      memory[46515] <=  8'h00;      memory[46516] <=  8'h00;      memory[46517] <=  8'h00;      memory[46518] <=  8'h00;      memory[46519] <=  8'h00;      memory[46520] <=  8'h00;      memory[46521] <=  8'h00;      memory[46522] <=  8'h00;      memory[46523] <=  8'h00;      memory[46524] <=  8'h00;      memory[46525] <=  8'h00;      memory[46526] <=  8'h00;      memory[46527] <=  8'h00;      memory[46528] <=  8'h00;      memory[46529] <=  8'h00;      memory[46530] <=  8'h00;      memory[46531] <=  8'h00;      memory[46532] <=  8'h00;      memory[46533] <=  8'h00;      memory[46534] <=  8'h00;      memory[46535] <=  8'h00;      memory[46536] <=  8'h00;      memory[46537] <=  8'h00;      memory[46538] <=  8'h00;      memory[46539] <=  8'h00;      memory[46540] <=  8'h00;      memory[46541] <=  8'h00;      memory[46542] <=  8'h00;      memory[46543] <=  8'h00;      memory[46544] <=  8'h00;      memory[46545] <=  8'h00;      memory[46546] <=  8'h00;      memory[46547] <=  8'h00;      memory[46548] <=  8'h00;      memory[46549] <=  8'h00;      memory[46550] <=  8'h00;      memory[46551] <=  8'h00;      memory[46552] <=  8'h00;      memory[46553] <=  8'h00;      memory[46554] <=  8'h00;      memory[46555] <=  8'h00;      memory[46556] <=  8'h00;      memory[46557] <=  8'h00;      memory[46558] <=  8'h00;      memory[46559] <=  8'h00;      memory[46560] <=  8'h00;      memory[46561] <=  8'h00;      memory[46562] <=  8'h00;      memory[46563] <=  8'h00;      memory[46564] <=  8'h00;      memory[46565] <=  8'h00;      memory[46566] <=  8'h00;      memory[46567] <=  8'h00;      memory[46568] <=  8'h00;      memory[46569] <=  8'h00;      memory[46570] <=  8'h00;      memory[46571] <=  8'h00;      memory[46572] <=  8'h00;      memory[46573] <=  8'h00;      memory[46574] <=  8'h00;      memory[46575] <=  8'h00;      memory[46576] <=  8'h00;      memory[46577] <=  8'h00;      memory[46578] <=  8'h00;      memory[46579] <=  8'h00;      memory[46580] <=  8'h00;      memory[46581] <=  8'h00;      memory[46582] <=  8'h00;      memory[46583] <=  8'h00;      memory[46584] <=  8'h00;      memory[46585] <=  8'h00;      memory[46586] <=  8'h00;      memory[46587] <=  8'h00;      memory[46588] <=  8'h00;      memory[46589] <=  8'h00;      memory[46590] <=  8'h00;      memory[46591] <=  8'h00;      memory[46592] <=  8'h00;      memory[46593] <=  8'h00;      memory[46594] <=  8'h00;      memory[46595] <=  8'h00;      memory[46596] <=  8'h00;      memory[46597] <=  8'h00;      memory[46598] <=  8'h00;      memory[46599] <=  8'h00;      memory[46600] <=  8'h00;      memory[46601] <=  8'h00;      memory[46602] <=  8'h00;      memory[46603] <=  8'h00;      memory[46604] <=  8'h00;      memory[46605] <=  8'h00;      memory[46606] <=  8'h00;      memory[46607] <=  8'h00;      memory[46608] <=  8'h00;      memory[46609] <=  8'h00;      memory[46610] <=  8'h00;      memory[46611] <=  8'h00;      memory[46612] <=  8'h00;      memory[46613] <=  8'h00;      memory[46614] <=  8'h00;      memory[46615] <=  8'h00;      memory[46616] <=  8'h00;      memory[46617] <=  8'h00;      memory[46618] <=  8'h00;      memory[46619] <=  8'h00;      memory[46620] <=  8'h00;      memory[46621] <=  8'h00;      memory[46622] <=  8'h00;      memory[46623] <=  8'h00;      memory[46624] <=  8'h00;      memory[46625] <=  8'h00;      memory[46626] <=  8'h00;      memory[46627] <=  8'h00;      memory[46628] <=  8'h00;      memory[46629] <=  8'h00;      memory[46630] <=  8'h00;      memory[46631] <=  8'h00;      memory[46632] <=  8'h00;      memory[46633] <=  8'h00;      memory[46634] <=  8'h00;      memory[46635] <=  8'h00;      memory[46636] <=  8'h00;      memory[46637] <=  8'h00;      memory[46638] <=  8'h00;      memory[46639] <=  8'h00;      memory[46640] <=  8'h00;      memory[46641] <=  8'h00;      memory[46642] <=  8'h00;      memory[46643] <=  8'h00;      memory[46644] <=  8'h00;      memory[46645] <=  8'h00;      memory[46646] <=  8'h00;      memory[46647] <=  8'h00;      memory[46648] <=  8'h00;      memory[46649] <=  8'h00;      memory[46650] <=  8'h00;      memory[46651] <=  8'h00;      memory[46652] <=  8'h00;      memory[46653] <=  8'h00;      memory[46654] <=  8'h00;      memory[46655] <=  8'h00;      memory[46656] <=  8'h00;      memory[46657] <=  8'h00;      memory[46658] <=  8'h00;      memory[46659] <=  8'h00;      memory[46660] <=  8'h00;      memory[46661] <=  8'h00;      memory[46662] <=  8'h00;      memory[46663] <=  8'h00;      memory[46664] <=  8'h00;      memory[46665] <=  8'h00;      memory[46666] <=  8'h00;      memory[46667] <=  8'h00;      memory[46668] <=  8'h00;      memory[46669] <=  8'h00;      memory[46670] <=  8'h00;      memory[46671] <=  8'h00;      memory[46672] <=  8'h00;      memory[46673] <=  8'h00;      memory[46674] <=  8'h00;      memory[46675] <=  8'h00;      memory[46676] <=  8'h00;      memory[46677] <=  8'h00;      memory[46678] <=  8'h00;      memory[46679] <=  8'h00;      memory[46680] <=  8'h00;      memory[46681] <=  8'h00;      memory[46682] <=  8'h00;      memory[46683] <=  8'h00;      memory[46684] <=  8'h00;      memory[46685] <=  8'h00;      memory[46686] <=  8'h00;      memory[46687] <=  8'h00;      memory[46688] <=  8'h00;      memory[46689] <=  8'h00;      memory[46690] <=  8'h00;      memory[46691] <=  8'h00;      memory[46692] <=  8'h00;      memory[46693] <=  8'h00;      memory[46694] <=  8'h00;      memory[46695] <=  8'h00;      memory[46696] <=  8'h00;      memory[46697] <=  8'h00;      memory[46698] <=  8'h00;      memory[46699] <=  8'h00;      memory[46700] <=  8'h00;      memory[46701] <=  8'h00;      memory[46702] <=  8'h00;      memory[46703] <=  8'h00;      memory[46704] <=  8'h00;      memory[46705] <=  8'h00;      memory[46706] <=  8'h00;      memory[46707] <=  8'h00;      memory[46708] <=  8'h00;      memory[46709] <=  8'h00;      memory[46710] <=  8'h00;      memory[46711] <=  8'h00;      memory[46712] <=  8'h00;      memory[46713] <=  8'h00;      memory[46714] <=  8'h00;      memory[46715] <=  8'h00;      memory[46716] <=  8'h00;      memory[46717] <=  8'h00;      memory[46718] <=  8'h00;      memory[46719] <=  8'h00;      memory[46720] <=  8'h00;      memory[46721] <=  8'h00;      memory[46722] <=  8'h00;      memory[46723] <=  8'h00;      memory[46724] <=  8'h00;      memory[46725] <=  8'h00;      memory[46726] <=  8'h00;      memory[46727] <=  8'h00;      memory[46728] <=  8'h00;      memory[46729] <=  8'h00;      memory[46730] <=  8'h00;      memory[46731] <=  8'h00;      memory[46732] <=  8'h00;      memory[46733] <=  8'h00;      memory[46734] <=  8'h00;      memory[46735] <=  8'h00;      memory[46736] <=  8'h00;      memory[46737] <=  8'h00;      memory[46738] <=  8'h00;      memory[46739] <=  8'h00;      memory[46740] <=  8'h00;      memory[46741] <=  8'h00;      memory[46742] <=  8'h00;      memory[46743] <=  8'h00;      memory[46744] <=  8'h00;      memory[46745] <=  8'h00;      memory[46746] <=  8'h00;      memory[46747] <=  8'h00;      memory[46748] <=  8'h00;      memory[46749] <=  8'h00;      memory[46750] <=  8'h00;      memory[46751] <=  8'h00;      memory[46752] <=  8'h00;      memory[46753] <=  8'h00;      memory[46754] <=  8'h00;      memory[46755] <=  8'h00;      memory[46756] <=  8'h00;      memory[46757] <=  8'h00;      memory[46758] <=  8'h00;      memory[46759] <=  8'h00;      memory[46760] <=  8'h00;      memory[46761] <=  8'h00;      memory[46762] <=  8'h00;      memory[46763] <=  8'h00;      memory[46764] <=  8'h00;      memory[46765] <=  8'h00;      memory[46766] <=  8'h00;      memory[46767] <=  8'h00;      memory[46768] <=  8'h00;      memory[46769] <=  8'h00;      memory[46770] <=  8'h00;      memory[46771] <=  8'h00;      memory[46772] <=  8'h00;      memory[46773] <=  8'h00;      memory[46774] <=  8'h00;      memory[46775] <=  8'h00;      memory[46776] <=  8'h00;      memory[46777] <=  8'h00;      memory[46778] <=  8'h00;      memory[46779] <=  8'h00;      memory[46780] <=  8'h00;      memory[46781] <=  8'h00;      memory[46782] <=  8'h00;      memory[46783] <=  8'h00;      memory[46784] <=  8'h00;      memory[46785] <=  8'h00;      memory[46786] <=  8'h00;      memory[46787] <=  8'h00;      memory[46788] <=  8'h00;      memory[46789] <=  8'h00;      memory[46790] <=  8'h00;      memory[46791] <=  8'h00;      memory[46792] <=  8'h00;      memory[46793] <=  8'h00;      memory[46794] <=  8'h00;      memory[46795] <=  8'h00;      memory[46796] <=  8'h00;      memory[46797] <=  8'h00;      memory[46798] <=  8'h00;      memory[46799] <=  8'h00;      memory[46800] <=  8'h00;      memory[46801] <=  8'h00;      memory[46802] <=  8'h00;      memory[46803] <=  8'h00;      memory[46804] <=  8'h00;      memory[46805] <=  8'h00;      memory[46806] <=  8'h00;      memory[46807] <=  8'h00;      memory[46808] <=  8'h00;      memory[46809] <=  8'h00;      memory[46810] <=  8'h00;      memory[46811] <=  8'h00;      memory[46812] <=  8'h00;      memory[46813] <=  8'h00;      memory[46814] <=  8'h00;      memory[46815] <=  8'h00;      memory[46816] <=  8'h00;      memory[46817] <=  8'h00;      memory[46818] <=  8'h00;      memory[46819] <=  8'h00;      memory[46820] <=  8'h00;      memory[46821] <=  8'h00;      memory[46822] <=  8'h00;      memory[46823] <=  8'h00;      memory[46824] <=  8'h00;      memory[46825] <=  8'h00;      memory[46826] <=  8'h00;      memory[46827] <=  8'h00;      memory[46828] <=  8'h00;      memory[46829] <=  8'h00;      memory[46830] <=  8'h00;      memory[46831] <=  8'h00;      memory[46832] <=  8'h00;      memory[46833] <=  8'h00;      memory[46834] <=  8'h00;      memory[46835] <=  8'h00;      memory[46836] <=  8'h00;      memory[46837] <=  8'h00;      memory[46838] <=  8'h00;      memory[46839] <=  8'h00;      memory[46840] <=  8'h00;      memory[46841] <=  8'h00;      memory[46842] <=  8'h00;      memory[46843] <=  8'h00;      memory[46844] <=  8'h00;      memory[46845] <=  8'h00;      memory[46846] <=  8'h00;      memory[46847] <=  8'h00;      memory[46848] <=  8'h00;      memory[46849] <=  8'h00;      memory[46850] <=  8'h00;      memory[46851] <=  8'h00;      memory[46852] <=  8'h00;      memory[46853] <=  8'h00;      memory[46854] <=  8'h00;      memory[46855] <=  8'h00;      memory[46856] <=  8'h00;      memory[46857] <=  8'h00;      memory[46858] <=  8'h00;      memory[46859] <=  8'h00;      memory[46860] <=  8'h00;      memory[46861] <=  8'h00;      memory[46862] <=  8'h00;      memory[46863] <=  8'h00;      memory[46864] <=  8'h00;      memory[46865] <=  8'h00;      memory[46866] <=  8'h00;      memory[46867] <=  8'h00;      memory[46868] <=  8'h00;      memory[46869] <=  8'h00;      memory[46870] <=  8'h00;      memory[46871] <=  8'h00;      memory[46872] <=  8'h00;      memory[46873] <=  8'h00;      memory[46874] <=  8'h00;      memory[46875] <=  8'h00;      memory[46876] <=  8'h00;      memory[46877] <=  8'h00;      memory[46878] <=  8'h00;      memory[46879] <=  8'h00;      memory[46880] <=  8'h00;      memory[46881] <=  8'h00;      memory[46882] <=  8'h00;      memory[46883] <=  8'h00;      memory[46884] <=  8'h00;      memory[46885] <=  8'h00;      memory[46886] <=  8'h00;      memory[46887] <=  8'h00;      memory[46888] <=  8'h00;      memory[46889] <=  8'h00;      memory[46890] <=  8'h00;      memory[46891] <=  8'h00;      memory[46892] <=  8'h00;      memory[46893] <=  8'h00;      memory[46894] <=  8'h00;      memory[46895] <=  8'h00;      memory[46896] <=  8'h00;      memory[46897] <=  8'h00;      memory[46898] <=  8'h00;      memory[46899] <=  8'h00;      memory[46900] <=  8'h00;      memory[46901] <=  8'h00;      memory[46902] <=  8'h00;      memory[46903] <=  8'h00;      memory[46904] <=  8'h00;      memory[46905] <=  8'h00;      memory[46906] <=  8'h00;      memory[46907] <=  8'h00;      memory[46908] <=  8'h00;      memory[46909] <=  8'h00;      memory[46910] <=  8'h00;      memory[46911] <=  8'h00;      memory[46912] <=  8'h00;      memory[46913] <=  8'h00;      memory[46914] <=  8'h00;      memory[46915] <=  8'h00;      memory[46916] <=  8'h00;      memory[46917] <=  8'h00;      memory[46918] <=  8'h00;      memory[46919] <=  8'h00;      memory[46920] <=  8'h00;      memory[46921] <=  8'h00;      memory[46922] <=  8'h00;      memory[46923] <=  8'h00;      memory[46924] <=  8'h00;      memory[46925] <=  8'h00;      memory[46926] <=  8'h00;      memory[46927] <=  8'h00;      memory[46928] <=  8'h00;      memory[46929] <=  8'h00;      memory[46930] <=  8'h00;      memory[46931] <=  8'h00;      memory[46932] <=  8'h00;      memory[46933] <=  8'h00;      memory[46934] <=  8'h00;      memory[46935] <=  8'h00;      memory[46936] <=  8'h00;      memory[46937] <=  8'h00;      memory[46938] <=  8'h00;      memory[46939] <=  8'h00;      memory[46940] <=  8'h00;      memory[46941] <=  8'h00;      memory[46942] <=  8'h00;      memory[46943] <=  8'h00;      memory[46944] <=  8'h00;      memory[46945] <=  8'h00;      memory[46946] <=  8'h00;      memory[46947] <=  8'h00;      memory[46948] <=  8'h00;      memory[46949] <=  8'h00;      memory[46950] <=  8'h00;      memory[46951] <=  8'h00;      memory[46952] <=  8'h00;      memory[46953] <=  8'h00;      memory[46954] <=  8'h00;      memory[46955] <=  8'h00;      memory[46956] <=  8'h00;      memory[46957] <=  8'h00;      memory[46958] <=  8'h00;      memory[46959] <=  8'h00;      memory[46960] <=  8'h00;      memory[46961] <=  8'h00;      memory[46962] <=  8'h00;      memory[46963] <=  8'h00;      memory[46964] <=  8'h00;      memory[46965] <=  8'h00;      memory[46966] <=  8'h00;      memory[46967] <=  8'h00;      memory[46968] <=  8'h00;      memory[46969] <=  8'h00;      memory[46970] <=  8'h00;      memory[46971] <=  8'h00;      memory[46972] <=  8'h00;      memory[46973] <=  8'h00;      memory[46974] <=  8'h00;      memory[46975] <=  8'h00;      memory[46976] <=  8'h00;      memory[46977] <=  8'h00;      memory[46978] <=  8'h00;      memory[46979] <=  8'h00;      memory[46980] <=  8'h00;      memory[46981] <=  8'h00;      memory[46982] <=  8'h00;      memory[46983] <=  8'h00;      memory[46984] <=  8'h00;      memory[46985] <=  8'h00;      memory[46986] <=  8'h00;      memory[46987] <=  8'h00;      memory[46988] <=  8'h00;      memory[46989] <=  8'h00;      memory[46990] <=  8'h00;      memory[46991] <=  8'h00;      memory[46992] <=  8'h00;      memory[46993] <=  8'h00;      memory[46994] <=  8'h00;      memory[46995] <=  8'h00;      memory[46996] <=  8'h00;      memory[46997] <=  8'h00;      memory[46998] <=  8'h00;      memory[46999] <=  8'h00;      memory[47000] <=  8'h00;      memory[47001] <=  8'h00;      memory[47002] <=  8'h00;      memory[47003] <=  8'h00;      memory[47004] <=  8'h00;      memory[47005] <=  8'h00;      memory[47006] <=  8'h00;      memory[47007] <=  8'h00;      memory[47008] <=  8'h00;      memory[47009] <=  8'h00;      memory[47010] <=  8'h00;      memory[47011] <=  8'h00;      memory[47012] <=  8'h00;      memory[47013] <=  8'h00;      memory[47014] <=  8'h00;      memory[47015] <=  8'h00;      memory[47016] <=  8'h00;      memory[47017] <=  8'h00;      memory[47018] <=  8'h00;      memory[47019] <=  8'h00;      memory[47020] <=  8'h00;      memory[47021] <=  8'h00;      memory[47022] <=  8'h00;      memory[47023] <=  8'h00;      memory[47024] <=  8'h00;      memory[47025] <=  8'h00;      memory[47026] <=  8'h00;      memory[47027] <=  8'h00;      memory[47028] <=  8'h00;      memory[47029] <=  8'h00;      memory[47030] <=  8'h00;      memory[47031] <=  8'h00;      memory[47032] <=  8'h00;      memory[47033] <=  8'h00;      memory[47034] <=  8'h00;      memory[47035] <=  8'h00;      memory[47036] <=  8'h00;      memory[47037] <=  8'h00;      memory[47038] <=  8'h00;      memory[47039] <=  8'h00;      memory[47040] <=  8'h00;      memory[47041] <=  8'h00;      memory[47042] <=  8'h00;      memory[47043] <=  8'h00;      memory[47044] <=  8'h00;      memory[47045] <=  8'h00;      memory[47046] <=  8'h00;      memory[47047] <=  8'h00;      memory[47048] <=  8'h00;      memory[47049] <=  8'h00;      memory[47050] <=  8'h00;      memory[47051] <=  8'h00;      memory[47052] <=  8'h00;      memory[47053] <=  8'h00;      memory[47054] <=  8'h00;      memory[47055] <=  8'h00;      memory[47056] <=  8'h00;      memory[47057] <=  8'h00;      memory[47058] <=  8'h00;      memory[47059] <=  8'h00;      memory[47060] <=  8'h00;      memory[47061] <=  8'h00;      memory[47062] <=  8'h00;      memory[47063] <=  8'h00;      memory[47064] <=  8'h00;      memory[47065] <=  8'h00;      memory[47066] <=  8'h00;      memory[47067] <=  8'h00;      memory[47068] <=  8'h00;      memory[47069] <=  8'h00;      memory[47070] <=  8'h00;      memory[47071] <=  8'h00;      memory[47072] <=  8'h00;      memory[47073] <=  8'h00;      memory[47074] <=  8'h00;      memory[47075] <=  8'h00;      memory[47076] <=  8'h00;      memory[47077] <=  8'h00;      memory[47078] <=  8'h00;      memory[47079] <=  8'h00;      memory[47080] <=  8'h00;      memory[47081] <=  8'h00;      memory[47082] <=  8'h00;      memory[47083] <=  8'h00;      memory[47084] <=  8'h00;      memory[47085] <=  8'h00;      memory[47086] <=  8'h00;      memory[47087] <=  8'h00;      memory[47088] <=  8'h00;      memory[47089] <=  8'h00;      memory[47090] <=  8'h00;      memory[47091] <=  8'h00;      memory[47092] <=  8'h00;      memory[47093] <=  8'h00;      memory[47094] <=  8'h00;      memory[47095] <=  8'h00;      memory[47096] <=  8'h00;      memory[47097] <=  8'h00;      memory[47098] <=  8'h00;      memory[47099] <=  8'h00;      memory[47100] <=  8'h00;      memory[47101] <=  8'h00;      memory[47102] <=  8'h00;      memory[47103] <=  8'h00;      memory[47104] <=  8'h00;      memory[47105] <=  8'h00;      memory[47106] <=  8'h00;      memory[47107] <=  8'h00;      memory[47108] <=  8'h00;      memory[47109] <=  8'h00;      memory[47110] <=  8'h00;      memory[47111] <=  8'h00;      memory[47112] <=  8'h00;      memory[47113] <=  8'h00;      memory[47114] <=  8'h00;      memory[47115] <=  8'h00;      memory[47116] <=  8'h00;      memory[47117] <=  8'h00;      memory[47118] <=  8'h00;      memory[47119] <=  8'h00;      memory[47120] <=  8'h00;      memory[47121] <=  8'h00;      memory[47122] <=  8'h00;      memory[47123] <=  8'h00;      memory[47124] <=  8'h00;      memory[47125] <=  8'h00;      memory[47126] <=  8'h00;      memory[47127] <=  8'h00;      memory[47128] <=  8'h00;      memory[47129] <=  8'h00;      memory[47130] <=  8'h00;      memory[47131] <=  8'h00;      memory[47132] <=  8'h00;      memory[47133] <=  8'h00;      memory[47134] <=  8'h00;      memory[47135] <=  8'h00;      memory[47136] <=  8'h00;      memory[47137] <=  8'h00;      memory[47138] <=  8'h00;      memory[47139] <=  8'h00;      memory[47140] <=  8'h00;      memory[47141] <=  8'h00;      memory[47142] <=  8'h00;      memory[47143] <=  8'h00;      memory[47144] <=  8'h00;      memory[47145] <=  8'h00;      memory[47146] <=  8'h00;      memory[47147] <=  8'h00;      memory[47148] <=  8'h00;      memory[47149] <=  8'h00;      memory[47150] <=  8'h00;      memory[47151] <=  8'h00;      memory[47152] <=  8'h00;      memory[47153] <=  8'h00;      memory[47154] <=  8'h00;      memory[47155] <=  8'h00;      memory[47156] <=  8'h00;      memory[47157] <=  8'h00;      memory[47158] <=  8'h00;      memory[47159] <=  8'h00;      memory[47160] <=  8'h00;      memory[47161] <=  8'h00;      memory[47162] <=  8'h00;      memory[47163] <=  8'h00;      memory[47164] <=  8'h00;      memory[47165] <=  8'h00;      memory[47166] <=  8'h00;      memory[47167] <=  8'h00;      memory[47168] <=  8'h00;      memory[47169] <=  8'h00;      memory[47170] <=  8'h00;      memory[47171] <=  8'h00;      memory[47172] <=  8'h00;      memory[47173] <=  8'h00;      memory[47174] <=  8'h00;      memory[47175] <=  8'h00;      memory[47176] <=  8'h00;      memory[47177] <=  8'h00;      memory[47178] <=  8'h00;      memory[47179] <=  8'h00;      memory[47180] <=  8'h00;      memory[47181] <=  8'h00;      memory[47182] <=  8'h00;      memory[47183] <=  8'h00;      memory[47184] <=  8'h00;      memory[47185] <=  8'h00;      memory[47186] <=  8'h00;      memory[47187] <=  8'h00;      memory[47188] <=  8'h00;      memory[47189] <=  8'h00;      memory[47190] <=  8'h00;      memory[47191] <=  8'h00;      memory[47192] <=  8'h00;      memory[47193] <=  8'h00;      memory[47194] <=  8'h00;      memory[47195] <=  8'h00;      memory[47196] <=  8'h00;      memory[47197] <=  8'h00;      memory[47198] <=  8'h00;      memory[47199] <=  8'h00;      memory[47200] <=  8'h00;      memory[47201] <=  8'h00;      memory[47202] <=  8'h00;      memory[47203] <=  8'h00;      memory[47204] <=  8'h00;      memory[47205] <=  8'h00;      memory[47206] <=  8'h00;      memory[47207] <=  8'h00;      memory[47208] <=  8'h00;      memory[47209] <=  8'h00;      memory[47210] <=  8'h00;      memory[47211] <=  8'h00;      memory[47212] <=  8'h00;      memory[47213] <=  8'h00;      memory[47214] <=  8'h00;      memory[47215] <=  8'h00;      memory[47216] <=  8'h00;      memory[47217] <=  8'h00;      memory[47218] <=  8'h00;      memory[47219] <=  8'h00;      memory[47220] <=  8'h00;      memory[47221] <=  8'h00;      memory[47222] <=  8'h00;      memory[47223] <=  8'h00;      memory[47224] <=  8'h00;      memory[47225] <=  8'h00;      memory[47226] <=  8'h00;      memory[47227] <=  8'h00;      memory[47228] <=  8'h00;      memory[47229] <=  8'h00;      memory[47230] <=  8'h00;      memory[47231] <=  8'h00;      memory[47232] <=  8'h00;      memory[47233] <=  8'h00;      memory[47234] <=  8'h00;      memory[47235] <=  8'h00;      memory[47236] <=  8'h00;      memory[47237] <=  8'h00;      memory[47238] <=  8'h00;      memory[47239] <=  8'h00;      memory[47240] <=  8'h00;      memory[47241] <=  8'h00;      memory[47242] <=  8'h00;      memory[47243] <=  8'h00;      memory[47244] <=  8'h00;      memory[47245] <=  8'h00;      memory[47246] <=  8'h00;      memory[47247] <=  8'h00;      memory[47248] <=  8'h00;      memory[47249] <=  8'h00;      memory[47250] <=  8'h00;      memory[47251] <=  8'h00;      memory[47252] <=  8'h00;      memory[47253] <=  8'h00;      memory[47254] <=  8'h00;      memory[47255] <=  8'h00;      memory[47256] <=  8'h00;      memory[47257] <=  8'h00;      memory[47258] <=  8'h00;      memory[47259] <=  8'h00;      memory[47260] <=  8'h00;      memory[47261] <=  8'h00;      memory[47262] <=  8'h00;      memory[47263] <=  8'h00;      memory[47264] <=  8'h00;      memory[47265] <=  8'h00;      memory[47266] <=  8'h00;      memory[47267] <=  8'h00;      memory[47268] <=  8'h00;      memory[47269] <=  8'h00;      memory[47270] <=  8'h00;      memory[47271] <=  8'h00;      memory[47272] <=  8'h00;      memory[47273] <=  8'h00;      memory[47274] <=  8'h00;      memory[47275] <=  8'h00;      memory[47276] <=  8'h00;      memory[47277] <=  8'h00;      memory[47278] <=  8'h00;      memory[47279] <=  8'h00;      memory[47280] <=  8'h00;      memory[47281] <=  8'h00;      memory[47282] <=  8'h00;      memory[47283] <=  8'h00;      memory[47284] <=  8'h00;      memory[47285] <=  8'h00;      memory[47286] <=  8'h00;      memory[47287] <=  8'h00;      memory[47288] <=  8'h00;      memory[47289] <=  8'h00;      memory[47290] <=  8'h00;      memory[47291] <=  8'h00;      memory[47292] <=  8'h00;      memory[47293] <=  8'h00;      memory[47294] <=  8'h00;      memory[47295] <=  8'h00;      memory[47296] <=  8'h00;      memory[47297] <=  8'h00;      memory[47298] <=  8'h00;      memory[47299] <=  8'h00;      memory[47300] <=  8'h00;      memory[47301] <=  8'h00;      memory[47302] <=  8'h00;      memory[47303] <=  8'h00;      memory[47304] <=  8'h00;      memory[47305] <=  8'h00;      memory[47306] <=  8'h00;      memory[47307] <=  8'h00;      memory[47308] <=  8'h00;      memory[47309] <=  8'h00;      memory[47310] <=  8'h00;      memory[47311] <=  8'h00;      memory[47312] <=  8'h00;      memory[47313] <=  8'h00;      memory[47314] <=  8'h00;      memory[47315] <=  8'h00;      memory[47316] <=  8'h00;      memory[47317] <=  8'h00;      memory[47318] <=  8'h00;      memory[47319] <=  8'h00;      memory[47320] <=  8'h00;      memory[47321] <=  8'h00;      memory[47322] <=  8'h00;      memory[47323] <=  8'h00;      memory[47324] <=  8'h00;      memory[47325] <=  8'h00;      memory[47326] <=  8'h00;      memory[47327] <=  8'h00;      memory[47328] <=  8'h00;      memory[47329] <=  8'h00;      memory[47330] <=  8'h00;      memory[47331] <=  8'h00;      memory[47332] <=  8'h00;      memory[47333] <=  8'h00;      memory[47334] <=  8'h00;      memory[47335] <=  8'h00;      memory[47336] <=  8'h00;      memory[47337] <=  8'h00;      memory[47338] <=  8'h00;      memory[47339] <=  8'h00;      memory[47340] <=  8'h00;      memory[47341] <=  8'h00;      memory[47342] <=  8'h00;      memory[47343] <=  8'h00;      memory[47344] <=  8'h00;      memory[47345] <=  8'h00;      memory[47346] <=  8'h00;      memory[47347] <=  8'h00;      memory[47348] <=  8'h00;      memory[47349] <=  8'h00;      memory[47350] <=  8'h00;      memory[47351] <=  8'h00;      memory[47352] <=  8'h00;      memory[47353] <=  8'h00;      memory[47354] <=  8'h00;      memory[47355] <=  8'h00;      memory[47356] <=  8'h00;      memory[47357] <=  8'h00;      memory[47358] <=  8'h00;      memory[47359] <=  8'h00;      memory[47360] <=  8'h00;      memory[47361] <=  8'h00;      memory[47362] <=  8'h00;      memory[47363] <=  8'h00;      memory[47364] <=  8'h00;      memory[47365] <=  8'h00;      memory[47366] <=  8'h00;      memory[47367] <=  8'h00;      memory[47368] <=  8'h00;      memory[47369] <=  8'h00;      memory[47370] <=  8'h00;      memory[47371] <=  8'h00;      memory[47372] <=  8'h00;      memory[47373] <=  8'h00;      memory[47374] <=  8'h00;      memory[47375] <=  8'h00;      memory[47376] <=  8'h00;      memory[47377] <=  8'h00;      memory[47378] <=  8'h00;      memory[47379] <=  8'h00;      memory[47380] <=  8'h00;      memory[47381] <=  8'h00;      memory[47382] <=  8'h00;      memory[47383] <=  8'h00;      memory[47384] <=  8'h00;      memory[47385] <=  8'h00;      memory[47386] <=  8'h00;      memory[47387] <=  8'h00;      memory[47388] <=  8'h00;      memory[47389] <=  8'h00;      memory[47390] <=  8'h00;      memory[47391] <=  8'h00;      memory[47392] <=  8'h00;      memory[47393] <=  8'h00;      memory[47394] <=  8'h00;      memory[47395] <=  8'h00;      memory[47396] <=  8'h00;      memory[47397] <=  8'h00;      memory[47398] <=  8'h00;      memory[47399] <=  8'h00;      memory[47400] <=  8'h00;      memory[47401] <=  8'h00;      memory[47402] <=  8'h00;      memory[47403] <=  8'h00;      memory[47404] <=  8'h00;      memory[47405] <=  8'h00;      memory[47406] <=  8'h00;      memory[47407] <=  8'h00;      memory[47408] <=  8'h00;      memory[47409] <=  8'h00;      memory[47410] <=  8'h00;      memory[47411] <=  8'h00;      memory[47412] <=  8'h00;      memory[47413] <=  8'h00;      memory[47414] <=  8'h00;      memory[47415] <=  8'h00;      memory[47416] <=  8'h00;      memory[47417] <=  8'h00;      memory[47418] <=  8'h00;      memory[47419] <=  8'h00;      memory[47420] <=  8'h00;      memory[47421] <=  8'h00;      memory[47422] <=  8'h00;      memory[47423] <=  8'h00;      memory[47424] <=  8'h00;      memory[47425] <=  8'h00;      memory[47426] <=  8'h00;      memory[47427] <=  8'h00;      memory[47428] <=  8'h00;      memory[47429] <=  8'h00;      memory[47430] <=  8'h00;      memory[47431] <=  8'h00;      memory[47432] <=  8'h00;      memory[47433] <=  8'h00;      memory[47434] <=  8'h00;      memory[47435] <=  8'h00;      memory[47436] <=  8'h00;      memory[47437] <=  8'h00;      memory[47438] <=  8'h00;      memory[47439] <=  8'h00;      memory[47440] <=  8'h00;      memory[47441] <=  8'h00;      memory[47442] <=  8'h00;      memory[47443] <=  8'h00;      memory[47444] <=  8'h00;      memory[47445] <=  8'h00;      memory[47446] <=  8'h00;      memory[47447] <=  8'h00;      memory[47448] <=  8'h00;      memory[47449] <=  8'h00;      memory[47450] <=  8'h00;      memory[47451] <=  8'h00;      memory[47452] <=  8'h00;      memory[47453] <=  8'h00;      memory[47454] <=  8'h00;      memory[47455] <=  8'h00;      memory[47456] <=  8'h00;      memory[47457] <=  8'h00;      memory[47458] <=  8'h00;      memory[47459] <=  8'h00;      memory[47460] <=  8'h00;      memory[47461] <=  8'h00;      memory[47462] <=  8'h00;      memory[47463] <=  8'h00;      memory[47464] <=  8'h00;      memory[47465] <=  8'h00;      memory[47466] <=  8'h00;      memory[47467] <=  8'h00;      memory[47468] <=  8'h00;      memory[47469] <=  8'h00;      memory[47470] <=  8'h00;      memory[47471] <=  8'h00;      memory[47472] <=  8'h00;      memory[47473] <=  8'h00;      memory[47474] <=  8'h00;      memory[47475] <=  8'h00;      memory[47476] <=  8'h00;      memory[47477] <=  8'h00;      memory[47478] <=  8'h00;      memory[47479] <=  8'h00;      memory[47480] <=  8'h00;      memory[47481] <=  8'h00;      memory[47482] <=  8'h00;      memory[47483] <=  8'h00;      memory[47484] <=  8'h00;      memory[47485] <=  8'h00;      memory[47486] <=  8'h00;      memory[47487] <=  8'h00;      memory[47488] <=  8'h00;      memory[47489] <=  8'h00;      memory[47490] <=  8'h00;      memory[47491] <=  8'h00;      memory[47492] <=  8'h00;      memory[47493] <=  8'h00;      memory[47494] <=  8'h00;      memory[47495] <=  8'h00;      memory[47496] <=  8'h00;      memory[47497] <=  8'h00;      memory[47498] <=  8'h00;      memory[47499] <=  8'h00;      memory[47500] <=  8'h00;      memory[47501] <=  8'h00;      memory[47502] <=  8'h00;      memory[47503] <=  8'h00;      memory[47504] <=  8'h00;      memory[47505] <=  8'h00;      memory[47506] <=  8'h00;      memory[47507] <=  8'h00;      memory[47508] <=  8'h00;      memory[47509] <=  8'h00;      memory[47510] <=  8'h00;      memory[47511] <=  8'h00;      memory[47512] <=  8'h00;      memory[47513] <=  8'h00;      memory[47514] <=  8'h00;      memory[47515] <=  8'h00;      memory[47516] <=  8'h00;      memory[47517] <=  8'h00;      memory[47518] <=  8'h00;      memory[47519] <=  8'h00;      memory[47520] <=  8'h00;      memory[47521] <=  8'h00;      memory[47522] <=  8'h00;      memory[47523] <=  8'h00;      memory[47524] <=  8'h00;      memory[47525] <=  8'h00;      memory[47526] <=  8'h00;      memory[47527] <=  8'h00;      memory[47528] <=  8'h00;      memory[47529] <=  8'h00;      memory[47530] <=  8'h00;      memory[47531] <=  8'h00;      memory[47532] <=  8'h00;      memory[47533] <=  8'h00;      memory[47534] <=  8'h00;      memory[47535] <=  8'h00;      memory[47536] <=  8'h00;      memory[47537] <=  8'h00;      memory[47538] <=  8'h00;      memory[47539] <=  8'h00;      memory[47540] <=  8'h00;      memory[47541] <=  8'h00;      memory[47542] <=  8'h00;      memory[47543] <=  8'h00;      memory[47544] <=  8'h00;      memory[47545] <=  8'h00;      memory[47546] <=  8'h00;      memory[47547] <=  8'h00;      memory[47548] <=  8'h00;      memory[47549] <=  8'h00;      memory[47550] <=  8'h00;      memory[47551] <=  8'h00;      memory[47552] <=  8'h00;      memory[47553] <=  8'h00;      memory[47554] <=  8'h00;      memory[47555] <=  8'h00;      memory[47556] <=  8'h00;      memory[47557] <=  8'h00;      memory[47558] <=  8'h00;      memory[47559] <=  8'h00;      memory[47560] <=  8'h00;      memory[47561] <=  8'h00;      memory[47562] <=  8'h00;      memory[47563] <=  8'h00;      memory[47564] <=  8'h00;      memory[47565] <=  8'h00;      memory[47566] <=  8'h00;      memory[47567] <=  8'h00;      memory[47568] <=  8'h00;      memory[47569] <=  8'h00;      memory[47570] <=  8'h00;      memory[47571] <=  8'h00;      memory[47572] <=  8'h00;      memory[47573] <=  8'h00;      memory[47574] <=  8'h00;      memory[47575] <=  8'h00;      memory[47576] <=  8'h00;      memory[47577] <=  8'h00;      memory[47578] <=  8'h00;      memory[47579] <=  8'h00;      memory[47580] <=  8'h00;      memory[47581] <=  8'h00;      memory[47582] <=  8'h00;      memory[47583] <=  8'h00;      memory[47584] <=  8'h00;      memory[47585] <=  8'h00;      memory[47586] <=  8'h00;      memory[47587] <=  8'h00;      memory[47588] <=  8'h00;      memory[47589] <=  8'h00;      memory[47590] <=  8'h00;      memory[47591] <=  8'h00;      memory[47592] <=  8'h00;      memory[47593] <=  8'h00;      memory[47594] <=  8'h00;      memory[47595] <=  8'h00;      memory[47596] <=  8'h00;      memory[47597] <=  8'h00;      memory[47598] <=  8'h00;      memory[47599] <=  8'h00;      memory[47600] <=  8'h00;      memory[47601] <=  8'h00;      memory[47602] <=  8'h00;      memory[47603] <=  8'h00;      memory[47604] <=  8'h00;      memory[47605] <=  8'h00;      memory[47606] <=  8'h00;      memory[47607] <=  8'h00;      memory[47608] <=  8'h00;      memory[47609] <=  8'h00;      memory[47610] <=  8'h00;      memory[47611] <=  8'h00;      memory[47612] <=  8'h00;      memory[47613] <=  8'h00;      memory[47614] <=  8'h00;      memory[47615] <=  8'h00;      memory[47616] <=  8'h00;      memory[47617] <=  8'h00;      memory[47618] <=  8'h00;      memory[47619] <=  8'h00;      memory[47620] <=  8'h00;      memory[47621] <=  8'h00;      memory[47622] <=  8'h00;      memory[47623] <=  8'h00;      memory[47624] <=  8'h00;      memory[47625] <=  8'h00;      memory[47626] <=  8'h00;      memory[47627] <=  8'h00;      memory[47628] <=  8'h00;      memory[47629] <=  8'h00;      memory[47630] <=  8'h00;      memory[47631] <=  8'h00;      memory[47632] <=  8'h00;      memory[47633] <=  8'h00;      memory[47634] <=  8'h00;      memory[47635] <=  8'h00;      memory[47636] <=  8'h00;      memory[47637] <=  8'h00;      memory[47638] <=  8'h00;      memory[47639] <=  8'h00;      memory[47640] <=  8'h00;      memory[47641] <=  8'h00;      memory[47642] <=  8'h00;      memory[47643] <=  8'h00;      memory[47644] <=  8'h00;      memory[47645] <=  8'h00;      memory[47646] <=  8'h00;      memory[47647] <=  8'h00;      memory[47648] <=  8'h00;      memory[47649] <=  8'h00;      memory[47650] <=  8'h00;      memory[47651] <=  8'h00;      memory[47652] <=  8'h00;      memory[47653] <=  8'h00;      memory[47654] <=  8'h00;      memory[47655] <=  8'h00;      memory[47656] <=  8'h00;      memory[47657] <=  8'h00;      memory[47658] <=  8'h00;      memory[47659] <=  8'h00;      memory[47660] <=  8'h00;      memory[47661] <=  8'h00;      memory[47662] <=  8'h00;      memory[47663] <=  8'h00;      memory[47664] <=  8'h00;      memory[47665] <=  8'h00;      memory[47666] <=  8'h00;      memory[47667] <=  8'h00;      memory[47668] <=  8'h00;      memory[47669] <=  8'h00;      memory[47670] <=  8'h00;      memory[47671] <=  8'h00;      memory[47672] <=  8'h00;      memory[47673] <=  8'h00;      memory[47674] <=  8'h00;      memory[47675] <=  8'h00;      memory[47676] <=  8'h00;      memory[47677] <=  8'h00;      memory[47678] <=  8'h00;      memory[47679] <=  8'h00;      memory[47680] <=  8'h00;      memory[47681] <=  8'h00;      memory[47682] <=  8'h00;      memory[47683] <=  8'h00;      memory[47684] <=  8'h00;      memory[47685] <=  8'h00;      memory[47686] <=  8'h00;      memory[47687] <=  8'h00;      memory[47688] <=  8'h00;      memory[47689] <=  8'h00;      memory[47690] <=  8'h00;      memory[47691] <=  8'h00;      memory[47692] <=  8'h00;      memory[47693] <=  8'h00;      memory[47694] <=  8'h00;      memory[47695] <=  8'h00;      memory[47696] <=  8'h00;      memory[47697] <=  8'h00;      memory[47698] <=  8'h00;      memory[47699] <=  8'h00;      memory[47700] <=  8'h00;      memory[47701] <=  8'h00;      memory[47702] <=  8'h00;      memory[47703] <=  8'h00;      memory[47704] <=  8'h00;      memory[47705] <=  8'h00;      memory[47706] <=  8'h00;      memory[47707] <=  8'h00;      memory[47708] <=  8'h00;      memory[47709] <=  8'h00;      memory[47710] <=  8'h00;      memory[47711] <=  8'h00;      memory[47712] <=  8'h00;      memory[47713] <=  8'h00;      memory[47714] <=  8'h00;      memory[47715] <=  8'h00;      memory[47716] <=  8'h00;      memory[47717] <=  8'h00;      memory[47718] <=  8'h00;      memory[47719] <=  8'h00;      memory[47720] <=  8'h00;      memory[47721] <=  8'h00;      memory[47722] <=  8'h00;      memory[47723] <=  8'h00;      memory[47724] <=  8'h00;      memory[47725] <=  8'h00;      memory[47726] <=  8'h00;      memory[47727] <=  8'h00;      memory[47728] <=  8'h00;      memory[47729] <=  8'h00;      memory[47730] <=  8'h00;      memory[47731] <=  8'h00;      memory[47732] <=  8'h00;      memory[47733] <=  8'h00;      memory[47734] <=  8'h00;      memory[47735] <=  8'h00;      memory[47736] <=  8'h00;      memory[47737] <=  8'h00;      memory[47738] <=  8'h00;      memory[47739] <=  8'h00;      memory[47740] <=  8'h00;      memory[47741] <=  8'h00;      memory[47742] <=  8'h00;      memory[47743] <=  8'h00;      memory[47744] <=  8'h00;      memory[47745] <=  8'h00;      memory[47746] <=  8'h00;      memory[47747] <=  8'h00;      memory[47748] <=  8'h00;      memory[47749] <=  8'h00;      memory[47750] <=  8'h00;      memory[47751] <=  8'h00;      memory[47752] <=  8'h00;      memory[47753] <=  8'h00;      memory[47754] <=  8'h00;      memory[47755] <=  8'h00;      memory[47756] <=  8'h00;      memory[47757] <=  8'h00;      memory[47758] <=  8'h00;      memory[47759] <=  8'h00;      memory[47760] <=  8'h00;      memory[47761] <=  8'h00;      memory[47762] <=  8'h00;      memory[47763] <=  8'h00;      memory[47764] <=  8'h00;      memory[47765] <=  8'h00;      memory[47766] <=  8'h00;      memory[47767] <=  8'h00;      memory[47768] <=  8'h00;      memory[47769] <=  8'h00;      memory[47770] <=  8'h00;      memory[47771] <=  8'h00;      memory[47772] <=  8'h00;      memory[47773] <=  8'h00;      memory[47774] <=  8'h00;      memory[47775] <=  8'h00;      memory[47776] <=  8'h00;      memory[47777] <=  8'h00;      memory[47778] <=  8'h00;      memory[47779] <=  8'h00;      memory[47780] <=  8'h00;      memory[47781] <=  8'h00;      memory[47782] <=  8'h00;      memory[47783] <=  8'h00;      memory[47784] <=  8'h00;      memory[47785] <=  8'h00;      memory[47786] <=  8'h00;      memory[47787] <=  8'h00;      memory[47788] <=  8'h00;      memory[47789] <=  8'h00;      memory[47790] <=  8'h00;      memory[47791] <=  8'h00;      memory[47792] <=  8'h00;      memory[47793] <=  8'h00;      memory[47794] <=  8'h00;      memory[47795] <=  8'h00;      memory[47796] <=  8'h00;      memory[47797] <=  8'h00;      memory[47798] <=  8'h00;      memory[47799] <=  8'h00;      memory[47800] <=  8'h00;      memory[47801] <=  8'h00;      memory[47802] <=  8'h00;      memory[47803] <=  8'h00;      memory[47804] <=  8'h00;      memory[47805] <=  8'h00;      memory[47806] <=  8'h00;      memory[47807] <=  8'h00;      memory[47808] <=  8'h00;      memory[47809] <=  8'h00;      memory[47810] <=  8'h00;      memory[47811] <=  8'h00;      memory[47812] <=  8'h00;      memory[47813] <=  8'h00;      memory[47814] <=  8'h00;      memory[47815] <=  8'h00;      memory[47816] <=  8'h00;      memory[47817] <=  8'h00;      memory[47818] <=  8'h00;      memory[47819] <=  8'h00;      memory[47820] <=  8'h00;      memory[47821] <=  8'h00;      memory[47822] <=  8'h00;      memory[47823] <=  8'h00;      memory[47824] <=  8'h00;      memory[47825] <=  8'h00;      memory[47826] <=  8'h00;      memory[47827] <=  8'h00;      memory[47828] <=  8'h00;      memory[47829] <=  8'h00;      memory[47830] <=  8'h00;      memory[47831] <=  8'h00;      memory[47832] <=  8'h00;      memory[47833] <=  8'h00;      memory[47834] <=  8'h00;      memory[47835] <=  8'h00;      memory[47836] <=  8'h00;      memory[47837] <=  8'h00;      memory[47838] <=  8'h00;      memory[47839] <=  8'h00;      memory[47840] <=  8'h00;      memory[47841] <=  8'h00;      memory[47842] <=  8'h00;      memory[47843] <=  8'h00;      memory[47844] <=  8'h00;      memory[47845] <=  8'h00;      memory[47846] <=  8'h00;      memory[47847] <=  8'h00;      memory[47848] <=  8'h00;      memory[47849] <=  8'h00;      memory[47850] <=  8'h00;      memory[47851] <=  8'h00;      memory[47852] <=  8'h00;      memory[47853] <=  8'h00;      memory[47854] <=  8'h00;      memory[47855] <=  8'h00;      memory[47856] <=  8'h00;      memory[47857] <=  8'h00;      memory[47858] <=  8'h00;      memory[47859] <=  8'h00;      memory[47860] <=  8'h00;      memory[47861] <=  8'h00;      memory[47862] <=  8'h00;      memory[47863] <=  8'h00;      memory[47864] <=  8'h00;      memory[47865] <=  8'h00;      memory[47866] <=  8'h00;      memory[47867] <=  8'h00;      memory[47868] <=  8'h00;      memory[47869] <=  8'h00;      memory[47870] <=  8'h00;      memory[47871] <=  8'h00;      memory[47872] <=  8'h00;      memory[47873] <=  8'h00;      memory[47874] <=  8'h00;      memory[47875] <=  8'h00;      memory[47876] <=  8'h00;      memory[47877] <=  8'h00;      memory[47878] <=  8'h00;      memory[47879] <=  8'h00;      memory[47880] <=  8'h00;      memory[47881] <=  8'h00;      memory[47882] <=  8'h00;      memory[47883] <=  8'h00;      memory[47884] <=  8'h00;      memory[47885] <=  8'h00;      memory[47886] <=  8'h00;      memory[47887] <=  8'h00;      memory[47888] <=  8'h00;      memory[47889] <=  8'h00;      memory[47890] <=  8'h00;      memory[47891] <=  8'h00;      memory[47892] <=  8'h00;      memory[47893] <=  8'h00;      memory[47894] <=  8'h00;      memory[47895] <=  8'h00;      memory[47896] <=  8'h00;      memory[47897] <=  8'h00;      memory[47898] <=  8'h00;      memory[47899] <=  8'h00;      memory[47900] <=  8'h00;      memory[47901] <=  8'h00;      memory[47902] <=  8'h00;      memory[47903] <=  8'h00;      memory[47904] <=  8'h00;      memory[47905] <=  8'h00;      memory[47906] <=  8'h00;      memory[47907] <=  8'h00;      memory[47908] <=  8'h00;      memory[47909] <=  8'h00;      memory[47910] <=  8'h00;      memory[47911] <=  8'h00;      memory[47912] <=  8'h00;      memory[47913] <=  8'h00;      memory[47914] <=  8'h00;      memory[47915] <=  8'h00;      memory[47916] <=  8'h00;      memory[47917] <=  8'h00;      memory[47918] <=  8'h00;      memory[47919] <=  8'h00;      memory[47920] <=  8'h00;      memory[47921] <=  8'h00;      memory[47922] <=  8'h00;      memory[47923] <=  8'h00;      memory[47924] <=  8'h00;      memory[47925] <=  8'h00;      memory[47926] <=  8'h00;      memory[47927] <=  8'h00;      memory[47928] <=  8'h00;      memory[47929] <=  8'h00;      memory[47930] <=  8'h00;      memory[47931] <=  8'h00;      memory[47932] <=  8'h00;      memory[47933] <=  8'h00;      memory[47934] <=  8'h00;      memory[47935] <=  8'h00;      memory[47936] <=  8'h00;      memory[47937] <=  8'h00;      memory[47938] <=  8'h00;      memory[47939] <=  8'h00;      memory[47940] <=  8'h00;      memory[47941] <=  8'h00;      memory[47942] <=  8'h00;      memory[47943] <=  8'h00;      memory[47944] <=  8'h00;      memory[47945] <=  8'h00;      memory[47946] <=  8'h00;      memory[47947] <=  8'h00;      memory[47948] <=  8'h00;      memory[47949] <=  8'h00;      memory[47950] <=  8'h00;      memory[47951] <=  8'h00;      memory[47952] <=  8'h00;      memory[47953] <=  8'h00;      memory[47954] <=  8'h00;      memory[47955] <=  8'h00;      memory[47956] <=  8'h00;      memory[47957] <=  8'h00;      memory[47958] <=  8'h00;      memory[47959] <=  8'h00;      memory[47960] <=  8'h00;      memory[47961] <=  8'h00;      memory[47962] <=  8'h00;      memory[47963] <=  8'h00;      memory[47964] <=  8'h00;      memory[47965] <=  8'h00;      memory[47966] <=  8'h00;      memory[47967] <=  8'h00;      memory[47968] <=  8'h00;      memory[47969] <=  8'h00;      memory[47970] <=  8'h00;      memory[47971] <=  8'h00;      memory[47972] <=  8'h00;      memory[47973] <=  8'h00;      memory[47974] <=  8'h00;      memory[47975] <=  8'h00;      memory[47976] <=  8'h00;      memory[47977] <=  8'h00;      memory[47978] <=  8'h00;      memory[47979] <=  8'h00;      memory[47980] <=  8'h00;      memory[47981] <=  8'h00;      memory[47982] <=  8'h00;      memory[47983] <=  8'h00;      memory[47984] <=  8'h00;      memory[47985] <=  8'h00;      memory[47986] <=  8'h00;      memory[47987] <=  8'h00;      memory[47988] <=  8'h00;      memory[47989] <=  8'h00;      memory[47990] <=  8'h00;      memory[47991] <=  8'h00;      memory[47992] <=  8'h00;      memory[47993] <=  8'h00;      memory[47994] <=  8'h00;      memory[47995] <=  8'h00;      memory[47996] <=  8'h00;      memory[47997] <=  8'h00;      memory[47998] <=  8'h00;      memory[47999] <=  8'h00;      memory[48000] <=  8'h00;      memory[48001] <=  8'h00;      memory[48002] <=  8'h00;      memory[48003] <=  8'h00;      memory[48004] <=  8'h00;      memory[48005] <=  8'h00;      memory[48006] <=  8'h00;      memory[48007] <=  8'h00;      memory[48008] <=  8'h00;      memory[48009] <=  8'h00;      memory[48010] <=  8'h00;      memory[48011] <=  8'h00;      memory[48012] <=  8'h00;      memory[48013] <=  8'h00;      memory[48014] <=  8'h00;      memory[48015] <=  8'h00;      memory[48016] <=  8'h00;      memory[48017] <=  8'h00;      memory[48018] <=  8'h00;      memory[48019] <=  8'h00;      memory[48020] <=  8'h00;      memory[48021] <=  8'h00;      memory[48022] <=  8'h00;      memory[48023] <=  8'h00;      memory[48024] <=  8'h00;      memory[48025] <=  8'h00;      memory[48026] <=  8'h00;      memory[48027] <=  8'h00;      memory[48028] <=  8'h00;      memory[48029] <=  8'h00;      memory[48030] <=  8'h00;      memory[48031] <=  8'h00;      memory[48032] <=  8'h00;      memory[48033] <=  8'h00;      memory[48034] <=  8'h00;      memory[48035] <=  8'h00;      memory[48036] <=  8'h00;      memory[48037] <=  8'h00;      memory[48038] <=  8'h00;      memory[48039] <=  8'h00;      memory[48040] <=  8'h00;      memory[48041] <=  8'h00;      memory[48042] <=  8'h00;      memory[48043] <=  8'h00;      memory[48044] <=  8'h00;      memory[48045] <=  8'h00;      memory[48046] <=  8'h00;      memory[48047] <=  8'h00;      memory[48048] <=  8'h00;      memory[48049] <=  8'h00;      memory[48050] <=  8'h00;      memory[48051] <=  8'h00;      memory[48052] <=  8'h00;      memory[48053] <=  8'h00;      memory[48054] <=  8'h00;      memory[48055] <=  8'h00;      memory[48056] <=  8'h00;      memory[48057] <=  8'h00;      memory[48058] <=  8'h00;      memory[48059] <=  8'h00;      memory[48060] <=  8'h00;      memory[48061] <=  8'h00;      memory[48062] <=  8'h00;      memory[48063] <=  8'h00;      memory[48064] <=  8'h00;      memory[48065] <=  8'h00;      memory[48066] <=  8'h00;      memory[48067] <=  8'h00;      memory[48068] <=  8'h00;      memory[48069] <=  8'h00;      memory[48070] <=  8'h00;      memory[48071] <=  8'h00;      memory[48072] <=  8'h00;      memory[48073] <=  8'h00;      memory[48074] <=  8'h00;      memory[48075] <=  8'h00;      memory[48076] <=  8'h00;      memory[48077] <=  8'h00;      memory[48078] <=  8'h00;      memory[48079] <=  8'h00;      memory[48080] <=  8'h00;      memory[48081] <=  8'h00;      memory[48082] <=  8'h00;      memory[48083] <=  8'h00;      memory[48084] <=  8'h00;      memory[48085] <=  8'h00;      memory[48086] <=  8'h00;      memory[48087] <=  8'h00;      memory[48088] <=  8'h00;      memory[48089] <=  8'h00;      memory[48090] <=  8'h00;      memory[48091] <=  8'h00;      memory[48092] <=  8'h00;      memory[48093] <=  8'h00;      memory[48094] <=  8'h00;      memory[48095] <=  8'h00;      memory[48096] <=  8'h00;      memory[48097] <=  8'h00;      memory[48098] <=  8'h00;      memory[48099] <=  8'h00;      memory[48100] <=  8'h00;      memory[48101] <=  8'h00;      memory[48102] <=  8'h00;      memory[48103] <=  8'h00;      memory[48104] <=  8'h00;      memory[48105] <=  8'h00;      memory[48106] <=  8'h00;      memory[48107] <=  8'h00;      memory[48108] <=  8'h00;      memory[48109] <=  8'h00;      memory[48110] <=  8'h00;      memory[48111] <=  8'h00;      memory[48112] <=  8'h00;      memory[48113] <=  8'h00;      memory[48114] <=  8'h00;      memory[48115] <=  8'h00;      memory[48116] <=  8'h00;      memory[48117] <=  8'h00;      memory[48118] <=  8'h00;      memory[48119] <=  8'h00;      memory[48120] <=  8'h00;      memory[48121] <=  8'h00;      memory[48122] <=  8'h00;      memory[48123] <=  8'h00;      memory[48124] <=  8'h00;      memory[48125] <=  8'h00;      memory[48126] <=  8'h00;      memory[48127] <=  8'h00;      memory[48128] <=  8'h00;      memory[48129] <=  8'h00;      memory[48130] <=  8'h00;      memory[48131] <=  8'h00;      memory[48132] <=  8'h00;      memory[48133] <=  8'h00;      memory[48134] <=  8'h00;      memory[48135] <=  8'h00;      memory[48136] <=  8'h00;      memory[48137] <=  8'h00;      memory[48138] <=  8'h00;      memory[48139] <=  8'h00;      memory[48140] <=  8'h00;      memory[48141] <=  8'h00;      memory[48142] <=  8'h00;      memory[48143] <=  8'h00;      memory[48144] <=  8'h00;      memory[48145] <=  8'h00;      memory[48146] <=  8'h00;      memory[48147] <=  8'h00;      memory[48148] <=  8'h00;      memory[48149] <=  8'h00;      memory[48150] <=  8'h00;      memory[48151] <=  8'h00;      memory[48152] <=  8'h00;      memory[48153] <=  8'h00;      memory[48154] <=  8'h00;      memory[48155] <=  8'h00;      memory[48156] <=  8'h00;      memory[48157] <=  8'h00;      memory[48158] <=  8'h00;      memory[48159] <=  8'h00;      memory[48160] <=  8'h00;      memory[48161] <=  8'h00;      memory[48162] <=  8'h00;      memory[48163] <=  8'h00;      memory[48164] <=  8'h00;      memory[48165] <=  8'h00;      memory[48166] <=  8'h00;      memory[48167] <=  8'h00;      memory[48168] <=  8'h00;      memory[48169] <=  8'h00;      memory[48170] <=  8'h00;      memory[48171] <=  8'h00;      memory[48172] <=  8'h00;      memory[48173] <=  8'h00;      memory[48174] <=  8'h00;      memory[48175] <=  8'h00;      memory[48176] <=  8'h00;      memory[48177] <=  8'h00;      memory[48178] <=  8'h00;      memory[48179] <=  8'h00;      memory[48180] <=  8'h00;      memory[48181] <=  8'h00;      memory[48182] <=  8'h00;      memory[48183] <=  8'h00;      memory[48184] <=  8'h00;      memory[48185] <=  8'h00;      memory[48186] <=  8'h00;      memory[48187] <=  8'h00;      memory[48188] <=  8'h00;      memory[48189] <=  8'h00;      memory[48190] <=  8'h00;      memory[48191] <=  8'h00;      memory[48192] <=  8'h00;      memory[48193] <=  8'h00;      memory[48194] <=  8'h00;      memory[48195] <=  8'h00;      memory[48196] <=  8'h00;      memory[48197] <=  8'h00;      memory[48198] <=  8'h00;      memory[48199] <=  8'h00;      memory[48200] <=  8'h00;      memory[48201] <=  8'h00;      memory[48202] <=  8'h00;      memory[48203] <=  8'h00;      memory[48204] <=  8'h00;      memory[48205] <=  8'h00;      memory[48206] <=  8'h00;      memory[48207] <=  8'h00;      memory[48208] <=  8'h00;      memory[48209] <=  8'h00;      memory[48210] <=  8'h00;      memory[48211] <=  8'h00;      memory[48212] <=  8'h00;      memory[48213] <=  8'h00;      memory[48214] <=  8'h00;      memory[48215] <=  8'h00;      memory[48216] <=  8'h00;      memory[48217] <=  8'h00;      memory[48218] <=  8'h00;      memory[48219] <=  8'h00;      memory[48220] <=  8'h00;      memory[48221] <=  8'h00;      memory[48222] <=  8'h00;      memory[48223] <=  8'h00;      memory[48224] <=  8'h00;      memory[48225] <=  8'h00;      memory[48226] <=  8'h00;      memory[48227] <=  8'h00;      memory[48228] <=  8'h00;      memory[48229] <=  8'h00;      memory[48230] <=  8'h00;      memory[48231] <=  8'h00;      memory[48232] <=  8'h00;      memory[48233] <=  8'h00;      memory[48234] <=  8'h00;      memory[48235] <=  8'h00;      memory[48236] <=  8'h00;      memory[48237] <=  8'h00;      memory[48238] <=  8'h00;      memory[48239] <=  8'h00;      memory[48240] <=  8'h00;      memory[48241] <=  8'h00;      memory[48242] <=  8'h00;      memory[48243] <=  8'h00;      memory[48244] <=  8'h00;      memory[48245] <=  8'h00;      memory[48246] <=  8'h00;      memory[48247] <=  8'h00;      memory[48248] <=  8'h00;      memory[48249] <=  8'h00;      memory[48250] <=  8'h00;      memory[48251] <=  8'h00;      memory[48252] <=  8'h00;      memory[48253] <=  8'h00;      memory[48254] <=  8'h00;      memory[48255] <=  8'h00;      memory[48256] <=  8'h00;      memory[48257] <=  8'h00;      memory[48258] <=  8'h00;      memory[48259] <=  8'h00;      memory[48260] <=  8'h00;      memory[48261] <=  8'h00;      memory[48262] <=  8'h00;      memory[48263] <=  8'h00;      memory[48264] <=  8'h00;      memory[48265] <=  8'h00;      memory[48266] <=  8'h00;      memory[48267] <=  8'h00;      memory[48268] <=  8'h00;      memory[48269] <=  8'h00;      memory[48270] <=  8'h00;      memory[48271] <=  8'h00;      memory[48272] <=  8'h00;      memory[48273] <=  8'h00;      memory[48274] <=  8'h00;      memory[48275] <=  8'h00;      memory[48276] <=  8'h00;      memory[48277] <=  8'h00;      memory[48278] <=  8'h00;      memory[48279] <=  8'h00;      memory[48280] <=  8'h00;      memory[48281] <=  8'h00;      memory[48282] <=  8'h00;      memory[48283] <=  8'h00;      memory[48284] <=  8'h00;      memory[48285] <=  8'h00;      memory[48286] <=  8'h00;      memory[48287] <=  8'h00;      memory[48288] <=  8'h00;      memory[48289] <=  8'h00;      memory[48290] <=  8'h00;      memory[48291] <=  8'h00;      memory[48292] <=  8'h00;      memory[48293] <=  8'h00;      memory[48294] <=  8'h00;      memory[48295] <=  8'h00;      memory[48296] <=  8'h00;      memory[48297] <=  8'h00;      memory[48298] <=  8'h00;      memory[48299] <=  8'h00;      memory[48300] <=  8'h00;      memory[48301] <=  8'h00;      memory[48302] <=  8'h00;      memory[48303] <=  8'h00;      memory[48304] <=  8'h00;      memory[48305] <=  8'h00;      memory[48306] <=  8'h00;      memory[48307] <=  8'h00;      memory[48308] <=  8'h00;      memory[48309] <=  8'h00;      memory[48310] <=  8'h00;      memory[48311] <=  8'h00;      memory[48312] <=  8'h00;      memory[48313] <=  8'h00;      memory[48314] <=  8'h00;      memory[48315] <=  8'h00;      memory[48316] <=  8'h00;      memory[48317] <=  8'h00;      memory[48318] <=  8'h00;      memory[48319] <=  8'h00;      memory[48320] <=  8'h00;      memory[48321] <=  8'h00;      memory[48322] <=  8'h00;      memory[48323] <=  8'h00;      memory[48324] <=  8'h00;      memory[48325] <=  8'h00;      memory[48326] <=  8'h00;      memory[48327] <=  8'h00;      memory[48328] <=  8'h00;      memory[48329] <=  8'h00;      memory[48330] <=  8'h00;      memory[48331] <=  8'h00;      memory[48332] <=  8'h00;      memory[48333] <=  8'h00;      memory[48334] <=  8'h00;      memory[48335] <=  8'h00;      memory[48336] <=  8'h00;      memory[48337] <=  8'h00;      memory[48338] <=  8'h00;      memory[48339] <=  8'h00;      memory[48340] <=  8'h00;      memory[48341] <=  8'h00;      memory[48342] <=  8'h00;      memory[48343] <=  8'h00;      memory[48344] <=  8'h00;      memory[48345] <=  8'h00;      memory[48346] <=  8'h00;      memory[48347] <=  8'h00;      memory[48348] <=  8'h00;      memory[48349] <=  8'h00;      memory[48350] <=  8'h00;      memory[48351] <=  8'h00;      memory[48352] <=  8'h00;      memory[48353] <=  8'h00;      memory[48354] <=  8'h00;      memory[48355] <=  8'h00;      memory[48356] <=  8'h00;      memory[48357] <=  8'h00;      memory[48358] <=  8'h00;      memory[48359] <=  8'h00;      memory[48360] <=  8'h00;      memory[48361] <=  8'h00;      memory[48362] <=  8'h00;      memory[48363] <=  8'h00;      memory[48364] <=  8'h00;      memory[48365] <=  8'h00;      memory[48366] <=  8'h00;      memory[48367] <=  8'h00;      memory[48368] <=  8'h00;      memory[48369] <=  8'h00;      memory[48370] <=  8'h00;      memory[48371] <=  8'h00;      memory[48372] <=  8'h00;      memory[48373] <=  8'h00;      memory[48374] <=  8'h00;      memory[48375] <=  8'h00;      memory[48376] <=  8'h00;      memory[48377] <=  8'h00;      memory[48378] <=  8'h00;      memory[48379] <=  8'h00;      memory[48380] <=  8'h00;      memory[48381] <=  8'h00;      memory[48382] <=  8'h00;      memory[48383] <=  8'h00;      memory[48384] <=  8'h00;      memory[48385] <=  8'h00;      memory[48386] <=  8'h00;      memory[48387] <=  8'h00;      memory[48388] <=  8'h00;      memory[48389] <=  8'h00;      memory[48390] <=  8'h00;      memory[48391] <=  8'h00;      memory[48392] <=  8'h00;      memory[48393] <=  8'h00;      memory[48394] <=  8'h00;      memory[48395] <=  8'h00;      memory[48396] <=  8'h00;      memory[48397] <=  8'h00;      memory[48398] <=  8'h00;      memory[48399] <=  8'h00;      memory[48400] <=  8'h00;      memory[48401] <=  8'h00;      memory[48402] <=  8'h00;      memory[48403] <=  8'h00;      memory[48404] <=  8'h00;      memory[48405] <=  8'h00;      memory[48406] <=  8'h00;      memory[48407] <=  8'h00;      memory[48408] <=  8'h00;      memory[48409] <=  8'h00;      memory[48410] <=  8'h00;      memory[48411] <=  8'h00;      memory[48412] <=  8'h00;      memory[48413] <=  8'h00;      memory[48414] <=  8'h00;      memory[48415] <=  8'h00;      memory[48416] <=  8'h00;      memory[48417] <=  8'h00;      memory[48418] <=  8'h00;      memory[48419] <=  8'h00;      memory[48420] <=  8'h00;      memory[48421] <=  8'h00;      memory[48422] <=  8'h00;      memory[48423] <=  8'h00;      memory[48424] <=  8'h00;      memory[48425] <=  8'h00;      memory[48426] <=  8'h00;      memory[48427] <=  8'h00;      memory[48428] <=  8'h00;      memory[48429] <=  8'h00;      memory[48430] <=  8'h00;      memory[48431] <=  8'h00;      memory[48432] <=  8'h00;      memory[48433] <=  8'h00;      memory[48434] <=  8'h00;      memory[48435] <=  8'h00;      memory[48436] <=  8'h00;      memory[48437] <=  8'h00;      memory[48438] <=  8'h00;      memory[48439] <=  8'h00;      memory[48440] <=  8'h00;      memory[48441] <=  8'h00;      memory[48442] <=  8'h00;      memory[48443] <=  8'h00;      memory[48444] <=  8'h00;      memory[48445] <=  8'h00;      memory[48446] <=  8'h00;      memory[48447] <=  8'h00;      memory[48448] <=  8'h00;      memory[48449] <=  8'h00;      memory[48450] <=  8'h00;      memory[48451] <=  8'h00;      memory[48452] <=  8'h00;      memory[48453] <=  8'h00;      memory[48454] <=  8'h00;      memory[48455] <=  8'h00;      memory[48456] <=  8'h00;      memory[48457] <=  8'h00;      memory[48458] <=  8'h00;      memory[48459] <=  8'h00;      memory[48460] <=  8'h00;      memory[48461] <=  8'h00;      memory[48462] <=  8'h00;      memory[48463] <=  8'h00;      memory[48464] <=  8'h00;      memory[48465] <=  8'h00;      memory[48466] <=  8'h00;      memory[48467] <=  8'h00;      memory[48468] <=  8'h00;      memory[48469] <=  8'h00;      memory[48470] <=  8'h00;      memory[48471] <=  8'h00;      memory[48472] <=  8'h00;      memory[48473] <=  8'h00;      memory[48474] <=  8'h00;      memory[48475] <=  8'h00;      memory[48476] <=  8'h00;      memory[48477] <=  8'h00;      memory[48478] <=  8'h00;      memory[48479] <=  8'h00;      memory[48480] <=  8'h00;      memory[48481] <=  8'h00;      memory[48482] <=  8'h00;      memory[48483] <=  8'h00;      memory[48484] <=  8'h00;      memory[48485] <=  8'h00;      memory[48486] <=  8'h00;      memory[48487] <=  8'h00;      memory[48488] <=  8'h00;      memory[48489] <=  8'h00;      memory[48490] <=  8'h00;      memory[48491] <=  8'h00;      memory[48492] <=  8'h00;      memory[48493] <=  8'h00;      memory[48494] <=  8'h00;      memory[48495] <=  8'h00;      memory[48496] <=  8'h00;      memory[48497] <=  8'h00;      memory[48498] <=  8'h00;      memory[48499] <=  8'h00;      memory[48500] <=  8'h00;      memory[48501] <=  8'h00;      memory[48502] <=  8'h00;      memory[48503] <=  8'h00;      memory[48504] <=  8'h00;      memory[48505] <=  8'h00;      memory[48506] <=  8'h00;      memory[48507] <=  8'h00;      memory[48508] <=  8'h00;      memory[48509] <=  8'h00;      memory[48510] <=  8'h00;      memory[48511] <=  8'h00;      memory[48512] <=  8'h00;      memory[48513] <=  8'h00;      memory[48514] <=  8'h00;      memory[48515] <=  8'h00;      memory[48516] <=  8'h00;      memory[48517] <=  8'h00;      memory[48518] <=  8'h00;      memory[48519] <=  8'h00;      memory[48520] <=  8'h00;      memory[48521] <=  8'h00;      memory[48522] <=  8'h00;      memory[48523] <=  8'h00;      memory[48524] <=  8'h00;      memory[48525] <=  8'h00;      memory[48526] <=  8'h00;      memory[48527] <=  8'h00;      memory[48528] <=  8'h00;      memory[48529] <=  8'h00;      memory[48530] <=  8'h00;      memory[48531] <=  8'h00;      memory[48532] <=  8'h00;      memory[48533] <=  8'h00;      memory[48534] <=  8'h00;      memory[48535] <=  8'h00;      memory[48536] <=  8'h00;      memory[48537] <=  8'h00;      memory[48538] <=  8'h00;      memory[48539] <=  8'h00;      memory[48540] <=  8'h00;      memory[48541] <=  8'h00;      memory[48542] <=  8'h00;      memory[48543] <=  8'h00;      memory[48544] <=  8'h00;      memory[48545] <=  8'h00;      memory[48546] <=  8'h00;      memory[48547] <=  8'h00;      memory[48548] <=  8'h00;      memory[48549] <=  8'h00;      memory[48550] <=  8'h00;      memory[48551] <=  8'h00;      memory[48552] <=  8'h00;      memory[48553] <=  8'h00;      memory[48554] <=  8'h00;      memory[48555] <=  8'h00;      memory[48556] <=  8'h00;      memory[48557] <=  8'h00;      memory[48558] <=  8'h00;      memory[48559] <=  8'h00;      memory[48560] <=  8'h00;      memory[48561] <=  8'h00;      memory[48562] <=  8'h00;      memory[48563] <=  8'h00;      memory[48564] <=  8'h00;      memory[48565] <=  8'h00;      memory[48566] <=  8'h00;      memory[48567] <=  8'h00;      memory[48568] <=  8'h00;      memory[48569] <=  8'h00;      memory[48570] <=  8'h00;      memory[48571] <=  8'h00;      memory[48572] <=  8'h00;      memory[48573] <=  8'h00;      memory[48574] <=  8'h00;      memory[48575] <=  8'h00;      memory[48576] <=  8'h00;      memory[48577] <=  8'h00;      memory[48578] <=  8'h00;      memory[48579] <=  8'h00;      memory[48580] <=  8'h00;      memory[48581] <=  8'h00;      memory[48582] <=  8'h00;      memory[48583] <=  8'h00;      memory[48584] <=  8'h00;      memory[48585] <=  8'h00;      memory[48586] <=  8'h00;      memory[48587] <=  8'h00;      memory[48588] <=  8'h00;      memory[48589] <=  8'h00;      memory[48590] <=  8'h00;      memory[48591] <=  8'h00;      memory[48592] <=  8'h00;      memory[48593] <=  8'h00;      memory[48594] <=  8'h00;      memory[48595] <=  8'h00;      memory[48596] <=  8'h00;      memory[48597] <=  8'h00;      memory[48598] <=  8'h00;      memory[48599] <=  8'h00;      memory[48600] <=  8'h00;      memory[48601] <=  8'h00;      memory[48602] <=  8'h00;      memory[48603] <=  8'h00;      memory[48604] <=  8'h00;      memory[48605] <=  8'h00;      memory[48606] <=  8'h00;      memory[48607] <=  8'h00;      memory[48608] <=  8'h00;      memory[48609] <=  8'h00;      memory[48610] <=  8'h00;      memory[48611] <=  8'h00;      memory[48612] <=  8'h00;      memory[48613] <=  8'h00;      memory[48614] <=  8'h00;      memory[48615] <=  8'h00;      memory[48616] <=  8'h00;      memory[48617] <=  8'h00;      memory[48618] <=  8'h00;      memory[48619] <=  8'h00;      memory[48620] <=  8'h00;      memory[48621] <=  8'h00;      memory[48622] <=  8'h00;      memory[48623] <=  8'h00;      memory[48624] <=  8'h00;      memory[48625] <=  8'h00;      memory[48626] <=  8'h00;      memory[48627] <=  8'h00;      memory[48628] <=  8'h00;      memory[48629] <=  8'h00;      memory[48630] <=  8'h00;      memory[48631] <=  8'h00;      memory[48632] <=  8'h00;      memory[48633] <=  8'h00;      memory[48634] <=  8'h00;      memory[48635] <=  8'h00;      memory[48636] <=  8'h00;      memory[48637] <=  8'h00;      memory[48638] <=  8'h00;      memory[48639] <=  8'h00;      memory[48640] <=  8'h00;      memory[48641] <=  8'h00;      memory[48642] <=  8'h00;      memory[48643] <=  8'h00;      memory[48644] <=  8'h00;      memory[48645] <=  8'h00;      memory[48646] <=  8'h00;      memory[48647] <=  8'h00;      memory[48648] <=  8'h00;      memory[48649] <=  8'h00;      memory[48650] <=  8'h00;      memory[48651] <=  8'h00;      memory[48652] <=  8'h00;      memory[48653] <=  8'h00;      memory[48654] <=  8'h00;      memory[48655] <=  8'h00;      memory[48656] <=  8'h00;      memory[48657] <=  8'h00;      memory[48658] <=  8'h00;      memory[48659] <=  8'h00;      memory[48660] <=  8'h00;      memory[48661] <=  8'h00;      memory[48662] <=  8'h00;      memory[48663] <=  8'h00;      memory[48664] <=  8'h00;      memory[48665] <=  8'h00;      memory[48666] <=  8'h00;      memory[48667] <=  8'h00;      memory[48668] <=  8'h00;      memory[48669] <=  8'h00;      memory[48670] <=  8'h00;      memory[48671] <=  8'h00;      memory[48672] <=  8'h00;      memory[48673] <=  8'h00;      memory[48674] <=  8'h00;      memory[48675] <=  8'h00;      memory[48676] <=  8'h00;      memory[48677] <=  8'h00;      memory[48678] <=  8'h00;      memory[48679] <=  8'h00;      memory[48680] <=  8'h00;      memory[48681] <=  8'h00;      memory[48682] <=  8'h00;      memory[48683] <=  8'h00;      memory[48684] <=  8'h00;      memory[48685] <=  8'h00;      memory[48686] <=  8'h00;      memory[48687] <=  8'h00;      memory[48688] <=  8'h00;      memory[48689] <=  8'h00;      memory[48690] <=  8'h00;      memory[48691] <=  8'h00;      memory[48692] <=  8'h00;      memory[48693] <=  8'h00;      memory[48694] <=  8'h00;      memory[48695] <=  8'h00;      memory[48696] <=  8'h00;      memory[48697] <=  8'h00;      memory[48698] <=  8'h00;      memory[48699] <=  8'h00;      memory[48700] <=  8'h00;      memory[48701] <=  8'h00;      memory[48702] <=  8'h00;      memory[48703] <=  8'h00;      memory[48704] <=  8'h00;      memory[48705] <=  8'h00;      memory[48706] <=  8'h00;      memory[48707] <=  8'h00;      memory[48708] <=  8'h00;      memory[48709] <=  8'h00;      memory[48710] <=  8'h00;      memory[48711] <=  8'h00;      memory[48712] <=  8'h00;      memory[48713] <=  8'h00;      memory[48714] <=  8'h00;      memory[48715] <=  8'h00;      memory[48716] <=  8'h00;      memory[48717] <=  8'h00;      memory[48718] <=  8'h00;      memory[48719] <=  8'h00;      memory[48720] <=  8'h00;      memory[48721] <=  8'h00;      memory[48722] <=  8'h00;      memory[48723] <=  8'h00;      memory[48724] <=  8'h00;      memory[48725] <=  8'h00;      memory[48726] <=  8'h00;      memory[48727] <=  8'h00;      memory[48728] <=  8'h00;      memory[48729] <=  8'h00;      memory[48730] <=  8'h00;      memory[48731] <=  8'h00;      memory[48732] <=  8'h00;      memory[48733] <=  8'h00;      memory[48734] <=  8'h00;      memory[48735] <=  8'h00;      memory[48736] <=  8'h00;      memory[48737] <=  8'h00;      memory[48738] <=  8'h00;      memory[48739] <=  8'h00;      memory[48740] <=  8'h00;      memory[48741] <=  8'h00;      memory[48742] <=  8'h00;      memory[48743] <=  8'h00;      memory[48744] <=  8'h00;      memory[48745] <=  8'h00;      memory[48746] <=  8'h00;      memory[48747] <=  8'h00;      memory[48748] <=  8'h00;      memory[48749] <=  8'h00;      memory[48750] <=  8'h00;      memory[48751] <=  8'h00;      memory[48752] <=  8'h00;      memory[48753] <=  8'h00;      memory[48754] <=  8'h00;      memory[48755] <=  8'h00;      memory[48756] <=  8'h00;      memory[48757] <=  8'h00;      memory[48758] <=  8'h00;      memory[48759] <=  8'h00;      memory[48760] <=  8'h00;      memory[48761] <=  8'h00;      memory[48762] <=  8'h00;      memory[48763] <=  8'h00;      memory[48764] <=  8'h00;      memory[48765] <=  8'h00;      memory[48766] <=  8'h00;      memory[48767] <=  8'h00;      memory[48768] <=  8'h00;      memory[48769] <=  8'h00;      memory[48770] <=  8'h00;      memory[48771] <=  8'h00;      memory[48772] <=  8'h00;      memory[48773] <=  8'h00;      memory[48774] <=  8'h00;      memory[48775] <=  8'h00;      memory[48776] <=  8'h00;      memory[48777] <=  8'h00;      memory[48778] <=  8'h00;      memory[48779] <=  8'h00;      memory[48780] <=  8'h00;      memory[48781] <=  8'h00;      memory[48782] <=  8'h00;      memory[48783] <=  8'h00;      memory[48784] <=  8'h00;      memory[48785] <=  8'h00;      memory[48786] <=  8'h00;      memory[48787] <=  8'h00;      memory[48788] <=  8'h00;      memory[48789] <=  8'h00;      memory[48790] <=  8'h00;      memory[48791] <=  8'h00;      memory[48792] <=  8'h00;      memory[48793] <=  8'h00;      memory[48794] <=  8'h00;      memory[48795] <=  8'h00;      memory[48796] <=  8'h00;      memory[48797] <=  8'h00;      memory[48798] <=  8'h00;      memory[48799] <=  8'h00;      memory[48800] <=  8'h00;      memory[48801] <=  8'h00;      memory[48802] <=  8'h00;      memory[48803] <=  8'h00;      memory[48804] <=  8'h00;      memory[48805] <=  8'h00;      memory[48806] <=  8'h00;      memory[48807] <=  8'h00;      memory[48808] <=  8'h00;      memory[48809] <=  8'h00;      memory[48810] <=  8'h00;      memory[48811] <=  8'h00;      memory[48812] <=  8'h00;      memory[48813] <=  8'h00;      memory[48814] <=  8'h00;      memory[48815] <=  8'h00;      memory[48816] <=  8'h00;      memory[48817] <=  8'h00;      memory[48818] <=  8'h00;      memory[48819] <=  8'h00;      memory[48820] <=  8'h00;      memory[48821] <=  8'h00;      memory[48822] <=  8'h00;      memory[48823] <=  8'h00;      memory[48824] <=  8'h00;      memory[48825] <=  8'h00;      memory[48826] <=  8'h00;      memory[48827] <=  8'h00;      memory[48828] <=  8'h00;      memory[48829] <=  8'h00;      memory[48830] <=  8'h00;      memory[48831] <=  8'h00;      memory[48832] <=  8'h00;      memory[48833] <=  8'h00;      memory[48834] <=  8'h00;      memory[48835] <=  8'h00;      memory[48836] <=  8'h00;      memory[48837] <=  8'h00;      memory[48838] <=  8'h00;      memory[48839] <=  8'h00;      memory[48840] <=  8'h00;      memory[48841] <=  8'h00;      memory[48842] <=  8'h00;      memory[48843] <=  8'h00;      memory[48844] <=  8'h00;      memory[48845] <=  8'h00;      memory[48846] <=  8'h00;      memory[48847] <=  8'h00;      memory[48848] <=  8'h00;      memory[48849] <=  8'h00;      memory[48850] <=  8'h00;      memory[48851] <=  8'h00;      memory[48852] <=  8'h00;      memory[48853] <=  8'h00;      memory[48854] <=  8'h00;      memory[48855] <=  8'h00;      memory[48856] <=  8'h00;      memory[48857] <=  8'h00;      memory[48858] <=  8'h00;      memory[48859] <=  8'h00;      memory[48860] <=  8'h00;      memory[48861] <=  8'h00;      memory[48862] <=  8'h00;      memory[48863] <=  8'h00;      memory[48864] <=  8'h00;      memory[48865] <=  8'h00;      memory[48866] <=  8'h00;      memory[48867] <=  8'h00;      memory[48868] <=  8'h00;      memory[48869] <=  8'h00;      memory[48870] <=  8'h00;      memory[48871] <=  8'h00;      memory[48872] <=  8'h00;      memory[48873] <=  8'h00;      memory[48874] <=  8'h00;      memory[48875] <=  8'h00;      memory[48876] <=  8'h00;      memory[48877] <=  8'h00;      memory[48878] <=  8'h00;      memory[48879] <=  8'h00;      memory[48880] <=  8'h00;      memory[48881] <=  8'h00;      memory[48882] <=  8'h00;      memory[48883] <=  8'h00;      memory[48884] <=  8'h00;      memory[48885] <=  8'h00;      memory[48886] <=  8'h00;      memory[48887] <=  8'h00;      memory[48888] <=  8'h00;      memory[48889] <=  8'h00;      memory[48890] <=  8'h00;      memory[48891] <=  8'h00;      memory[48892] <=  8'h00;      memory[48893] <=  8'h00;      memory[48894] <=  8'h00;      memory[48895] <=  8'h00;      memory[48896] <=  8'h00;      memory[48897] <=  8'h00;      memory[48898] <=  8'h00;      memory[48899] <=  8'h00;      memory[48900] <=  8'h00;      memory[48901] <=  8'h00;      memory[48902] <=  8'h00;      memory[48903] <=  8'h00;      memory[48904] <=  8'h00;      memory[48905] <=  8'h00;      memory[48906] <=  8'h00;      memory[48907] <=  8'h00;      memory[48908] <=  8'h00;      memory[48909] <=  8'h00;      memory[48910] <=  8'h00;      memory[48911] <=  8'h00;      memory[48912] <=  8'h00;      memory[48913] <=  8'h00;      memory[48914] <=  8'h00;      memory[48915] <=  8'h00;      memory[48916] <=  8'h00;      memory[48917] <=  8'h00;      memory[48918] <=  8'h00;      memory[48919] <=  8'h00;      memory[48920] <=  8'h00;      memory[48921] <=  8'h00;      memory[48922] <=  8'h00;      memory[48923] <=  8'h00;      memory[48924] <=  8'h00;      memory[48925] <=  8'h00;      memory[48926] <=  8'h00;      memory[48927] <=  8'h00;      memory[48928] <=  8'h00;      memory[48929] <=  8'h00;      memory[48930] <=  8'h00;      memory[48931] <=  8'h00;      memory[48932] <=  8'h00;      memory[48933] <=  8'h00;      memory[48934] <=  8'h00;      memory[48935] <=  8'h00;      memory[48936] <=  8'h00;      memory[48937] <=  8'h00;      memory[48938] <=  8'h00;      memory[48939] <=  8'h00;      memory[48940] <=  8'h00;      memory[48941] <=  8'h00;      memory[48942] <=  8'h00;      memory[48943] <=  8'h00;      memory[48944] <=  8'h00;      memory[48945] <=  8'h00;      memory[48946] <=  8'h00;      memory[48947] <=  8'h00;      memory[48948] <=  8'h00;      memory[48949] <=  8'h00;      memory[48950] <=  8'h00;      memory[48951] <=  8'h00;      memory[48952] <=  8'h00;      memory[48953] <=  8'h00;      memory[48954] <=  8'h00;      memory[48955] <=  8'h00;      memory[48956] <=  8'h00;      memory[48957] <=  8'h00;      memory[48958] <=  8'h00;      memory[48959] <=  8'h00;      memory[48960] <=  8'h00;      memory[48961] <=  8'h00;      memory[48962] <=  8'h00;      memory[48963] <=  8'h00;      memory[48964] <=  8'h00;      memory[48965] <=  8'h00;      memory[48966] <=  8'h00;      memory[48967] <=  8'h00;      memory[48968] <=  8'h00;      memory[48969] <=  8'h00;      memory[48970] <=  8'h00;      memory[48971] <=  8'h00;      memory[48972] <=  8'h00;      memory[48973] <=  8'h00;      memory[48974] <=  8'h00;      memory[48975] <=  8'h00;      memory[48976] <=  8'h00;      memory[48977] <=  8'h00;      memory[48978] <=  8'h00;      memory[48979] <=  8'h00;      memory[48980] <=  8'h00;      memory[48981] <=  8'h00;      memory[48982] <=  8'h00;      memory[48983] <=  8'h00;      memory[48984] <=  8'h00;      memory[48985] <=  8'h00;      memory[48986] <=  8'h00;      memory[48987] <=  8'h00;      memory[48988] <=  8'h00;      memory[48989] <=  8'h00;      memory[48990] <=  8'h00;      memory[48991] <=  8'h00;      memory[48992] <=  8'h00;      memory[48993] <=  8'h00;      memory[48994] <=  8'h00;      memory[48995] <=  8'h00;      memory[48996] <=  8'h00;      memory[48997] <=  8'h00;      memory[48998] <=  8'h00;      memory[48999] <=  8'h00;      memory[49000] <=  8'h00;      memory[49001] <=  8'h00;      memory[49002] <=  8'h00;      memory[49003] <=  8'h00;      memory[49004] <=  8'h00;      memory[49005] <=  8'h00;      memory[49006] <=  8'h00;      memory[49007] <=  8'h00;      memory[49008] <=  8'h00;      memory[49009] <=  8'h00;      memory[49010] <=  8'h00;      memory[49011] <=  8'h00;      memory[49012] <=  8'h00;      memory[49013] <=  8'h00;      memory[49014] <=  8'h00;      memory[49015] <=  8'h00;      memory[49016] <=  8'h00;      memory[49017] <=  8'h00;      memory[49018] <=  8'h00;      memory[49019] <=  8'h00;      memory[49020] <=  8'h00;      memory[49021] <=  8'h00;      memory[49022] <=  8'h00;      memory[49023] <=  8'h00;      memory[49024] <=  8'h00;      memory[49025] <=  8'h00;      memory[49026] <=  8'h00;      memory[49027] <=  8'h00;      memory[49028] <=  8'h00;      memory[49029] <=  8'h00;      memory[49030] <=  8'h00;      memory[49031] <=  8'h00;      memory[49032] <=  8'h00;      memory[49033] <=  8'h00;      memory[49034] <=  8'h00;      memory[49035] <=  8'h00;      memory[49036] <=  8'h00;      memory[49037] <=  8'h00;      memory[49038] <=  8'h00;      memory[49039] <=  8'h00;      memory[49040] <=  8'h00;      memory[49041] <=  8'h00;      memory[49042] <=  8'h00;      memory[49043] <=  8'h00;      memory[49044] <=  8'h00;      memory[49045] <=  8'h00;      memory[49046] <=  8'h00;      memory[49047] <=  8'h00;      memory[49048] <=  8'h00;      memory[49049] <=  8'h00;      memory[49050] <=  8'h00;      memory[49051] <=  8'h00;      memory[49052] <=  8'h00;      memory[49053] <=  8'h00;      memory[49054] <=  8'h00;      memory[49055] <=  8'h00;      memory[49056] <=  8'h00;      memory[49057] <=  8'h00;      memory[49058] <=  8'h00;      memory[49059] <=  8'h00;      memory[49060] <=  8'h00;      memory[49061] <=  8'h00;      memory[49062] <=  8'h00;      memory[49063] <=  8'h00;      memory[49064] <=  8'h00;      memory[49065] <=  8'h00;      memory[49066] <=  8'h00;      memory[49067] <=  8'h00;      memory[49068] <=  8'h00;      memory[49069] <=  8'h00;      memory[49070] <=  8'h00;      memory[49071] <=  8'h00;      memory[49072] <=  8'h00;      memory[49073] <=  8'h00;      memory[49074] <=  8'h00;      memory[49075] <=  8'h00;      memory[49076] <=  8'h00;      memory[49077] <=  8'h00;      memory[49078] <=  8'h00;      memory[49079] <=  8'h00;      memory[49080] <=  8'h00;      memory[49081] <=  8'h00;      memory[49082] <=  8'h00;      memory[49083] <=  8'h00;      memory[49084] <=  8'h00;      memory[49085] <=  8'h00;      memory[49086] <=  8'h00;      memory[49087] <=  8'h00;      memory[49088] <=  8'h00;      memory[49089] <=  8'h00;      memory[49090] <=  8'h00;      memory[49091] <=  8'h00;      memory[49092] <=  8'h00;      memory[49093] <=  8'h00;      memory[49094] <=  8'h00;      memory[49095] <=  8'h00;      memory[49096] <=  8'h00;      memory[49097] <=  8'h00;      memory[49098] <=  8'h00;      memory[49099] <=  8'h00;      memory[49100] <=  8'h00;      memory[49101] <=  8'h00;      memory[49102] <=  8'h00;      memory[49103] <=  8'h00;      memory[49104] <=  8'h00;      memory[49105] <=  8'h00;      memory[49106] <=  8'h00;      memory[49107] <=  8'h00;      memory[49108] <=  8'h00;      memory[49109] <=  8'h00;      memory[49110] <=  8'h00;      memory[49111] <=  8'h00;      memory[49112] <=  8'h00;      memory[49113] <=  8'h00;      memory[49114] <=  8'h00;      memory[49115] <=  8'h00;      memory[49116] <=  8'h00;      memory[49117] <=  8'h00;      memory[49118] <=  8'h00;      memory[49119] <=  8'h00;      memory[49120] <=  8'h00;      memory[49121] <=  8'h00;      memory[49122] <=  8'h00;      memory[49123] <=  8'h00;      memory[49124] <=  8'h00;      memory[49125] <=  8'h00;      memory[49126] <=  8'h00;      memory[49127] <=  8'h00;      memory[49128] <=  8'h00;      memory[49129] <=  8'h00;      memory[49130] <=  8'h00;      memory[49131] <=  8'h00;      memory[49132] <=  8'h00;      memory[49133] <=  8'h00;      memory[49134] <=  8'h00;      memory[49135] <=  8'h00;      memory[49136] <=  8'h00;      memory[49137] <=  8'h00;      memory[49138] <=  8'h00;      memory[49139] <=  8'h00;      memory[49140] <=  8'h00;      memory[49141] <=  8'h00;      memory[49142] <=  8'h00;      memory[49143] <=  8'h00;      memory[49144] <=  8'h00;      memory[49145] <=  8'h00;      memory[49146] <=  8'h00;      memory[49147] <=  8'h00;      memory[49148] <=  8'h00;      memory[49149] <=  8'h00;      memory[49150] <=  8'h00;      memory[49151] <=  8'h00;      memory[49152] <=  8'h00;      memory[49153] <=  8'h00;      memory[49154] <=  8'h00;      memory[49155] <=  8'h00;      memory[49156] <=  8'h00;      memory[49157] <=  8'h00;      memory[49158] <=  8'h00;      memory[49159] <=  8'h00;      memory[49160] <=  8'h00;      memory[49161] <=  8'h00;      memory[49162] <=  8'h00;      memory[49163] <=  8'h00;      memory[49164] <=  8'h00;      memory[49165] <=  8'h00;      memory[49166] <=  8'h00;      memory[49167] <=  8'h00;      memory[49168] <=  8'h00;      memory[49169] <=  8'h00;      memory[49170] <=  8'h00;      memory[49171] <=  8'h00;      memory[49172] <=  8'h00;      memory[49173] <=  8'h00;      memory[49174] <=  8'h00;      memory[49175] <=  8'h00;      memory[49176] <=  8'h00;      memory[49177] <=  8'h00;      memory[49178] <=  8'h00;      memory[49179] <=  8'h00;      memory[49180] <=  8'h00;      memory[49181] <=  8'h00;      memory[49182] <=  8'h00;      memory[49183] <=  8'h00;      memory[49184] <=  8'h00;      memory[49185] <=  8'h00;      memory[49186] <=  8'h00;      memory[49187] <=  8'h00;      memory[49188] <=  8'h00;      memory[49189] <=  8'h00;      memory[49190] <=  8'h00;      memory[49191] <=  8'h00;      memory[49192] <=  8'h00;      memory[49193] <=  8'h00;      memory[49194] <=  8'h00;      memory[49195] <=  8'h00;      memory[49196] <=  8'h00;      memory[49197] <=  8'h00;      memory[49198] <=  8'h00;      memory[49199] <=  8'h00;      memory[49200] <=  8'h00;      memory[49201] <=  8'h00;      memory[49202] <=  8'h00;      memory[49203] <=  8'h00;      memory[49204] <=  8'h00;      memory[49205] <=  8'h00;      memory[49206] <=  8'h00;      memory[49207] <=  8'h00;      memory[49208] <=  8'h00;      memory[49209] <=  8'h00;      memory[49210] <=  8'h00;      memory[49211] <=  8'h00;      memory[49212] <=  8'h00;      memory[49213] <=  8'h00;      memory[49214] <=  8'h00;      memory[49215] <=  8'h00;      memory[49216] <=  8'h00;      memory[49217] <=  8'h00;      memory[49218] <=  8'h00;      memory[49219] <=  8'h00;      memory[49220] <=  8'h00;      memory[49221] <=  8'h00;      memory[49222] <=  8'h00;      memory[49223] <=  8'h00;      memory[49224] <=  8'h00;      memory[49225] <=  8'h00;      memory[49226] <=  8'h00;      memory[49227] <=  8'h00;      memory[49228] <=  8'h00;      memory[49229] <=  8'h00;      memory[49230] <=  8'h00;      memory[49231] <=  8'h00;      memory[49232] <=  8'h00;      memory[49233] <=  8'h00;      memory[49234] <=  8'h00;      memory[49235] <=  8'h00;      memory[49236] <=  8'h00;      memory[49237] <=  8'h00;      memory[49238] <=  8'h00;      memory[49239] <=  8'h00;      memory[49240] <=  8'h00;      memory[49241] <=  8'h00;      memory[49242] <=  8'h00;      memory[49243] <=  8'h00;      memory[49244] <=  8'h00;      memory[49245] <=  8'h00;      memory[49246] <=  8'h00;      memory[49247] <=  8'h00;      memory[49248] <=  8'h00;      memory[49249] <=  8'h00;      memory[49250] <=  8'h00;      memory[49251] <=  8'h00;      memory[49252] <=  8'h00;      memory[49253] <=  8'h00;      memory[49254] <=  8'h00;      memory[49255] <=  8'h00;      memory[49256] <=  8'h00;      memory[49257] <=  8'h00;      memory[49258] <=  8'h00;      memory[49259] <=  8'h00;      memory[49260] <=  8'h00;      memory[49261] <=  8'h00;      memory[49262] <=  8'h00;      memory[49263] <=  8'h00;      memory[49264] <=  8'h00;      memory[49265] <=  8'h00;      memory[49266] <=  8'h00;      memory[49267] <=  8'h00;      memory[49268] <=  8'h00;      memory[49269] <=  8'h00;      memory[49270] <=  8'h00;      memory[49271] <=  8'h00;      memory[49272] <=  8'h00;      memory[49273] <=  8'h00;      memory[49274] <=  8'h00;      memory[49275] <=  8'h00;      memory[49276] <=  8'h00;      memory[49277] <=  8'h00;      memory[49278] <=  8'h00;      memory[49279] <=  8'h00;      memory[49280] <=  8'h00;      memory[49281] <=  8'h00;      memory[49282] <=  8'h00;      memory[49283] <=  8'h00;      memory[49284] <=  8'h00;      memory[49285] <=  8'h00;      memory[49286] <=  8'h00;      memory[49287] <=  8'h00;      memory[49288] <=  8'h00;      memory[49289] <=  8'h00;      memory[49290] <=  8'h00;      memory[49291] <=  8'h00;      memory[49292] <=  8'h00;      memory[49293] <=  8'h00;      memory[49294] <=  8'h00;      memory[49295] <=  8'h00;      memory[49296] <=  8'h00;      memory[49297] <=  8'h00;      memory[49298] <=  8'h00;      memory[49299] <=  8'h00;      memory[49300] <=  8'h00;      memory[49301] <=  8'h00;      memory[49302] <=  8'h00;      memory[49303] <=  8'h00;      memory[49304] <=  8'h00;      memory[49305] <=  8'h00;      memory[49306] <=  8'h00;      memory[49307] <=  8'h00;      memory[49308] <=  8'h00;      memory[49309] <=  8'h00;      memory[49310] <=  8'h00;      memory[49311] <=  8'h00;      memory[49312] <=  8'h00;      memory[49313] <=  8'h00;      memory[49314] <=  8'h00;      memory[49315] <=  8'h00;      memory[49316] <=  8'h00;      memory[49317] <=  8'h00;      memory[49318] <=  8'h00;      memory[49319] <=  8'h00;      memory[49320] <=  8'h00;      memory[49321] <=  8'h00;      memory[49322] <=  8'h00;      memory[49323] <=  8'h00;      memory[49324] <=  8'h00;      memory[49325] <=  8'h00;      memory[49326] <=  8'h00;      memory[49327] <=  8'h00;      memory[49328] <=  8'h00;      memory[49329] <=  8'h00;      memory[49330] <=  8'h00;      memory[49331] <=  8'h00;      memory[49332] <=  8'h00;      memory[49333] <=  8'h00;      memory[49334] <=  8'h00;      memory[49335] <=  8'h00;      memory[49336] <=  8'h00;      memory[49337] <=  8'h00;      memory[49338] <=  8'h00;      memory[49339] <=  8'h00;      memory[49340] <=  8'h00;      memory[49341] <=  8'h00;      memory[49342] <=  8'h00;      memory[49343] <=  8'h00;      memory[49344] <=  8'h00;      memory[49345] <=  8'h00;      memory[49346] <=  8'h00;      memory[49347] <=  8'h00;      memory[49348] <=  8'h00;      memory[49349] <=  8'h00;      memory[49350] <=  8'h00;      memory[49351] <=  8'h00;      memory[49352] <=  8'h00;      memory[49353] <=  8'h00;      memory[49354] <=  8'h00;      memory[49355] <=  8'h00;      memory[49356] <=  8'h00;      memory[49357] <=  8'h00;      memory[49358] <=  8'h00;      memory[49359] <=  8'h00;      memory[49360] <=  8'h00;      memory[49361] <=  8'h00;      memory[49362] <=  8'h00;      memory[49363] <=  8'h00;      memory[49364] <=  8'h00;      memory[49365] <=  8'h00;      memory[49366] <=  8'h00;      memory[49367] <=  8'h00;      memory[49368] <=  8'h00;      memory[49369] <=  8'h00;      memory[49370] <=  8'h00;      memory[49371] <=  8'h00;      memory[49372] <=  8'h00;      memory[49373] <=  8'h00;      memory[49374] <=  8'h00;      memory[49375] <=  8'h00;      memory[49376] <=  8'h00;      memory[49377] <=  8'h00;      memory[49378] <=  8'h00;      memory[49379] <=  8'h00;      memory[49380] <=  8'h00;      memory[49381] <=  8'h00;      memory[49382] <=  8'h00;      memory[49383] <=  8'h00;      memory[49384] <=  8'h00;      memory[49385] <=  8'h00;      memory[49386] <=  8'h00;      memory[49387] <=  8'h00;      memory[49388] <=  8'h00;      memory[49389] <=  8'h00;      memory[49390] <=  8'h00;      memory[49391] <=  8'h00;      memory[49392] <=  8'h00;      memory[49393] <=  8'h00;      memory[49394] <=  8'h00;      memory[49395] <=  8'h00;      memory[49396] <=  8'h00;      memory[49397] <=  8'h00;      memory[49398] <=  8'h00;      memory[49399] <=  8'h00;      memory[49400] <=  8'h00;      memory[49401] <=  8'h00;      memory[49402] <=  8'h00;      memory[49403] <=  8'h00;      memory[49404] <=  8'h00;      memory[49405] <=  8'h00;      memory[49406] <=  8'h00;      memory[49407] <=  8'h00;      memory[49408] <=  8'h00;      memory[49409] <=  8'h00;      memory[49410] <=  8'h00;      memory[49411] <=  8'h00;      memory[49412] <=  8'h00;      memory[49413] <=  8'h00;      memory[49414] <=  8'h00;      memory[49415] <=  8'h00;      memory[49416] <=  8'h00;      memory[49417] <=  8'h00;      memory[49418] <=  8'h00;      memory[49419] <=  8'h00;      memory[49420] <=  8'h00;      memory[49421] <=  8'h00;      memory[49422] <=  8'h00;      memory[49423] <=  8'h00;      memory[49424] <=  8'h00;      memory[49425] <=  8'h00;      memory[49426] <=  8'h00;      memory[49427] <=  8'h00;      memory[49428] <=  8'h00;      memory[49429] <=  8'h00;      memory[49430] <=  8'h00;      memory[49431] <=  8'h00;      memory[49432] <=  8'h00;      memory[49433] <=  8'h00;      memory[49434] <=  8'h00;      memory[49435] <=  8'h00;      memory[49436] <=  8'h00;      memory[49437] <=  8'h00;      memory[49438] <=  8'h00;      memory[49439] <=  8'h00;      memory[49440] <=  8'h00;      memory[49441] <=  8'h00;      memory[49442] <=  8'h00;      memory[49443] <=  8'h00;      memory[49444] <=  8'h00;      memory[49445] <=  8'h00;      memory[49446] <=  8'h00;      memory[49447] <=  8'h00;      memory[49448] <=  8'h00;      memory[49449] <=  8'h00;      memory[49450] <=  8'h00;      memory[49451] <=  8'h00;      memory[49452] <=  8'h00;      memory[49453] <=  8'h00;      memory[49454] <=  8'h00;      memory[49455] <=  8'h00;      memory[49456] <=  8'h00;      memory[49457] <=  8'h00;      memory[49458] <=  8'h00;      memory[49459] <=  8'h00;      memory[49460] <=  8'h00;      memory[49461] <=  8'h00;      memory[49462] <=  8'h00;      memory[49463] <=  8'h00;      memory[49464] <=  8'h00;      memory[49465] <=  8'h00;      memory[49466] <=  8'h00;      memory[49467] <=  8'h00;      memory[49468] <=  8'h00;      memory[49469] <=  8'h00;      memory[49470] <=  8'h00;      memory[49471] <=  8'h00;      memory[49472] <=  8'h00;      memory[49473] <=  8'h00;      memory[49474] <=  8'h00;      memory[49475] <=  8'h00;      memory[49476] <=  8'h00;      memory[49477] <=  8'h00;      memory[49478] <=  8'h00;      memory[49479] <=  8'h00;      memory[49480] <=  8'h00;      memory[49481] <=  8'h00;      memory[49482] <=  8'h00;      memory[49483] <=  8'h00;      memory[49484] <=  8'h00;      memory[49485] <=  8'h00;      memory[49486] <=  8'h00;      memory[49487] <=  8'h00;      memory[49488] <=  8'h00;      memory[49489] <=  8'h00;      memory[49490] <=  8'h00;      memory[49491] <=  8'h00;      memory[49492] <=  8'h00;      memory[49493] <=  8'h00;      memory[49494] <=  8'h00;      memory[49495] <=  8'h00;      memory[49496] <=  8'h00;      memory[49497] <=  8'h00;      memory[49498] <=  8'h00;      memory[49499] <=  8'h00;      memory[49500] <=  8'h00;      memory[49501] <=  8'h00;      memory[49502] <=  8'h00;      memory[49503] <=  8'h00;      memory[49504] <=  8'h00;      memory[49505] <=  8'h00;      memory[49506] <=  8'h00;      memory[49507] <=  8'h00;      memory[49508] <=  8'h00;      memory[49509] <=  8'h00;      memory[49510] <=  8'h00;      memory[49511] <=  8'h00;      memory[49512] <=  8'h00;      memory[49513] <=  8'h00;      memory[49514] <=  8'h00;      memory[49515] <=  8'h00;      memory[49516] <=  8'h00;      memory[49517] <=  8'h00;      memory[49518] <=  8'h00;      memory[49519] <=  8'h00;      memory[49520] <=  8'h00;      memory[49521] <=  8'h00;      memory[49522] <=  8'h00;      memory[49523] <=  8'h00;      memory[49524] <=  8'h00;      memory[49525] <=  8'h00;      memory[49526] <=  8'h00;      memory[49527] <=  8'h00;      memory[49528] <=  8'h00;      memory[49529] <=  8'h00;      memory[49530] <=  8'h00;      memory[49531] <=  8'h00;      memory[49532] <=  8'h00;      memory[49533] <=  8'h00;      memory[49534] <=  8'h00;      memory[49535] <=  8'h00;      memory[49536] <=  8'h00;      memory[49537] <=  8'h00;      memory[49538] <=  8'h00;      memory[49539] <=  8'h00;      memory[49540] <=  8'h00;      memory[49541] <=  8'h00;      memory[49542] <=  8'h00;      memory[49543] <=  8'h00;      memory[49544] <=  8'h00;      memory[49545] <=  8'h00;      memory[49546] <=  8'h00;      memory[49547] <=  8'h00;      memory[49548] <=  8'h00;      memory[49549] <=  8'h00;      memory[49550] <=  8'h00;      memory[49551] <=  8'h00;      memory[49552] <=  8'h00;      memory[49553] <=  8'h00;      memory[49554] <=  8'h00;      memory[49555] <=  8'h00;      memory[49556] <=  8'h00;      memory[49557] <=  8'h00;      memory[49558] <=  8'h00;      memory[49559] <=  8'h00;      memory[49560] <=  8'h00;      memory[49561] <=  8'h00;      memory[49562] <=  8'h00;      memory[49563] <=  8'h00;      memory[49564] <=  8'h00;      memory[49565] <=  8'h00;      memory[49566] <=  8'h00;      memory[49567] <=  8'h00;      memory[49568] <=  8'h00;      memory[49569] <=  8'h00;      memory[49570] <=  8'h00;      memory[49571] <=  8'h00;      memory[49572] <=  8'h00;      memory[49573] <=  8'h00;      memory[49574] <=  8'h00;      memory[49575] <=  8'h00;      memory[49576] <=  8'h00;      memory[49577] <=  8'h00;      memory[49578] <=  8'h00;      memory[49579] <=  8'h00;      memory[49580] <=  8'h00;      memory[49581] <=  8'h00;      memory[49582] <=  8'h00;      memory[49583] <=  8'h00;      memory[49584] <=  8'h00;      memory[49585] <=  8'h00;      memory[49586] <=  8'h00;      memory[49587] <=  8'h00;      memory[49588] <=  8'h00;      memory[49589] <=  8'h00;      memory[49590] <=  8'h00;      memory[49591] <=  8'h00;      memory[49592] <=  8'h00;      memory[49593] <=  8'h00;      memory[49594] <=  8'h00;      memory[49595] <=  8'h00;      memory[49596] <=  8'h00;      memory[49597] <=  8'h00;      memory[49598] <=  8'h00;      memory[49599] <=  8'h00;      memory[49600] <=  8'h00;      memory[49601] <=  8'h00;      memory[49602] <=  8'h00;      memory[49603] <=  8'h00;      memory[49604] <=  8'h00;      memory[49605] <=  8'h00;      memory[49606] <=  8'h00;      memory[49607] <=  8'h00;      memory[49608] <=  8'h00;      memory[49609] <=  8'h00;      memory[49610] <=  8'h00;      memory[49611] <=  8'h00;      memory[49612] <=  8'h00;      memory[49613] <=  8'h00;      memory[49614] <=  8'h00;      memory[49615] <=  8'h00;      memory[49616] <=  8'h00;      memory[49617] <=  8'h00;      memory[49618] <=  8'h00;      memory[49619] <=  8'h00;      memory[49620] <=  8'h00;      memory[49621] <=  8'h00;      memory[49622] <=  8'h00;      memory[49623] <=  8'h00;      memory[49624] <=  8'h00;      memory[49625] <=  8'h00;      memory[49626] <=  8'h00;      memory[49627] <=  8'h00;      memory[49628] <=  8'h00;      memory[49629] <=  8'h00;      memory[49630] <=  8'h00;      memory[49631] <=  8'h00;      memory[49632] <=  8'h00;      memory[49633] <=  8'h00;      memory[49634] <=  8'h00;      memory[49635] <=  8'h00;      memory[49636] <=  8'h00;      memory[49637] <=  8'h00;      memory[49638] <=  8'h00;      memory[49639] <=  8'h00;      memory[49640] <=  8'h00;      memory[49641] <=  8'h00;      memory[49642] <=  8'h00;      memory[49643] <=  8'h00;      memory[49644] <=  8'h00;      memory[49645] <=  8'h00;      memory[49646] <=  8'h00;      memory[49647] <=  8'h00;      memory[49648] <=  8'h00;      memory[49649] <=  8'h00;      memory[49650] <=  8'h00;      memory[49651] <=  8'h00;      memory[49652] <=  8'h00;      memory[49653] <=  8'h00;      memory[49654] <=  8'h00;      memory[49655] <=  8'h00;      memory[49656] <=  8'h00;      memory[49657] <=  8'h00;      memory[49658] <=  8'h00;      memory[49659] <=  8'h00;      memory[49660] <=  8'h00;      memory[49661] <=  8'h00;      memory[49662] <=  8'h00;      memory[49663] <=  8'h00;      memory[49664] <=  8'h00;      memory[49665] <=  8'h00;      memory[49666] <=  8'h00;      memory[49667] <=  8'h00;      memory[49668] <=  8'h00;      memory[49669] <=  8'h00;      memory[49670] <=  8'h00;      memory[49671] <=  8'h00;      memory[49672] <=  8'h00;      memory[49673] <=  8'h00;      memory[49674] <=  8'h00;      memory[49675] <=  8'h00;      memory[49676] <=  8'h00;      memory[49677] <=  8'h00;      memory[49678] <=  8'h00;      memory[49679] <=  8'h00;      memory[49680] <=  8'h00;      memory[49681] <=  8'h00;      memory[49682] <=  8'h00;      memory[49683] <=  8'h00;      memory[49684] <=  8'h00;      memory[49685] <=  8'h00;      memory[49686] <=  8'h00;      memory[49687] <=  8'h00;      memory[49688] <=  8'h00;      memory[49689] <=  8'h00;      memory[49690] <=  8'h00;      memory[49691] <=  8'h00;      memory[49692] <=  8'h00;      memory[49693] <=  8'h00;      memory[49694] <=  8'h00;      memory[49695] <=  8'h00;      memory[49696] <=  8'h00;      memory[49697] <=  8'h00;      memory[49698] <=  8'h00;      memory[49699] <=  8'h00;      memory[49700] <=  8'h00;      memory[49701] <=  8'h00;      memory[49702] <=  8'h00;      memory[49703] <=  8'h00;      memory[49704] <=  8'h00;      memory[49705] <=  8'h00;      memory[49706] <=  8'h00;      memory[49707] <=  8'h00;      memory[49708] <=  8'h00;      memory[49709] <=  8'h00;      memory[49710] <=  8'h00;      memory[49711] <=  8'h00;      memory[49712] <=  8'h00;      memory[49713] <=  8'h00;      memory[49714] <=  8'h00;      memory[49715] <=  8'h00;      memory[49716] <=  8'h00;      memory[49717] <=  8'h00;      memory[49718] <=  8'h00;      memory[49719] <=  8'h00;      memory[49720] <=  8'h00;      memory[49721] <=  8'h00;      memory[49722] <=  8'h00;      memory[49723] <=  8'h00;      memory[49724] <=  8'h00;      memory[49725] <=  8'h00;      memory[49726] <=  8'h00;      memory[49727] <=  8'h00;      memory[49728] <=  8'h00;      memory[49729] <=  8'h00;      memory[49730] <=  8'h00;      memory[49731] <=  8'h00;      memory[49732] <=  8'h00;      memory[49733] <=  8'h00;      memory[49734] <=  8'h00;      memory[49735] <=  8'h00;      memory[49736] <=  8'h00;      memory[49737] <=  8'h00;      memory[49738] <=  8'h00;      memory[49739] <=  8'h00;      memory[49740] <=  8'h00;      memory[49741] <=  8'h00;      memory[49742] <=  8'h00;      memory[49743] <=  8'h00;      memory[49744] <=  8'h00;      memory[49745] <=  8'h00;      memory[49746] <=  8'h00;      memory[49747] <=  8'h00;      memory[49748] <=  8'h00;      memory[49749] <=  8'h00;      memory[49750] <=  8'h00;      memory[49751] <=  8'h00;      memory[49752] <=  8'h00;      memory[49753] <=  8'h00;      memory[49754] <=  8'h00;      memory[49755] <=  8'h00;      memory[49756] <=  8'h00;      memory[49757] <=  8'h00;      memory[49758] <=  8'h00;      memory[49759] <=  8'h00;      memory[49760] <=  8'h00;      memory[49761] <=  8'h00;      memory[49762] <=  8'h00;      memory[49763] <=  8'h00;      memory[49764] <=  8'h00;      memory[49765] <=  8'h00;      memory[49766] <=  8'h00;      memory[49767] <=  8'h00;      memory[49768] <=  8'h00;      memory[49769] <=  8'h00;      memory[49770] <=  8'h00;      memory[49771] <=  8'h00;      memory[49772] <=  8'h00;      memory[49773] <=  8'h00;      memory[49774] <=  8'h00;      memory[49775] <=  8'h00;      memory[49776] <=  8'h00;      memory[49777] <=  8'h00;      memory[49778] <=  8'h00;      memory[49779] <=  8'h00;      memory[49780] <=  8'h00;      memory[49781] <=  8'h00;      memory[49782] <=  8'h00;      memory[49783] <=  8'h00;      memory[49784] <=  8'h00;      memory[49785] <=  8'h00;      memory[49786] <=  8'h00;      memory[49787] <=  8'h00;      memory[49788] <=  8'h00;      memory[49789] <=  8'h00;      memory[49790] <=  8'h00;      memory[49791] <=  8'h00;      memory[49792] <=  8'h00;      memory[49793] <=  8'h00;      memory[49794] <=  8'h00;      memory[49795] <=  8'h00;      memory[49796] <=  8'h00;      memory[49797] <=  8'h00;      memory[49798] <=  8'h00;      memory[49799] <=  8'h00;      memory[49800] <=  8'h00;      memory[49801] <=  8'h00;      memory[49802] <=  8'h00;      memory[49803] <=  8'h00;      memory[49804] <=  8'h00;      memory[49805] <=  8'h00;      memory[49806] <=  8'h00;      memory[49807] <=  8'h00;      memory[49808] <=  8'h00;      memory[49809] <=  8'h00;      memory[49810] <=  8'h00;      memory[49811] <=  8'h00;      memory[49812] <=  8'h00;      memory[49813] <=  8'h00;      memory[49814] <=  8'h00;      memory[49815] <=  8'h00;      memory[49816] <=  8'h00;      memory[49817] <=  8'h00;      memory[49818] <=  8'h00;      memory[49819] <=  8'h00;      memory[49820] <=  8'h00;      memory[49821] <=  8'h00;      memory[49822] <=  8'h00;      memory[49823] <=  8'h00;      memory[49824] <=  8'h00;      memory[49825] <=  8'h00;      memory[49826] <=  8'h00;      memory[49827] <=  8'h00;      memory[49828] <=  8'h00;      memory[49829] <=  8'h00;      memory[49830] <=  8'h00;      memory[49831] <=  8'h00;      memory[49832] <=  8'h00;      memory[49833] <=  8'h00;      memory[49834] <=  8'h00;      memory[49835] <=  8'h00;      memory[49836] <=  8'h00;      memory[49837] <=  8'h00;      memory[49838] <=  8'h00;      memory[49839] <=  8'h00;      memory[49840] <=  8'h00;      memory[49841] <=  8'h00;      memory[49842] <=  8'h00;      memory[49843] <=  8'h00;      memory[49844] <=  8'h00;      memory[49845] <=  8'h00;      memory[49846] <=  8'h00;      memory[49847] <=  8'h00;      memory[49848] <=  8'h00;      memory[49849] <=  8'h00;      memory[49850] <=  8'h00;      memory[49851] <=  8'h00;      memory[49852] <=  8'h00;      memory[49853] <=  8'h00;      memory[49854] <=  8'h00;      memory[49855] <=  8'h00;      memory[49856] <=  8'h00;      memory[49857] <=  8'h00;      memory[49858] <=  8'h00;      memory[49859] <=  8'h00;      memory[49860] <=  8'h00;      memory[49861] <=  8'h00;      memory[49862] <=  8'h00;      memory[49863] <=  8'h00;      memory[49864] <=  8'h00;      memory[49865] <=  8'h00;      memory[49866] <=  8'h00;      memory[49867] <=  8'h00;      memory[49868] <=  8'h00;      memory[49869] <=  8'h00;      memory[49870] <=  8'h00;      memory[49871] <=  8'h00;      memory[49872] <=  8'h00;      memory[49873] <=  8'h00;      memory[49874] <=  8'h00;      memory[49875] <=  8'h00;      memory[49876] <=  8'h00;      memory[49877] <=  8'h00;      memory[49878] <=  8'h00;      memory[49879] <=  8'h00;      memory[49880] <=  8'h00;      memory[49881] <=  8'h00;      memory[49882] <=  8'h00;      memory[49883] <=  8'h00;      memory[49884] <=  8'h00;      memory[49885] <=  8'h00;      memory[49886] <=  8'h00;      memory[49887] <=  8'h00;      memory[49888] <=  8'h00;      memory[49889] <=  8'h00;      memory[49890] <=  8'h00;      memory[49891] <=  8'h00;      memory[49892] <=  8'h00;      memory[49893] <=  8'h00;      memory[49894] <=  8'h00;      memory[49895] <=  8'h00;      memory[49896] <=  8'h00;      memory[49897] <=  8'h00;      memory[49898] <=  8'h00;      memory[49899] <=  8'h00;      memory[49900] <=  8'h00;      memory[49901] <=  8'h00;      memory[49902] <=  8'h00;      memory[49903] <=  8'h00;      memory[49904] <=  8'h00;      memory[49905] <=  8'h00;      memory[49906] <=  8'h00;      memory[49907] <=  8'h00;      memory[49908] <=  8'h00;      memory[49909] <=  8'h00;      memory[49910] <=  8'h00;      memory[49911] <=  8'h00;      memory[49912] <=  8'h00;      memory[49913] <=  8'h00;      memory[49914] <=  8'h00;      memory[49915] <=  8'h00;      memory[49916] <=  8'h00;      memory[49917] <=  8'h00;      memory[49918] <=  8'h00;      memory[49919] <=  8'h00;      memory[49920] <=  8'h00;      memory[49921] <=  8'h00;      memory[49922] <=  8'h00;      memory[49923] <=  8'h00;      memory[49924] <=  8'h00;      memory[49925] <=  8'h00;      memory[49926] <=  8'h00;      memory[49927] <=  8'h00;      memory[49928] <=  8'h00;      memory[49929] <=  8'h00;      memory[49930] <=  8'h00;      memory[49931] <=  8'h00;      memory[49932] <=  8'h00;      memory[49933] <=  8'h00;      memory[49934] <=  8'h00;      memory[49935] <=  8'h00;      memory[49936] <=  8'h00;      memory[49937] <=  8'h00;      memory[49938] <=  8'h00;      memory[49939] <=  8'h00;      memory[49940] <=  8'h00;      memory[49941] <=  8'h00;      memory[49942] <=  8'h00;      memory[49943] <=  8'h00;      memory[49944] <=  8'h00;      memory[49945] <=  8'h00;      memory[49946] <=  8'h00;      memory[49947] <=  8'h00;      memory[49948] <=  8'h00;      memory[49949] <=  8'h00;      memory[49950] <=  8'h00;      memory[49951] <=  8'h00;      memory[49952] <=  8'h00;      memory[49953] <=  8'h00;      memory[49954] <=  8'h00;      memory[49955] <=  8'h00;      memory[49956] <=  8'h00;      memory[49957] <=  8'h00;      memory[49958] <=  8'h00;      memory[49959] <=  8'h00;      memory[49960] <=  8'h00;      memory[49961] <=  8'h00;      memory[49962] <=  8'h00;      memory[49963] <=  8'h00;      memory[49964] <=  8'h00;      memory[49965] <=  8'h00;      memory[49966] <=  8'h00;      memory[49967] <=  8'h00;      memory[49968] <=  8'h00;      memory[49969] <=  8'h00;      memory[49970] <=  8'h00;      memory[49971] <=  8'h00;      memory[49972] <=  8'h00;      memory[49973] <=  8'h00;      memory[49974] <=  8'h00;      memory[49975] <=  8'h00;      memory[49976] <=  8'h00;      memory[49977] <=  8'h00;      memory[49978] <=  8'h00;      memory[49979] <=  8'h00;      memory[49980] <=  8'h00;      memory[49981] <=  8'h00;      memory[49982] <=  8'h00;      memory[49983] <=  8'h00;      memory[49984] <=  8'h00;      memory[49985] <=  8'h00;      memory[49986] <=  8'h00;      memory[49987] <=  8'h00;      memory[49988] <=  8'h00;      memory[49989] <=  8'h00;      memory[49990] <=  8'h00;      memory[49991] <=  8'h00;      memory[49992] <=  8'h00;      memory[49993] <=  8'h00;      memory[49994] <=  8'h00;      memory[49995] <=  8'h00;      memory[49996] <=  8'h00;      memory[49997] <=  8'h00;      memory[49998] <=  8'h00;      memory[49999] <=  8'h00;      memory[50000] <=  8'h00;      memory[50001] <=  8'h00;      memory[50002] <=  8'h00;      memory[50003] <=  8'h00;      memory[50004] <=  8'h00;      memory[50005] <=  8'h00;      memory[50006] <=  8'h00;      memory[50007] <=  8'h00;      memory[50008] <=  8'h00;      memory[50009] <=  8'h00;      memory[50010] <=  8'h00;      memory[50011] <=  8'h00;      memory[50012] <=  8'h00;      memory[50013] <=  8'h00;      memory[50014] <=  8'h00;      memory[50015] <=  8'h00;      memory[50016] <=  8'h00;      memory[50017] <=  8'h00;      memory[50018] <=  8'h00;      memory[50019] <=  8'h00;      memory[50020] <=  8'h00;      memory[50021] <=  8'h00;      memory[50022] <=  8'h00;      memory[50023] <=  8'h00;      memory[50024] <=  8'h00;      memory[50025] <=  8'h00;      memory[50026] <=  8'h00;      memory[50027] <=  8'h00;      memory[50028] <=  8'h00;      memory[50029] <=  8'h00;      memory[50030] <=  8'h00;      memory[50031] <=  8'h00;      memory[50032] <=  8'h00;      memory[50033] <=  8'h00;      memory[50034] <=  8'h00;      memory[50035] <=  8'h00;      memory[50036] <=  8'h00;      memory[50037] <=  8'h00;      memory[50038] <=  8'h00;      memory[50039] <=  8'h00;      memory[50040] <=  8'h00;      memory[50041] <=  8'h00;      memory[50042] <=  8'h00;      memory[50043] <=  8'h00;      memory[50044] <=  8'h00;      memory[50045] <=  8'h00;      memory[50046] <=  8'h00;      memory[50047] <=  8'h00;      memory[50048] <=  8'h00;      memory[50049] <=  8'h00;      memory[50050] <=  8'h00;      memory[50051] <=  8'h00;      memory[50052] <=  8'h00;      memory[50053] <=  8'h00;      memory[50054] <=  8'h00;      memory[50055] <=  8'h00;      memory[50056] <=  8'h00;      memory[50057] <=  8'h00;      memory[50058] <=  8'h00;      memory[50059] <=  8'h00;      memory[50060] <=  8'h00;      memory[50061] <=  8'h00;      memory[50062] <=  8'h00;      memory[50063] <=  8'h00;      memory[50064] <=  8'h00;      memory[50065] <=  8'h00;      memory[50066] <=  8'h00;      memory[50067] <=  8'h00;      memory[50068] <=  8'h00;      memory[50069] <=  8'h00;      memory[50070] <=  8'h00;      memory[50071] <=  8'h00;      memory[50072] <=  8'h00;      memory[50073] <=  8'h00;      memory[50074] <=  8'h00;      memory[50075] <=  8'h00;      memory[50076] <=  8'h00;      memory[50077] <=  8'h00;      memory[50078] <=  8'h00;      memory[50079] <=  8'h00;      memory[50080] <=  8'h00;      memory[50081] <=  8'h00;      memory[50082] <=  8'h00;      memory[50083] <=  8'h00;      memory[50084] <=  8'h00;      memory[50085] <=  8'h00;      memory[50086] <=  8'h00;      memory[50087] <=  8'h00;      memory[50088] <=  8'h00;      memory[50089] <=  8'h00;      memory[50090] <=  8'h00;      memory[50091] <=  8'h00;      memory[50092] <=  8'h00;      memory[50093] <=  8'h00;      memory[50094] <=  8'h00;      memory[50095] <=  8'h00;      memory[50096] <=  8'h00;      memory[50097] <=  8'h00;      memory[50098] <=  8'h00;      memory[50099] <=  8'h00;      memory[50100] <=  8'h00;      memory[50101] <=  8'h00;      memory[50102] <=  8'h00;      memory[50103] <=  8'h00;      memory[50104] <=  8'h00;      memory[50105] <=  8'h00;      memory[50106] <=  8'h00;      memory[50107] <=  8'h00;      memory[50108] <=  8'h00;      memory[50109] <=  8'h00;      memory[50110] <=  8'h00;      memory[50111] <=  8'h00;      memory[50112] <=  8'h00;      memory[50113] <=  8'h00;      memory[50114] <=  8'h00;      memory[50115] <=  8'h00;      memory[50116] <=  8'h00;      memory[50117] <=  8'h00;      memory[50118] <=  8'h00;      memory[50119] <=  8'h00;      memory[50120] <=  8'h00;      memory[50121] <=  8'h00;      memory[50122] <=  8'h00;      memory[50123] <=  8'h00;      memory[50124] <=  8'h00;      memory[50125] <=  8'h00;      memory[50126] <=  8'h00;      memory[50127] <=  8'h00;      memory[50128] <=  8'h00;      memory[50129] <=  8'h00;      memory[50130] <=  8'h00;      memory[50131] <=  8'h00;      memory[50132] <=  8'h00;      memory[50133] <=  8'h00;      memory[50134] <=  8'h00;      memory[50135] <=  8'h00;      memory[50136] <=  8'h00;      memory[50137] <=  8'h00;      memory[50138] <=  8'h00;      memory[50139] <=  8'h00;      memory[50140] <=  8'h00;      memory[50141] <=  8'h00;      memory[50142] <=  8'h00;      memory[50143] <=  8'h00;      memory[50144] <=  8'h00;      memory[50145] <=  8'h00;      memory[50146] <=  8'h00;      memory[50147] <=  8'h00;      memory[50148] <=  8'h00;      memory[50149] <=  8'h00;      memory[50150] <=  8'h00;      memory[50151] <=  8'h00;      memory[50152] <=  8'h00;      memory[50153] <=  8'h00;      memory[50154] <=  8'h00;      memory[50155] <=  8'h00;      memory[50156] <=  8'h00;      memory[50157] <=  8'h00;      memory[50158] <=  8'h00;      memory[50159] <=  8'h00;      memory[50160] <=  8'h00;      memory[50161] <=  8'h00;      memory[50162] <=  8'h00;      memory[50163] <=  8'h00;      memory[50164] <=  8'h00;      memory[50165] <=  8'h00;      memory[50166] <=  8'h00;      memory[50167] <=  8'h00;      memory[50168] <=  8'h00;      memory[50169] <=  8'h00;      memory[50170] <=  8'h00;      memory[50171] <=  8'h00;      memory[50172] <=  8'h00;      memory[50173] <=  8'h00;      memory[50174] <=  8'h00;      memory[50175] <=  8'h00;      memory[50176] <=  8'h00;      memory[50177] <=  8'h00;      memory[50178] <=  8'h00;      memory[50179] <=  8'h00;      memory[50180] <=  8'h00;      memory[50181] <=  8'h00;      memory[50182] <=  8'h00;      memory[50183] <=  8'h00;      memory[50184] <=  8'h00;      memory[50185] <=  8'h00;      memory[50186] <=  8'h00;      memory[50187] <=  8'h00;      memory[50188] <=  8'h00;      memory[50189] <=  8'h00;      memory[50190] <=  8'h00;      memory[50191] <=  8'h00;      memory[50192] <=  8'h00;      memory[50193] <=  8'h00;      memory[50194] <=  8'h00;      memory[50195] <=  8'h00;      memory[50196] <=  8'h00;      memory[50197] <=  8'h00;      memory[50198] <=  8'h00;      memory[50199] <=  8'h00;      memory[50200] <=  8'h00;      memory[50201] <=  8'h00;      memory[50202] <=  8'h00;      memory[50203] <=  8'h00;      memory[50204] <=  8'h00;      memory[50205] <=  8'h00;      memory[50206] <=  8'h00;      memory[50207] <=  8'h00;      memory[50208] <=  8'h00;      memory[50209] <=  8'h00;      memory[50210] <=  8'h00;      memory[50211] <=  8'h00;      memory[50212] <=  8'h00;      memory[50213] <=  8'h00;      memory[50214] <=  8'h00;      memory[50215] <=  8'h00;      memory[50216] <=  8'h00;      memory[50217] <=  8'h00;      memory[50218] <=  8'h00;      memory[50219] <=  8'h00;      memory[50220] <=  8'h00;      memory[50221] <=  8'h00;      memory[50222] <=  8'h00;      memory[50223] <=  8'h00;      memory[50224] <=  8'h00;      memory[50225] <=  8'h00;      memory[50226] <=  8'h00;      memory[50227] <=  8'h00;      memory[50228] <=  8'h00;      memory[50229] <=  8'h00;      memory[50230] <=  8'h00;      memory[50231] <=  8'h00;      memory[50232] <=  8'h00;      memory[50233] <=  8'h00;      memory[50234] <=  8'h00;      memory[50235] <=  8'h00;      memory[50236] <=  8'h00;      memory[50237] <=  8'h00;      memory[50238] <=  8'h00;      memory[50239] <=  8'h00;      memory[50240] <=  8'h00;      memory[50241] <=  8'h00;      memory[50242] <=  8'h00;      memory[50243] <=  8'h00;      memory[50244] <=  8'h00;      memory[50245] <=  8'h00;      memory[50246] <=  8'h00;      memory[50247] <=  8'h00;      memory[50248] <=  8'h00;      memory[50249] <=  8'h00;      memory[50250] <=  8'h00;      memory[50251] <=  8'h00;      memory[50252] <=  8'h00;      memory[50253] <=  8'h00;      memory[50254] <=  8'h00;      memory[50255] <=  8'h00;      memory[50256] <=  8'h00;      memory[50257] <=  8'h00;      memory[50258] <=  8'h00;      memory[50259] <=  8'h00;      memory[50260] <=  8'h00;      memory[50261] <=  8'h00;      memory[50262] <=  8'h00;      memory[50263] <=  8'h00;      memory[50264] <=  8'h00;      memory[50265] <=  8'h00;      memory[50266] <=  8'h00;      memory[50267] <=  8'h00;      memory[50268] <=  8'h00;      memory[50269] <=  8'h00;      memory[50270] <=  8'h00;      memory[50271] <=  8'h00;      memory[50272] <=  8'h00;      memory[50273] <=  8'h00;      memory[50274] <=  8'h00;      memory[50275] <=  8'h00;      memory[50276] <=  8'h00;      memory[50277] <=  8'h00;      memory[50278] <=  8'h00;      memory[50279] <=  8'h00;      memory[50280] <=  8'h00;      memory[50281] <=  8'h00;      memory[50282] <=  8'h00;      memory[50283] <=  8'h00;      memory[50284] <=  8'h00;      memory[50285] <=  8'h00;      memory[50286] <=  8'h00;      memory[50287] <=  8'h00;      memory[50288] <=  8'h00;      memory[50289] <=  8'h00;      memory[50290] <=  8'h00;      memory[50291] <=  8'h00;      memory[50292] <=  8'h00;      memory[50293] <=  8'h00;      memory[50294] <=  8'h00;      memory[50295] <=  8'h00;      memory[50296] <=  8'h00;      memory[50297] <=  8'h00;      memory[50298] <=  8'h00;      memory[50299] <=  8'h00;      memory[50300] <=  8'h00;      memory[50301] <=  8'h00;      memory[50302] <=  8'h00;      memory[50303] <=  8'h00;      memory[50304] <=  8'h00;      memory[50305] <=  8'h00;      memory[50306] <=  8'h00;      memory[50307] <=  8'h00;      memory[50308] <=  8'h00;      memory[50309] <=  8'h00;      memory[50310] <=  8'h00;      memory[50311] <=  8'h00;      memory[50312] <=  8'h00;      memory[50313] <=  8'h00;      memory[50314] <=  8'h00;      memory[50315] <=  8'h00;      memory[50316] <=  8'h00;      memory[50317] <=  8'h00;      memory[50318] <=  8'h00;      memory[50319] <=  8'h00;      memory[50320] <=  8'h00;      memory[50321] <=  8'h00;      memory[50322] <=  8'h00;      memory[50323] <=  8'h00;      memory[50324] <=  8'h00;      memory[50325] <=  8'h00;      memory[50326] <=  8'h00;      memory[50327] <=  8'h00;      memory[50328] <=  8'h00;      memory[50329] <=  8'h00;      memory[50330] <=  8'h00;      memory[50331] <=  8'h00;      memory[50332] <=  8'h00;      memory[50333] <=  8'h00;      memory[50334] <=  8'h00;      memory[50335] <=  8'h00;      memory[50336] <=  8'h00;      memory[50337] <=  8'h00;      memory[50338] <=  8'h00;      memory[50339] <=  8'h00;      memory[50340] <=  8'h00;      memory[50341] <=  8'h00;      memory[50342] <=  8'h00;      memory[50343] <=  8'h00;      memory[50344] <=  8'h00;      memory[50345] <=  8'h00;      memory[50346] <=  8'h00;      memory[50347] <=  8'h00;      memory[50348] <=  8'h00;      memory[50349] <=  8'h00;      memory[50350] <=  8'h00;      memory[50351] <=  8'h00;      memory[50352] <=  8'h00;      memory[50353] <=  8'h00;      memory[50354] <=  8'h00;      memory[50355] <=  8'h00;      memory[50356] <=  8'h00;      memory[50357] <=  8'h00;      memory[50358] <=  8'h00;      memory[50359] <=  8'h00;      memory[50360] <=  8'h00;      memory[50361] <=  8'h00;      memory[50362] <=  8'h00;      memory[50363] <=  8'h00;      memory[50364] <=  8'h00;      memory[50365] <=  8'h00;      memory[50366] <=  8'h00;      memory[50367] <=  8'h00;      memory[50368] <=  8'h00;      memory[50369] <=  8'h00;      memory[50370] <=  8'h00;      memory[50371] <=  8'h00;      memory[50372] <=  8'h00;      memory[50373] <=  8'h00;      memory[50374] <=  8'h00;      memory[50375] <=  8'h00;      memory[50376] <=  8'h00;      memory[50377] <=  8'h00;      memory[50378] <=  8'h00;      memory[50379] <=  8'h00;      memory[50380] <=  8'h00;      memory[50381] <=  8'h00;      memory[50382] <=  8'h00;      memory[50383] <=  8'h00;      memory[50384] <=  8'h00;      memory[50385] <=  8'h00;      memory[50386] <=  8'h00;      memory[50387] <=  8'h00;      memory[50388] <=  8'h00;      memory[50389] <=  8'h00;      memory[50390] <=  8'h00;      memory[50391] <=  8'h00;      memory[50392] <=  8'h00;      memory[50393] <=  8'h00;      memory[50394] <=  8'h00;      memory[50395] <=  8'h00;      memory[50396] <=  8'h00;      memory[50397] <=  8'h00;      memory[50398] <=  8'h00;      memory[50399] <=  8'h00;      memory[50400] <=  8'h00;      memory[50401] <=  8'h00;      memory[50402] <=  8'h00;      memory[50403] <=  8'h00;      memory[50404] <=  8'h00;      memory[50405] <=  8'h00;      memory[50406] <=  8'h00;      memory[50407] <=  8'h00;      memory[50408] <=  8'h00;      memory[50409] <=  8'h00;      memory[50410] <=  8'h00;      memory[50411] <=  8'h00;      memory[50412] <=  8'h00;      memory[50413] <=  8'h00;      memory[50414] <=  8'h00;      memory[50415] <=  8'h00;      memory[50416] <=  8'h00;      memory[50417] <=  8'h00;      memory[50418] <=  8'h00;      memory[50419] <=  8'h00;      memory[50420] <=  8'h00;      memory[50421] <=  8'h00;      memory[50422] <=  8'h00;      memory[50423] <=  8'h00;      memory[50424] <=  8'h00;      memory[50425] <=  8'h00;      memory[50426] <=  8'h00;      memory[50427] <=  8'h00;      memory[50428] <=  8'h00;      memory[50429] <=  8'h00;      memory[50430] <=  8'h00;      memory[50431] <=  8'h00;      memory[50432] <=  8'h00;      memory[50433] <=  8'h00;      memory[50434] <=  8'h00;      memory[50435] <=  8'h00;      memory[50436] <=  8'h00;      memory[50437] <=  8'h00;      memory[50438] <=  8'h00;      memory[50439] <=  8'h00;      memory[50440] <=  8'h00;      memory[50441] <=  8'h00;      memory[50442] <=  8'h00;      memory[50443] <=  8'h00;      memory[50444] <=  8'h00;      memory[50445] <=  8'h00;      memory[50446] <=  8'h00;      memory[50447] <=  8'h00;      memory[50448] <=  8'h00;      memory[50449] <=  8'h00;      memory[50450] <=  8'h00;      memory[50451] <=  8'h00;      memory[50452] <=  8'h00;      memory[50453] <=  8'h00;      memory[50454] <=  8'h00;      memory[50455] <=  8'h00;      memory[50456] <=  8'h00;      memory[50457] <=  8'h00;      memory[50458] <=  8'h00;      memory[50459] <=  8'h00;      memory[50460] <=  8'h00;      memory[50461] <=  8'h00;      memory[50462] <=  8'h00;      memory[50463] <=  8'h00;      memory[50464] <=  8'h00;      memory[50465] <=  8'h00;      memory[50466] <=  8'h00;      memory[50467] <=  8'h00;      memory[50468] <=  8'h00;      memory[50469] <=  8'h00;      memory[50470] <=  8'h00;      memory[50471] <=  8'h00;      memory[50472] <=  8'h00;      memory[50473] <=  8'h00;      memory[50474] <=  8'h00;      memory[50475] <=  8'h00;      memory[50476] <=  8'h00;      memory[50477] <=  8'h00;      memory[50478] <=  8'h00;      memory[50479] <=  8'h00;      memory[50480] <=  8'h00;      memory[50481] <=  8'h00;      memory[50482] <=  8'h00;      memory[50483] <=  8'h00;      memory[50484] <=  8'h00;      memory[50485] <=  8'h00;      memory[50486] <=  8'h00;      memory[50487] <=  8'h00;      memory[50488] <=  8'h00;      memory[50489] <=  8'h00;      memory[50490] <=  8'h00;      memory[50491] <=  8'h00;      memory[50492] <=  8'h00;      memory[50493] <=  8'h00;      memory[50494] <=  8'h00;      memory[50495] <=  8'h00;      memory[50496] <=  8'h00;      memory[50497] <=  8'h00;      memory[50498] <=  8'h00;      memory[50499] <=  8'h00;      memory[50500] <=  8'h00;      memory[50501] <=  8'h00;      memory[50502] <=  8'h00;      memory[50503] <=  8'h00;      memory[50504] <=  8'h00;      memory[50505] <=  8'h00;      memory[50506] <=  8'h00;      memory[50507] <=  8'h00;      memory[50508] <=  8'h00;      memory[50509] <=  8'h00;      memory[50510] <=  8'h00;      memory[50511] <=  8'h00;      memory[50512] <=  8'h00;      memory[50513] <=  8'h00;      memory[50514] <=  8'h00;      memory[50515] <=  8'h00;      memory[50516] <=  8'h00;      memory[50517] <=  8'h00;      memory[50518] <=  8'h00;      memory[50519] <=  8'h00;      memory[50520] <=  8'h00;      memory[50521] <=  8'h00;      memory[50522] <=  8'h00;      memory[50523] <=  8'h00;      memory[50524] <=  8'h00;      memory[50525] <=  8'h00;      memory[50526] <=  8'h00;      memory[50527] <=  8'h00;      memory[50528] <=  8'h00;      memory[50529] <=  8'h00;      memory[50530] <=  8'h00;      memory[50531] <=  8'h00;      memory[50532] <=  8'h00;      memory[50533] <=  8'h00;      memory[50534] <=  8'h00;      memory[50535] <=  8'h00;      memory[50536] <=  8'h00;      memory[50537] <=  8'h00;      memory[50538] <=  8'h00;      memory[50539] <=  8'h00;      memory[50540] <=  8'h00;      memory[50541] <=  8'h00;      memory[50542] <=  8'h00;      memory[50543] <=  8'h00;      memory[50544] <=  8'h00;      memory[50545] <=  8'h00;      memory[50546] <=  8'h00;      memory[50547] <=  8'h00;      memory[50548] <=  8'h00;      memory[50549] <=  8'h00;      memory[50550] <=  8'h00;      memory[50551] <=  8'h00;      memory[50552] <=  8'h00;      memory[50553] <=  8'h00;      memory[50554] <=  8'h00;      memory[50555] <=  8'h00;      memory[50556] <=  8'h00;      memory[50557] <=  8'h00;      memory[50558] <=  8'h00;      memory[50559] <=  8'h00;      memory[50560] <=  8'h00;      memory[50561] <=  8'h00;      memory[50562] <=  8'h00;      memory[50563] <=  8'h00;      memory[50564] <=  8'h00;      memory[50565] <=  8'h00;      memory[50566] <=  8'h00;      memory[50567] <=  8'h00;      memory[50568] <=  8'h00;      memory[50569] <=  8'h00;      memory[50570] <=  8'h00;      memory[50571] <=  8'h00;      memory[50572] <=  8'h00;      memory[50573] <=  8'h00;      memory[50574] <=  8'h00;      memory[50575] <=  8'h00;      memory[50576] <=  8'h00;      memory[50577] <=  8'h00;      memory[50578] <=  8'h00;      memory[50579] <=  8'h00;      memory[50580] <=  8'h00;      memory[50581] <=  8'h00;      memory[50582] <=  8'h00;      memory[50583] <=  8'h00;      memory[50584] <=  8'h00;      memory[50585] <=  8'h00;      memory[50586] <=  8'h00;      memory[50587] <=  8'h00;      memory[50588] <=  8'h00;      memory[50589] <=  8'h00;      memory[50590] <=  8'h00;      memory[50591] <=  8'h00;      memory[50592] <=  8'h00;      memory[50593] <=  8'h00;      memory[50594] <=  8'h00;      memory[50595] <=  8'h00;      memory[50596] <=  8'h00;      memory[50597] <=  8'h00;      memory[50598] <=  8'h00;      memory[50599] <=  8'h00;      memory[50600] <=  8'h00;      memory[50601] <=  8'h00;      memory[50602] <=  8'h00;      memory[50603] <=  8'h00;      memory[50604] <=  8'h00;      memory[50605] <=  8'h00;      memory[50606] <=  8'h00;      memory[50607] <=  8'h00;      memory[50608] <=  8'h00;      memory[50609] <=  8'h00;      memory[50610] <=  8'h00;      memory[50611] <=  8'h00;      memory[50612] <=  8'h00;      memory[50613] <=  8'h00;      memory[50614] <=  8'h00;      memory[50615] <=  8'h00;      memory[50616] <=  8'h00;      memory[50617] <=  8'h00;      memory[50618] <=  8'h00;      memory[50619] <=  8'h00;      memory[50620] <=  8'h00;      memory[50621] <=  8'h00;      memory[50622] <=  8'h00;      memory[50623] <=  8'h00;      memory[50624] <=  8'h00;      memory[50625] <=  8'h00;      memory[50626] <=  8'h00;      memory[50627] <=  8'h00;      memory[50628] <=  8'h00;      memory[50629] <=  8'h00;      memory[50630] <=  8'h00;      memory[50631] <=  8'h00;      memory[50632] <=  8'h00;      memory[50633] <=  8'h00;      memory[50634] <=  8'h00;      memory[50635] <=  8'h00;      memory[50636] <=  8'h00;      memory[50637] <=  8'h00;      memory[50638] <=  8'h00;      memory[50639] <=  8'h00;      memory[50640] <=  8'h00;      memory[50641] <=  8'h00;      memory[50642] <=  8'h00;      memory[50643] <=  8'h00;      memory[50644] <=  8'h00;      memory[50645] <=  8'h00;      memory[50646] <=  8'h00;      memory[50647] <=  8'h00;      memory[50648] <=  8'h00;      memory[50649] <=  8'h00;      memory[50650] <=  8'h00;      memory[50651] <=  8'h00;      memory[50652] <=  8'h00;      memory[50653] <=  8'h00;      memory[50654] <=  8'h00;      memory[50655] <=  8'h00;      memory[50656] <=  8'h00;      memory[50657] <=  8'h00;      memory[50658] <=  8'h00;      memory[50659] <=  8'h00;      memory[50660] <=  8'h00;      memory[50661] <=  8'h00;      memory[50662] <=  8'h00;      memory[50663] <=  8'h00;      memory[50664] <=  8'h00;      memory[50665] <=  8'h00;      memory[50666] <=  8'h00;      memory[50667] <=  8'h00;      memory[50668] <=  8'h00;      memory[50669] <=  8'h00;      memory[50670] <=  8'h00;      memory[50671] <=  8'h00;      memory[50672] <=  8'h00;      memory[50673] <=  8'h00;      memory[50674] <=  8'h00;      memory[50675] <=  8'h00;      memory[50676] <=  8'h00;      memory[50677] <=  8'h00;      memory[50678] <=  8'h00;      memory[50679] <=  8'h00;      memory[50680] <=  8'h00;      memory[50681] <=  8'h00;      memory[50682] <=  8'h00;      memory[50683] <=  8'h00;      memory[50684] <=  8'h00;      memory[50685] <=  8'h00;      memory[50686] <=  8'h00;      memory[50687] <=  8'h00;      memory[50688] <=  8'h00;      memory[50689] <=  8'h00;      memory[50690] <=  8'h00;      memory[50691] <=  8'h00;      memory[50692] <=  8'h00;      memory[50693] <=  8'h00;      memory[50694] <=  8'h00;      memory[50695] <=  8'h00;      memory[50696] <=  8'h00;      memory[50697] <=  8'h00;      memory[50698] <=  8'h00;      memory[50699] <=  8'h00;      memory[50700] <=  8'h00;      memory[50701] <=  8'h00;      memory[50702] <=  8'h00;      memory[50703] <=  8'h00;      memory[50704] <=  8'h00;      memory[50705] <=  8'h00;      memory[50706] <=  8'h00;      memory[50707] <=  8'h00;      memory[50708] <=  8'h00;      memory[50709] <=  8'h00;      memory[50710] <=  8'h00;      memory[50711] <=  8'h00;      memory[50712] <=  8'h00;      memory[50713] <=  8'h00;      memory[50714] <=  8'h00;      memory[50715] <=  8'h00;      memory[50716] <=  8'h00;      memory[50717] <=  8'h00;      memory[50718] <=  8'h00;      memory[50719] <=  8'h00;      memory[50720] <=  8'h00;      memory[50721] <=  8'h00;      memory[50722] <=  8'h00;      memory[50723] <=  8'h00;      memory[50724] <=  8'h00;      memory[50725] <=  8'h00;      memory[50726] <=  8'h00;      memory[50727] <=  8'h00;      memory[50728] <=  8'h00;      memory[50729] <=  8'h00;      memory[50730] <=  8'h00;      memory[50731] <=  8'h00;      memory[50732] <=  8'h00;      memory[50733] <=  8'h00;      memory[50734] <=  8'h00;      memory[50735] <=  8'h00;      memory[50736] <=  8'h00;      memory[50737] <=  8'h00;      memory[50738] <=  8'h00;      memory[50739] <=  8'h00;      memory[50740] <=  8'h00;      memory[50741] <=  8'h00;      memory[50742] <=  8'h00;      memory[50743] <=  8'h00;      memory[50744] <=  8'h00;      memory[50745] <=  8'h00;      memory[50746] <=  8'h00;      memory[50747] <=  8'h00;      memory[50748] <=  8'h00;      memory[50749] <=  8'h00;      memory[50750] <=  8'h00;      memory[50751] <=  8'h00;      memory[50752] <=  8'h00;      memory[50753] <=  8'h00;      memory[50754] <=  8'h00;      memory[50755] <=  8'h00;      memory[50756] <=  8'h00;      memory[50757] <=  8'h00;      memory[50758] <=  8'h00;      memory[50759] <=  8'h00;      memory[50760] <=  8'h00;      memory[50761] <=  8'h00;      memory[50762] <=  8'h00;      memory[50763] <=  8'h00;      memory[50764] <=  8'h00;      memory[50765] <=  8'h00;      memory[50766] <=  8'h00;      memory[50767] <=  8'h00;      memory[50768] <=  8'h00;      memory[50769] <=  8'h00;      memory[50770] <=  8'h00;      memory[50771] <=  8'h00;      memory[50772] <=  8'h00;      memory[50773] <=  8'h00;      memory[50774] <=  8'h00;      memory[50775] <=  8'h00;      memory[50776] <=  8'h00;      memory[50777] <=  8'h00;      memory[50778] <=  8'h00;      memory[50779] <=  8'h00;      memory[50780] <=  8'h00;      memory[50781] <=  8'h00;      memory[50782] <=  8'h00;      memory[50783] <=  8'h00;      memory[50784] <=  8'h00;      memory[50785] <=  8'h00;      memory[50786] <=  8'h00;      memory[50787] <=  8'h00;      memory[50788] <=  8'h00;      memory[50789] <=  8'h00;      memory[50790] <=  8'h00;      memory[50791] <=  8'h00;      memory[50792] <=  8'h00;      memory[50793] <=  8'h00;      memory[50794] <=  8'h00;      memory[50795] <=  8'h00;      memory[50796] <=  8'h00;      memory[50797] <=  8'h00;      memory[50798] <=  8'h00;      memory[50799] <=  8'h00;      memory[50800] <=  8'h00;      memory[50801] <=  8'h00;      memory[50802] <=  8'h00;      memory[50803] <=  8'h00;      memory[50804] <=  8'h00;      memory[50805] <=  8'h00;      memory[50806] <=  8'h00;      memory[50807] <=  8'h00;      memory[50808] <=  8'h00;      memory[50809] <=  8'h00;      memory[50810] <=  8'h00;      memory[50811] <=  8'h00;      memory[50812] <=  8'h00;      memory[50813] <=  8'h00;      memory[50814] <=  8'h00;      memory[50815] <=  8'h00;      memory[50816] <=  8'h00;      memory[50817] <=  8'h00;      memory[50818] <=  8'h00;      memory[50819] <=  8'h00;      memory[50820] <=  8'h00;      memory[50821] <=  8'h00;      memory[50822] <=  8'h00;      memory[50823] <=  8'h00;      memory[50824] <=  8'h00;      memory[50825] <=  8'h00;      memory[50826] <=  8'h00;      memory[50827] <=  8'h00;      memory[50828] <=  8'h00;      memory[50829] <=  8'h00;      memory[50830] <=  8'h00;      memory[50831] <=  8'h00;      memory[50832] <=  8'h00;      memory[50833] <=  8'h00;      memory[50834] <=  8'h00;      memory[50835] <=  8'h00;      memory[50836] <=  8'h00;      memory[50837] <=  8'h00;      memory[50838] <=  8'h00;      memory[50839] <=  8'h00;      memory[50840] <=  8'h00;      memory[50841] <=  8'h00;      memory[50842] <=  8'h00;      memory[50843] <=  8'h00;      memory[50844] <=  8'h00;      memory[50845] <=  8'h00;      memory[50846] <=  8'h00;      memory[50847] <=  8'h00;      memory[50848] <=  8'h00;      memory[50849] <=  8'h00;      memory[50850] <=  8'h00;      memory[50851] <=  8'h00;      memory[50852] <=  8'h00;      memory[50853] <=  8'h00;      memory[50854] <=  8'h00;      memory[50855] <=  8'h00;      memory[50856] <=  8'h00;      memory[50857] <=  8'h00;      memory[50858] <=  8'h00;      memory[50859] <=  8'h00;      memory[50860] <=  8'h00;      memory[50861] <=  8'h00;      memory[50862] <=  8'h00;      memory[50863] <=  8'h00;      memory[50864] <=  8'h00;      memory[50865] <=  8'h00;      memory[50866] <=  8'h00;      memory[50867] <=  8'h00;      memory[50868] <=  8'h00;      memory[50869] <=  8'h00;      memory[50870] <=  8'h00;      memory[50871] <=  8'h00;      memory[50872] <=  8'h00;      memory[50873] <=  8'h00;      memory[50874] <=  8'h00;      memory[50875] <=  8'h00;      memory[50876] <=  8'h00;      memory[50877] <=  8'h00;      memory[50878] <=  8'h00;      memory[50879] <=  8'h00;      memory[50880] <=  8'h00;      memory[50881] <=  8'h00;      memory[50882] <=  8'h00;      memory[50883] <=  8'h00;      memory[50884] <=  8'h00;      memory[50885] <=  8'h00;      memory[50886] <=  8'h00;      memory[50887] <=  8'h00;      memory[50888] <=  8'h00;      memory[50889] <=  8'h00;      memory[50890] <=  8'h00;      memory[50891] <=  8'h00;      memory[50892] <=  8'h00;      memory[50893] <=  8'h00;      memory[50894] <=  8'h00;      memory[50895] <=  8'h00;      memory[50896] <=  8'h00;      memory[50897] <=  8'h00;      memory[50898] <=  8'h00;      memory[50899] <=  8'h00;      memory[50900] <=  8'h00;      memory[50901] <=  8'h00;      memory[50902] <=  8'h00;      memory[50903] <=  8'h00;      memory[50904] <=  8'h00;      memory[50905] <=  8'h00;      memory[50906] <=  8'h00;      memory[50907] <=  8'h00;      memory[50908] <=  8'h00;      memory[50909] <=  8'h00;      memory[50910] <=  8'h00;      memory[50911] <=  8'h00;      memory[50912] <=  8'h00;      memory[50913] <=  8'h00;      memory[50914] <=  8'h00;      memory[50915] <=  8'h00;      memory[50916] <=  8'h00;      memory[50917] <=  8'h00;      memory[50918] <=  8'h00;      memory[50919] <=  8'h00;      memory[50920] <=  8'h00;      memory[50921] <=  8'h00;      memory[50922] <=  8'h00;      memory[50923] <=  8'h00;      memory[50924] <=  8'h00;      memory[50925] <=  8'h00;      memory[50926] <=  8'h00;      memory[50927] <=  8'h00;      memory[50928] <=  8'h00;      memory[50929] <=  8'h00;      memory[50930] <=  8'h00;      memory[50931] <=  8'h00;      memory[50932] <=  8'h00;      memory[50933] <=  8'h00;      memory[50934] <=  8'h00;      memory[50935] <=  8'h00;      memory[50936] <=  8'h00;      memory[50937] <=  8'h00;      memory[50938] <=  8'h00;      memory[50939] <=  8'h00;      memory[50940] <=  8'h00;      memory[50941] <=  8'h00;      memory[50942] <=  8'h00;      memory[50943] <=  8'h00;      memory[50944] <=  8'h00;      memory[50945] <=  8'h00;      memory[50946] <=  8'h00;      memory[50947] <=  8'h00;      memory[50948] <=  8'h00;      memory[50949] <=  8'h00;      memory[50950] <=  8'h00;      memory[50951] <=  8'h00;      memory[50952] <=  8'h00;      memory[50953] <=  8'h00;      memory[50954] <=  8'h00;      memory[50955] <=  8'h00;      memory[50956] <=  8'h00;      memory[50957] <=  8'h00;      memory[50958] <=  8'h00;      memory[50959] <=  8'h00;      memory[50960] <=  8'h00;      memory[50961] <=  8'h00;      memory[50962] <=  8'h00;      memory[50963] <=  8'h00;      memory[50964] <=  8'h00;      memory[50965] <=  8'h00;      memory[50966] <=  8'h00;      memory[50967] <=  8'h00;      memory[50968] <=  8'h00;      memory[50969] <=  8'h00;      memory[50970] <=  8'h00;      memory[50971] <=  8'h00;      memory[50972] <=  8'h00;      memory[50973] <=  8'h00;      memory[50974] <=  8'h00;      memory[50975] <=  8'h00;      memory[50976] <=  8'h00;      memory[50977] <=  8'h00;      memory[50978] <=  8'h00;      memory[50979] <=  8'h00;      memory[50980] <=  8'h00;      memory[50981] <=  8'h00;      memory[50982] <=  8'h00;      memory[50983] <=  8'h00;      memory[50984] <=  8'h00;      memory[50985] <=  8'h00;      memory[50986] <=  8'h00;      memory[50987] <=  8'h00;      memory[50988] <=  8'h00;      memory[50989] <=  8'h00;      memory[50990] <=  8'h00;      memory[50991] <=  8'h00;      memory[50992] <=  8'h00;      memory[50993] <=  8'h00;      memory[50994] <=  8'h00;      memory[50995] <=  8'h00;      memory[50996] <=  8'h00;      memory[50997] <=  8'h00;      memory[50998] <=  8'h00;      memory[50999] <=  8'h00;      memory[51000] <=  8'h00;      memory[51001] <=  8'h00;      memory[51002] <=  8'h00;      memory[51003] <=  8'h00;      memory[51004] <=  8'h00;      memory[51005] <=  8'h00;      memory[51006] <=  8'h00;      memory[51007] <=  8'h00;      memory[51008] <=  8'h00;      memory[51009] <=  8'h00;      memory[51010] <=  8'h00;      memory[51011] <=  8'h00;      memory[51012] <=  8'h00;      memory[51013] <=  8'h00;      memory[51014] <=  8'h00;      memory[51015] <=  8'h00;      memory[51016] <=  8'h00;      memory[51017] <=  8'h00;      memory[51018] <=  8'h00;      memory[51019] <=  8'h00;      memory[51020] <=  8'h00;      memory[51021] <=  8'h00;      memory[51022] <=  8'h00;      memory[51023] <=  8'h00;      memory[51024] <=  8'h00;      memory[51025] <=  8'h00;      memory[51026] <=  8'h00;      memory[51027] <=  8'h00;      memory[51028] <=  8'h00;      memory[51029] <=  8'h00;      memory[51030] <=  8'h00;      memory[51031] <=  8'h00;      memory[51032] <=  8'h00;      memory[51033] <=  8'h00;      memory[51034] <=  8'h00;      memory[51035] <=  8'h00;      memory[51036] <=  8'h00;      memory[51037] <=  8'h00;      memory[51038] <=  8'h00;      memory[51039] <=  8'h00;      memory[51040] <=  8'h00;      memory[51041] <=  8'h00;      memory[51042] <=  8'h00;      memory[51043] <=  8'h00;      memory[51044] <=  8'h00;      memory[51045] <=  8'h00;      memory[51046] <=  8'h00;      memory[51047] <=  8'h00;      memory[51048] <=  8'h00;      memory[51049] <=  8'h00;      memory[51050] <=  8'h00;      memory[51051] <=  8'h00;      memory[51052] <=  8'h00;      memory[51053] <=  8'h00;      memory[51054] <=  8'h00;      memory[51055] <=  8'h00;      memory[51056] <=  8'h00;      memory[51057] <=  8'h00;      memory[51058] <=  8'h00;      memory[51059] <=  8'h00;      memory[51060] <=  8'h00;      memory[51061] <=  8'h00;      memory[51062] <=  8'h00;      memory[51063] <=  8'h00;      memory[51064] <=  8'h00;      memory[51065] <=  8'h00;      memory[51066] <=  8'h00;      memory[51067] <=  8'h00;      memory[51068] <=  8'h00;      memory[51069] <=  8'h00;      memory[51070] <=  8'h00;      memory[51071] <=  8'h00;      memory[51072] <=  8'h00;      memory[51073] <=  8'h00;      memory[51074] <=  8'h00;      memory[51075] <=  8'h00;      memory[51076] <=  8'h00;      memory[51077] <=  8'h00;      memory[51078] <=  8'h00;      memory[51079] <=  8'h00;      memory[51080] <=  8'h00;      memory[51081] <=  8'h00;      memory[51082] <=  8'h00;      memory[51083] <=  8'h00;      memory[51084] <=  8'h00;      memory[51085] <=  8'h00;      memory[51086] <=  8'h00;      memory[51087] <=  8'h00;      memory[51088] <=  8'h00;      memory[51089] <=  8'h00;      memory[51090] <=  8'h00;      memory[51091] <=  8'h00;      memory[51092] <=  8'h00;      memory[51093] <=  8'h00;      memory[51094] <=  8'h00;      memory[51095] <=  8'h00;      memory[51096] <=  8'h00;      memory[51097] <=  8'h00;      memory[51098] <=  8'h00;      memory[51099] <=  8'h00;      memory[51100] <=  8'h00;      memory[51101] <=  8'h00;      memory[51102] <=  8'h00;      memory[51103] <=  8'h00;      memory[51104] <=  8'h00;      memory[51105] <=  8'h00;      memory[51106] <=  8'h00;      memory[51107] <=  8'h00;      memory[51108] <=  8'h00;      memory[51109] <=  8'h00;      memory[51110] <=  8'h00;      memory[51111] <=  8'h00;      memory[51112] <=  8'h00;      memory[51113] <=  8'h00;      memory[51114] <=  8'h00;      memory[51115] <=  8'h00;      memory[51116] <=  8'h00;      memory[51117] <=  8'h00;      memory[51118] <=  8'h00;      memory[51119] <=  8'h00;      memory[51120] <=  8'h00;      memory[51121] <=  8'h00;      memory[51122] <=  8'h00;      memory[51123] <=  8'h00;      memory[51124] <=  8'h00;      memory[51125] <=  8'h00;      memory[51126] <=  8'h00;      memory[51127] <=  8'h00;      memory[51128] <=  8'h00;      memory[51129] <=  8'h00;      memory[51130] <=  8'h00;      memory[51131] <=  8'h00;      memory[51132] <=  8'h00;      memory[51133] <=  8'h00;      memory[51134] <=  8'h00;      memory[51135] <=  8'h00;      memory[51136] <=  8'h00;      memory[51137] <=  8'h00;      memory[51138] <=  8'h00;      memory[51139] <=  8'h00;      memory[51140] <=  8'h00;      memory[51141] <=  8'h00;      memory[51142] <=  8'h00;      memory[51143] <=  8'h00;      memory[51144] <=  8'h00;      memory[51145] <=  8'h00;      memory[51146] <=  8'h00;      memory[51147] <=  8'h00;      memory[51148] <=  8'h00;      memory[51149] <=  8'h00;      memory[51150] <=  8'h00;      memory[51151] <=  8'h00;      memory[51152] <=  8'h00;      memory[51153] <=  8'h00;      memory[51154] <=  8'h00;      memory[51155] <=  8'h00;      memory[51156] <=  8'h00;      memory[51157] <=  8'h00;      memory[51158] <=  8'h00;      memory[51159] <=  8'h00;      memory[51160] <=  8'h00;      memory[51161] <=  8'h00;      memory[51162] <=  8'h00;      memory[51163] <=  8'h00;      memory[51164] <=  8'h00;      memory[51165] <=  8'h00;      memory[51166] <=  8'h00;      memory[51167] <=  8'h00;      memory[51168] <=  8'h00;      memory[51169] <=  8'h00;      memory[51170] <=  8'h00;      memory[51171] <=  8'h00;      memory[51172] <=  8'h00;      memory[51173] <=  8'h00;      memory[51174] <=  8'h00;      memory[51175] <=  8'h00;      memory[51176] <=  8'h00;      memory[51177] <=  8'h00;      memory[51178] <=  8'h00;      memory[51179] <=  8'h00;      memory[51180] <=  8'h00;      memory[51181] <=  8'h00;      memory[51182] <=  8'h00;      memory[51183] <=  8'h00;      memory[51184] <=  8'h00;      memory[51185] <=  8'h00;      memory[51186] <=  8'h00;      memory[51187] <=  8'h00;      memory[51188] <=  8'h00;      memory[51189] <=  8'h00;      memory[51190] <=  8'h00;      memory[51191] <=  8'h00;      memory[51192] <=  8'h00;      memory[51193] <=  8'h00;      memory[51194] <=  8'h00;      memory[51195] <=  8'h00;      memory[51196] <=  8'h00;      memory[51197] <=  8'h00;      memory[51198] <=  8'h00;      memory[51199] <=  8'h00;      memory[51200] <=  8'h00;      memory[51201] <=  8'h00;      memory[51202] <=  8'h00;      memory[51203] <=  8'h00;      memory[51204] <=  8'h00;      memory[51205] <=  8'h00;      memory[51206] <=  8'h00;      memory[51207] <=  8'h00;      memory[51208] <=  8'h00;      memory[51209] <=  8'h00;      memory[51210] <=  8'h00;      memory[51211] <=  8'h00;      memory[51212] <=  8'h00;      memory[51213] <=  8'h00;      memory[51214] <=  8'h00;      memory[51215] <=  8'h00;      memory[51216] <=  8'h00;      memory[51217] <=  8'h00;      memory[51218] <=  8'h00;      memory[51219] <=  8'h00;      memory[51220] <=  8'h00;      memory[51221] <=  8'h00;      memory[51222] <=  8'h00;      memory[51223] <=  8'h00;      memory[51224] <=  8'h00;      memory[51225] <=  8'h00;      memory[51226] <=  8'h00;      memory[51227] <=  8'h00;      memory[51228] <=  8'h00;      memory[51229] <=  8'h00;      memory[51230] <=  8'h00;      memory[51231] <=  8'h00;      memory[51232] <=  8'h00;      memory[51233] <=  8'h00;      memory[51234] <=  8'h00;      memory[51235] <=  8'h00;      memory[51236] <=  8'h00;      memory[51237] <=  8'h00;      memory[51238] <=  8'h00;      memory[51239] <=  8'h00;      memory[51240] <=  8'h00;      memory[51241] <=  8'h00;      memory[51242] <=  8'h00;      memory[51243] <=  8'h00;      memory[51244] <=  8'h00;      memory[51245] <=  8'h00;      memory[51246] <=  8'h00;      memory[51247] <=  8'h00;      memory[51248] <=  8'h00;      memory[51249] <=  8'h00;      memory[51250] <=  8'h00;      memory[51251] <=  8'h00;      memory[51252] <=  8'h00;      memory[51253] <=  8'h00;      memory[51254] <=  8'h00;      memory[51255] <=  8'h00;      memory[51256] <=  8'h00;      memory[51257] <=  8'h00;      memory[51258] <=  8'h00;      memory[51259] <=  8'h00;      memory[51260] <=  8'h00;      memory[51261] <=  8'h00;      memory[51262] <=  8'h00;      memory[51263] <=  8'h00;      memory[51264] <=  8'h00;      memory[51265] <=  8'h00;      memory[51266] <=  8'h00;      memory[51267] <=  8'h00;      memory[51268] <=  8'h00;      memory[51269] <=  8'h00;      memory[51270] <=  8'h00;      memory[51271] <=  8'h00;      memory[51272] <=  8'h00;      memory[51273] <=  8'h00;      memory[51274] <=  8'h00;      memory[51275] <=  8'h00;      memory[51276] <=  8'h00;      memory[51277] <=  8'h00;      memory[51278] <=  8'h00;      memory[51279] <=  8'h00;      memory[51280] <=  8'h00;      memory[51281] <=  8'h00;      memory[51282] <=  8'h00;      memory[51283] <=  8'h00;      memory[51284] <=  8'h00;      memory[51285] <=  8'h00;      memory[51286] <=  8'h00;      memory[51287] <=  8'h00;      memory[51288] <=  8'h00;      memory[51289] <=  8'h00;      memory[51290] <=  8'h00;      memory[51291] <=  8'h00;      memory[51292] <=  8'h00;      memory[51293] <=  8'h00;      memory[51294] <=  8'h00;      memory[51295] <=  8'h00;      memory[51296] <=  8'h00;      memory[51297] <=  8'h00;      memory[51298] <=  8'h00;      memory[51299] <=  8'h00;      memory[51300] <=  8'h00;      memory[51301] <=  8'h00;      memory[51302] <=  8'h00;      memory[51303] <=  8'h00;      memory[51304] <=  8'h00;      memory[51305] <=  8'h00;      memory[51306] <=  8'h00;      memory[51307] <=  8'h00;      memory[51308] <=  8'h00;      memory[51309] <=  8'h00;      memory[51310] <=  8'h00;      memory[51311] <=  8'h00;      memory[51312] <=  8'h00;      memory[51313] <=  8'h00;      memory[51314] <=  8'h00;      memory[51315] <=  8'h00;      memory[51316] <=  8'h00;      memory[51317] <=  8'h00;      memory[51318] <=  8'h00;      memory[51319] <=  8'h00;      memory[51320] <=  8'h00;      memory[51321] <=  8'h00;      memory[51322] <=  8'h00;      memory[51323] <=  8'h00;      memory[51324] <=  8'h00;      memory[51325] <=  8'h00;      memory[51326] <=  8'h00;      memory[51327] <=  8'h00;      memory[51328] <=  8'h00;      memory[51329] <=  8'h00;      memory[51330] <=  8'h00;      memory[51331] <=  8'h00;      memory[51332] <=  8'h00;      memory[51333] <=  8'h00;      memory[51334] <=  8'h00;      memory[51335] <=  8'h00;      memory[51336] <=  8'h00;      memory[51337] <=  8'h00;      memory[51338] <=  8'h00;      memory[51339] <=  8'h00;      memory[51340] <=  8'h00;      memory[51341] <=  8'h00;      memory[51342] <=  8'h00;      memory[51343] <=  8'h00;      memory[51344] <=  8'h00;      memory[51345] <=  8'h00;      memory[51346] <=  8'h00;      memory[51347] <=  8'h00;      memory[51348] <=  8'h00;      memory[51349] <=  8'h00;      memory[51350] <=  8'h00;      memory[51351] <=  8'h00;      memory[51352] <=  8'h00;      memory[51353] <=  8'h00;      memory[51354] <=  8'h00;      memory[51355] <=  8'h00;      memory[51356] <=  8'h00;      memory[51357] <=  8'h00;      memory[51358] <=  8'h00;      memory[51359] <=  8'h00;      memory[51360] <=  8'h00;      memory[51361] <=  8'h00;      memory[51362] <=  8'h00;      memory[51363] <=  8'h00;      memory[51364] <=  8'h00;      memory[51365] <=  8'h00;      memory[51366] <=  8'h00;      memory[51367] <=  8'h00;      memory[51368] <=  8'h00;      memory[51369] <=  8'h00;      memory[51370] <=  8'h00;      memory[51371] <=  8'h00;      memory[51372] <=  8'h00;      memory[51373] <=  8'h00;      memory[51374] <=  8'h00;      memory[51375] <=  8'h00;      memory[51376] <=  8'h00;      memory[51377] <=  8'h00;      memory[51378] <=  8'h00;      memory[51379] <=  8'h00;      memory[51380] <=  8'h00;      memory[51381] <=  8'h00;      memory[51382] <=  8'h00;      memory[51383] <=  8'h00;      memory[51384] <=  8'h00;      memory[51385] <=  8'h00;      memory[51386] <=  8'h00;      memory[51387] <=  8'h00;      memory[51388] <=  8'h00;      memory[51389] <=  8'h00;      memory[51390] <=  8'h00;      memory[51391] <=  8'h00;      memory[51392] <=  8'h00;      memory[51393] <=  8'h00;      memory[51394] <=  8'h00;      memory[51395] <=  8'h00;      memory[51396] <=  8'h00;      memory[51397] <=  8'h00;      memory[51398] <=  8'h00;      memory[51399] <=  8'h00;      memory[51400] <=  8'h00;      memory[51401] <=  8'h00;      memory[51402] <=  8'h00;      memory[51403] <=  8'h00;      memory[51404] <=  8'h00;      memory[51405] <=  8'h00;      memory[51406] <=  8'h00;      memory[51407] <=  8'h00;      memory[51408] <=  8'h00;      memory[51409] <=  8'h00;      memory[51410] <=  8'h00;      memory[51411] <=  8'h00;      memory[51412] <=  8'h00;      memory[51413] <=  8'h00;      memory[51414] <=  8'h00;      memory[51415] <=  8'h00;      memory[51416] <=  8'h00;      memory[51417] <=  8'h00;      memory[51418] <=  8'h00;      memory[51419] <=  8'h00;      memory[51420] <=  8'h00;      memory[51421] <=  8'h00;      memory[51422] <=  8'h00;      memory[51423] <=  8'h00;      memory[51424] <=  8'h00;      memory[51425] <=  8'h00;      memory[51426] <=  8'h00;      memory[51427] <=  8'h00;      memory[51428] <=  8'h00;      memory[51429] <=  8'h00;      memory[51430] <=  8'h00;      memory[51431] <=  8'h00;      memory[51432] <=  8'h00;      memory[51433] <=  8'h00;      memory[51434] <=  8'h00;      memory[51435] <=  8'h00;      memory[51436] <=  8'h00;      memory[51437] <=  8'h00;      memory[51438] <=  8'h00;      memory[51439] <=  8'h00;      memory[51440] <=  8'h00;      memory[51441] <=  8'h00;      memory[51442] <=  8'h00;      memory[51443] <=  8'h00;      memory[51444] <=  8'h00;      memory[51445] <=  8'h00;      memory[51446] <=  8'h00;      memory[51447] <=  8'h00;      memory[51448] <=  8'h00;      memory[51449] <=  8'h00;      memory[51450] <=  8'h00;      memory[51451] <=  8'h00;      memory[51452] <=  8'h00;      memory[51453] <=  8'h00;      memory[51454] <=  8'h00;      memory[51455] <=  8'h00;      memory[51456] <=  8'h00;      memory[51457] <=  8'h00;      memory[51458] <=  8'h00;      memory[51459] <=  8'h00;      memory[51460] <=  8'h00;      memory[51461] <=  8'h00;      memory[51462] <=  8'h00;      memory[51463] <=  8'h00;      memory[51464] <=  8'h00;      memory[51465] <=  8'h00;      memory[51466] <=  8'h00;      memory[51467] <=  8'h00;      memory[51468] <=  8'h00;      memory[51469] <=  8'h00;      memory[51470] <=  8'h00;      memory[51471] <=  8'h00;      memory[51472] <=  8'h00;      memory[51473] <=  8'h00;      memory[51474] <=  8'h00;      memory[51475] <=  8'h00;      memory[51476] <=  8'h00;      memory[51477] <=  8'h00;      memory[51478] <=  8'h00;      memory[51479] <=  8'h00;      memory[51480] <=  8'h00;      memory[51481] <=  8'h00;      memory[51482] <=  8'h00;      memory[51483] <=  8'h00;      memory[51484] <=  8'h00;      memory[51485] <=  8'h00;      memory[51486] <=  8'h00;      memory[51487] <=  8'h00;      memory[51488] <=  8'h00;      memory[51489] <=  8'h00;      memory[51490] <=  8'h00;      memory[51491] <=  8'h00;      memory[51492] <=  8'h00;      memory[51493] <=  8'h00;      memory[51494] <=  8'h00;      memory[51495] <=  8'h00;      memory[51496] <=  8'h00;      memory[51497] <=  8'h00;      memory[51498] <=  8'h00;      memory[51499] <=  8'h00;      memory[51500] <=  8'h00;      memory[51501] <=  8'h00;      memory[51502] <=  8'h00;      memory[51503] <=  8'h00;      memory[51504] <=  8'h00;      memory[51505] <=  8'h00;      memory[51506] <=  8'h00;      memory[51507] <=  8'h00;      memory[51508] <=  8'h00;      memory[51509] <=  8'h00;      memory[51510] <=  8'h00;      memory[51511] <=  8'h00;      memory[51512] <=  8'h00;      memory[51513] <=  8'h00;      memory[51514] <=  8'h00;      memory[51515] <=  8'h00;      memory[51516] <=  8'h00;      memory[51517] <=  8'h00;      memory[51518] <=  8'h00;      memory[51519] <=  8'h00;      memory[51520] <=  8'h00;      memory[51521] <=  8'h00;      memory[51522] <=  8'h00;      memory[51523] <=  8'h00;      memory[51524] <=  8'h00;      memory[51525] <=  8'h00;      memory[51526] <=  8'h00;      memory[51527] <=  8'h00;      memory[51528] <=  8'h00;      memory[51529] <=  8'h00;      memory[51530] <=  8'h00;      memory[51531] <=  8'h00;      memory[51532] <=  8'h00;      memory[51533] <=  8'h00;      memory[51534] <=  8'h00;      memory[51535] <=  8'h00;      memory[51536] <=  8'h00;      memory[51537] <=  8'h00;      memory[51538] <=  8'h00;      memory[51539] <=  8'h00;      memory[51540] <=  8'h00;      memory[51541] <=  8'h00;      memory[51542] <=  8'h00;      memory[51543] <=  8'h00;      memory[51544] <=  8'h00;      memory[51545] <=  8'h00;      memory[51546] <=  8'h00;      memory[51547] <=  8'h00;      memory[51548] <=  8'h00;      memory[51549] <=  8'h00;      memory[51550] <=  8'h00;      memory[51551] <=  8'h00;      memory[51552] <=  8'h00;      memory[51553] <=  8'h00;      memory[51554] <=  8'h00;      memory[51555] <=  8'h00;      memory[51556] <=  8'h00;      memory[51557] <=  8'h00;      memory[51558] <=  8'h00;      memory[51559] <=  8'h00;      memory[51560] <=  8'h00;      memory[51561] <=  8'h00;      memory[51562] <=  8'h00;      memory[51563] <=  8'h00;      memory[51564] <=  8'h00;      memory[51565] <=  8'h00;      memory[51566] <=  8'h00;      memory[51567] <=  8'h00;      memory[51568] <=  8'h00;      memory[51569] <=  8'h00;      memory[51570] <=  8'h00;      memory[51571] <=  8'h00;      memory[51572] <=  8'h00;      memory[51573] <=  8'h00;      memory[51574] <=  8'h00;      memory[51575] <=  8'h00;      memory[51576] <=  8'h00;      memory[51577] <=  8'h00;      memory[51578] <=  8'h00;      memory[51579] <=  8'h00;      memory[51580] <=  8'h00;      memory[51581] <=  8'h00;      memory[51582] <=  8'h00;      memory[51583] <=  8'h00;      memory[51584] <=  8'h00;      memory[51585] <=  8'h00;      memory[51586] <=  8'h00;      memory[51587] <=  8'h00;      memory[51588] <=  8'h00;      memory[51589] <=  8'h00;      memory[51590] <=  8'h00;      memory[51591] <=  8'h00;      memory[51592] <=  8'h00;      memory[51593] <=  8'h00;      memory[51594] <=  8'h00;      memory[51595] <=  8'h00;      memory[51596] <=  8'h00;      memory[51597] <=  8'h00;      memory[51598] <=  8'h00;      memory[51599] <=  8'h00;      memory[51600] <=  8'h00;      memory[51601] <=  8'h00;      memory[51602] <=  8'h00;      memory[51603] <=  8'h00;      memory[51604] <=  8'h00;      memory[51605] <=  8'h00;      memory[51606] <=  8'h00;      memory[51607] <=  8'h00;      memory[51608] <=  8'h00;      memory[51609] <=  8'h00;      memory[51610] <=  8'h00;      memory[51611] <=  8'h00;      memory[51612] <=  8'h00;      memory[51613] <=  8'h00;      memory[51614] <=  8'h00;      memory[51615] <=  8'h00;      memory[51616] <=  8'h00;      memory[51617] <=  8'h00;      memory[51618] <=  8'h00;      memory[51619] <=  8'h00;      memory[51620] <=  8'h00;      memory[51621] <=  8'h00;      memory[51622] <=  8'h00;      memory[51623] <=  8'h00;      memory[51624] <=  8'h00;      memory[51625] <=  8'h00;      memory[51626] <=  8'h00;      memory[51627] <=  8'h00;      memory[51628] <=  8'h00;      memory[51629] <=  8'h00;      memory[51630] <=  8'h00;      memory[51631] <=  8'h00;      memory[51632] <=  8'h00;      memory[51633] <=  8'h00;      memory[51634] <=  8'h00;      memory[51635] <=  8'h00;      memory[51636] <=  8'h00;      memory[51637] <=  8'h00;      memory[51638] <=  8'h00;      memory[51639] <=  8'h00;      memory[51640] <=  8'h00;      memory[51641] <=  8'h00;      memory[51642] <=  8'h00;      memory[51643] <=  8'h00;      memory[51644] <=  8'h00;      memory[51645] <=  8'h00;      memory[51646] <=  8'h00;      memory[51647] <=  8'h00;      memory[51648] <=  8'h00;      memory[51649] <=  8'h00;      memory[51650] <=  8'h00;      memory[51651] <=  8'h00;      memory[51652] <=  8'h00;      memory[51653] <=  8'h00;      memory[51654] <=  8'h00;      memory[51655] <=  8'h00;      memory[51656] <=  8'h00;      memory[51657] <=  8'h00;      memory[51658] <=  8'h00;      memory[51659] <=  8'h00;      memory[51660] <=  8'h00;      memory[51661] <=  8'h00;      memory[51662] <=  8'h00;      memory[51663] <=  8'h00;      memory[51664] <=  8'h00;      memory[51665] <=  8'h00;      memory[51666] <=  8'h00;      memory[51667] <=  8'h00;      memory[51668] <=  8'h00;      memory[51669] <=  8'h00;      memory[51670] <=  8'h00;      memory[51671] <=  8'h00;      memory[51672] <=  8'h00;      memory[51673] <=  8'h00;      memory[51674] <=  8'h00;      memory[51675] <=  8'h00;      memory[51676] <=  8'h00;      memory[51677] <=  8'h00;      memory[51678] <=  8'h00;      memory[51679] <=  8'h00;      memory[51680] <=  8'h00;      memory[51681] <=  8'h00;      memory[51682] <=  8'h00;      memory[51683] <=  8'h00;      memory[51684] <=  8'h00;      memory[51685] <=  8'h00;      memory[51686] <=  8'h00;      memory[51687] <=  8'h00;      memory[51688] <=  8'h00;      memory[51689] <=  8'h00;      memory[51690] <=  8'h00;      memory[51691] <=  8'h00;      memory[51692] <=  8'h00;      memory[51693] <=  8'h00;      memory[51694] <=  8'h00;      memory[51695] <=  8'h00;      memory[51696] <=  8'h00;      memory[51697] <=  8'h00;      memory[51698] <=  8'h00;      memory[51699] <=  8'h00;      memory[51700] <=  8'h00;      memory[51701] <=  8'h00;      memory[51702] <=  8'h00;      memory[51703] <=  8'h00;      memory[51704] <=  8'h00;      memory[51705] <=  8'h00;      memory[51706] <=  8'h00;      memory[51707] <=  8'h00;      memory[51708] <=  8'h00;      memory[51709] <=  8'h00;      memory[51710] <=  8'h00;      memory[51711] <=  8'h00;      memory[51712] <=  8'h00;      memory[51713] <=  8'h00;      memory[51714] <=  8'h00;      memory[51715] <=  8'h00;      memory[51716] <=  8'h00;      memory[51717] <=  8'h00;      memory[51718] <=  8'h00;      memory[51719] <=  8'h00;      memory[51720] <=  8'h00;      memory[51721] <=  8'h00;      memory[51722] <=  8'h00;      memory[51723] <=  8'h00;      memory[51724] <=  8'h00;      memory[51725] <=  8'h00;      memory[51726] <=  8'h00;      memory[51727] <=  8'h00;      memory[51728] <=  8'h00;      memory[51729] <=  8'h00;      memory[51730] <=  8'h00;      memory[51731] <=  8'h00;      memory[51732] <=  8'h00;      memory[51733] <=  8'h00;      memory[51734] <=  8'h00;      memory[51735] <=  8'h00;      memory[51736] <=  8'h00;      memory[51737] <=  8'h00;      memory[51738] <=  8'h00;      memory[51739] <=  8'h00;      memory[51740] <=  8'h00;      memory[51741] <=  8'h00;      memory[51742] <=  8'h00;      memory[51743] <=  8'h00;      memory[51744] <=  8'h00;      memory[51745] <=  8'h00;      memory[51746] <=  8'h00;      memory[51747] <=  8'h00;      memory[51748] <=  8'h00;      memory[51749] <=  8'h00;      memory[51750] <=  8'h00;      memory[51751] <=  8'h00;      memory[51752] <=  8'h00;      memory[51753] <=  8'h00;      memory[51754] <=  8'h00;      memory[51755] <=  8'h00;      memory[51756] <=  8'h00;      memory[51757] <=  8'h00;      memory[51758] <=  8'h00;      memory[51759] <=  8'h00;      memory[51760] <=  8'h00;      memory[51761] <=  8'h00;      memory[51762] <=  8'h00;      memory[51763] <=  8'h00;      memory[51764] <=  8'h00;      memory[51765] <=  8'h00;      memory[51766] <=  8'h00;      memory[51767] <=  8'h00;      memory[51768] <=  8'h00;      memory[51769] <=  8'h00;      memory[51770] <=  8'h00;      memory[51771] <=  8'h00;      memory[51772] <=  8'h00;      memory[51773] <=  8'h00;      memory[51774] <=  8'h00;      memory[51775] <=  8'h00;      memory[51776] <=  8'h00;      memory[51777] <=  8'h00;      memory[51778] <=  8'h00;      memory[51779] <=  8'h00;      memory[51780] <=  8'h00;      memory[51781] <=  8'h00;      memory[51782] <=  8'h00;      memory[51783] <=  8'h00;      memory[51784] <=  8'h00;      memory[51785] <=  8'h00;      memory[51786] <=  8'h00;      memory[51787] <=  8'h00;      memory[51788] <=  8'h00;      memory[51789] <=  8'h00;      memory[51790] <=  8'h00;      memory[51791] <=  8'h00;      memory[51792] <=  8'h00;      memory[51793] <=  8'h00;      memory[51794] <=  8'h00;      memory[51795] <=  8'h00;      memory[51796] <=  8'h00;      memory[51797] <=  8'h00;      memory[51798] <=  8'h00;      memory[51799] <=  8'h00;      memory[51800] <=  8'h00;      memory[51801] <=  8'h00;      memory[51802] <=  8'h00;      memory[51803] <=  8'h00;      memory[51804] <=  8'h00;      memory[51805] <=  8'h00;      memory[51806] <=  8'h00;      memory[51807] <=  8'h00;      memory[51808] <=  8'h00;      memory[51809] <=  8'h00;      memory[51810] <=  8'h00;      memory[51811] <=  8'h00;      memory[51812] <=  8'h00;      memory[51813] <=  8'h00;      memory[51814] <=  8'h00;      memory[51815] <=  8'h00;      memory[51816] <=  8'h00;      memory[51817] <=  8'h00;      memory[51818] <=  8'h00;      memory[51819] <=  8'h00;      memory[51820] <=  8'h00;      memory[51821] <=  8'h00;      memory[51822] <=  8'h00;      memory[51823] <=  8'h00;      memory[51824] <=  8'h00;      memory[51825] <=  8'h00;      memory[51826] <=  8'h00;      memory[51827] <=  8'h00;      memory[51828] <=  8'h00;      memory[51829] <=  8'h00;      memory[51830] <=  8'h00;      memory[51831] <=  8'h00;      memory[51832] <=  8'h00;      memory[51833] <=  8'h00;      memory[51834] <=  8'h00;      memory[51835] <=  8'h00;      memory[51836] <=  8'h00;      memory[51837] <=  8'h00;      memory[51838] <=  8'h00;      memory[51839] <=  8'h00;      memory[51840] <=  8'h00;      memory[51841] <=  8'h00;      memory[51842] <=  8'h00;      memory[51843] <=  8'h00;      memory[51844] <=  8'h00;      memory[51845] <=  8'h00;      memory[51846] <=  8'h00;      memory[51847] <=  8'h00;      memory[51848] <=  8'h00;      memory[51849] <=  8'h00;      memory[51850] <=  8'h00;      memory[51851] <=  8'h00;      memory[51852] <=  8'h00;      memory[51853] <=  8'h00;      memory[51854] <=  8'h00;      memory[51855] <=  8'h00;      memory[51856] <=  8'h00;      memory[51857] <=  8'h00;      memory[51858] <=  8'h00;      memory[51859] <=  8'h00;      memory[51860] <=  8'h00;      memory[51861] <=  8'h00;      memory[51862] <=  8'h00;      memory[51863] <=  8'h00;      memory[51864] <=  8'h00;      memory[51865] <=  8'h00;      memory[51866] <=  8'h00;      memory[51867] <=  8'h00;      memory[51868] <=  8'h00;      memory[51869] <=  8'h00;      memory[51870] <=  8'h00;      memory[51871] <=  8'h00;      memory[51872] <=  8'h00;      memory[51873] <=  8'h00;      memory[51874] <=  8'h00;      memory[51875] <=  8'h00;      memory[51876] <=  8'h00;      memory[51877] <=  8'h00;      memory[51878] <=  8'h00;      memory[51879] <=  8'h00;      memory[51880] <=  8'h00;      memory[51881] <=  8'h00;      memory[51882] <=  8'h00;      memory[51883] <=  8'h00;      memory[51884] <=  8'h00;      memory[51885] <=  8'h00;      memory[51886] <=  8'h00;      memory[51887] <=  8'h00;      memory[51888] <=  8'h00;      memory[51889] <=  8'h00;      memory[51890] <=  8'h00;      memory[51891] <=  8'h00;      memory[51892] <=  8'h00;      memory[51893] <=  8'h00;      memory[51894] <=  8'h00;      memory[51895] <=  8'h00;      memory[51896] <=  8'h00;      memory[51897] <=  8'h00;      memory[51898] <=  8'h00;      memory[51899] <=  8'h00;      memory[51900] <=  8'h00;      memory[51901] <=  8'h00;      memory[51902] <=  8'h00;      memory[51903] <=  8'h00;      memory[51904] <=  8'h00;      memory[51905] <=  8'h00;      memory[51906] <=  8'h00;      memory[51907] <=  8'h00;      memory[51908] <=  8'h00;      memory[51909] <=  8'h00;      memory[51910] <=  8'h00;      memory[51911] <=  8'h00;      memory[51912] <=  8'h00;      memory[51913] <=  8'h00;      memory[51914] <=  8'h00;      memory[51915] <=  8'h00;      memory[51916] <=  8'h00;      memory[51917] <=  8'h00;      memory[51918] <=  8'h00;      memory[51919] <=  8'h00;      memory[51920] <=  8'h00;      memory[51921] <=  8'h00;      memory[51922] <=  8'h00;      memory[51923] <=  8'h00;      memory[51924] <=  8'h00;      memory[51925] <=  8'h00;      memory[51926] <=  8'h00;      memory[51927] <=  8'h00;      memory[51928] <=  8'h00;      memory[51929] <=  8'h00;      memory[51930] <=  8'h00;      memory[51931] <=  8'h00;      memory[51932] <=  8'h00;      memory[51933] <=  8'h00;      memory[51934] <=  8'h00;      memory[51935] <=  8'h00;      memory[51936] <=  8'h00;      memory[51937] <=  8'h00;      memory[51938] <=  8'h00;      memory[51939] <=  8'h00;      memory[51940] <=  8'h00;      memory[51941] <=  8'h00;      memory[51942] <=  8'h00;      memory[51943] <=  8'h00;      memory[51944] <=  8'h00;      memory[51945] <=  8'h00;      memory[51946] <=  8'h00;      memory[51947] <=  8'h00;      memory[51948] <=  8'h00;      memory[51949] <=  8'h00;      memory[51950] <=  8'h00;      memory[51951] <=  8'h00;      memory[51952] <=  8'h00;      memory[51953] <=  8'h00;      memory[51954] <=  8'h00;      memory[51955] <=  8'h00;      memory[51956] <=  8'h00;      memory[51957] <=  8'h00;      memory[51958] <=  8'h00;      memory[51959] <=  8'h00;      memory[51960] <=  8'h00;      memory[51961] <=  8'h00;      memory[51962] <=  8'h00;      memory[51963] <=  8'h00;      memory[51964] <=  8'h00;      memory[51965] <=  8'h00;      memory[51966] <=  8'h00;      memory[51967] <=  8'h00;      memory[51968] <=  8'h00;      memory[51969] <=  8'h00;      memory[51970] <=  8'h00;      memory[51971] <=  8'h00;      memory[51972] <=  8'h00;      memory[51973] <=  8'h00;      memory[51974] <=  8'h00;      memory[51975] <=  8'h00;      memory[51976] <=  8'h00;      memory[51977] <=  8'h00;      memory[51978] <=  8'h00;      memory[51979] <=  8'h00;      memory[51980] <=  8'h00;      memory[51981] <=  8'h00;      memory[51982] <=  8'h00;      memory[51983] <=  8'h00;      memory[51984] <=  8'h00;      memory[51985] <=  8'h00;      memory[51986] <=  8'h00;      memory[51987] <=  8'h00;      memory[51988] <=  8'h00;      memory[51989] <=  8'h00;      memory[51990] <=  8'h00;      memory[51991] <=  8'h00;      memory[51992] <=  8'h00;      memory[51993] <=  8'h00;      memory[51994] <=  8'h00;      memory[51995] <=  8'h00;      memory[51996] <=  8'h00;      memory[51997] <=  8'h00;      memory[51998] <=  8'h00;      memory[51999] <=  8'h00;      memory[52000] <=  8'h00;      memory[52001] <=  8'h00;      memory[52002] <=  8'h00;      memory[52003] <=  8'h00;      memory[52004] <=  8'h00;      memory[52005] <=  8'h00;      memory[52006] <=  8'h00;      memory[52007] <=  8'h00;      memory[52008] <=  8'h00;      memory[52009] <=  8'h00;      memory[52010] <=  8'h00;      memory[52011] <=  8'h00;      memory[52012] <=  8'h00;      memory[52013] <=  8'h00;      memory[52014] <=  8'h00;      memory[52015] <=  8'h00;      memory[52016] <=  8'h00;      memory[52017] <=  8'h00;      memory[52018] <=  8'h00;      memory[52019] <=  8'h00;      memory[52020] <=  8'h00;      memory[52021] <=  8'h00;      memory[52022] <=  8'h00;      memory[52023] <=  8'h00;      memory[52024] <=  8'h00;      memory[52025] <=  8'h00;      memory[52026] <=  8'h00;      memory[52027] <=  8'h00;      memory[52028] <=  8'h00;      memory[52029] <=  8'h00;      memory[52030] <=  8'h00;      memory[52031] <=  8'h00;      memory[52032] <=  8'h00;      memory[52033] <=  8'h00;      memory[52034] <=  8'h00;      memory[52035] <=  8'h00;      memory[52036] <=  8'h00;      memory[52037] <=  8'h00;      memory[52038] <=  8'h00;      memory[52039] <=  8'h00;      memory[52040] <=  8'h00;      memory[52041] <=  8'h00;      memory[52042] <=  8'h00;      memory[52043] <=  8'h00;      memory[52044] <=  8'h00;      memory[52045] <=  8'h00;      memory[52046] <=  8'h00;      memory[52047] <=  8'h00;      memory[52048] <=  8'h00;      memory[52049] <=  8'h00;      memory[52050] <=  8'h00;      memory[52051] <=  8'h00;      memory[52052] <=  8'h00;      memory[52053] <=  8'h00;      memory[52054] <=  8'h00;      memory[52055] <=  8'h00;      memory[52056] <=  8'h00;      memory[52057] <=  8'h00;      memory[52058] <=  8'h00;      memory[52059] <=  8'h00;      memory[52060] <=  8'h00;      memory[52061] <=  8'h00;      memory[52062] <=  8'h00;      memory[52063] <=  8'h00;      memory[52064] <=  8'h00;      memory[52065] <=  8'h00;      memory[52066] <=  8'h00;      memory[52067] <=  8'h00;      memory[52068] <=  8'h00;      memory[52069] <=  8'h00;      memory[52070] <=  8'h00;      memory[52071] <=  8'h00;      memory[52072] <=  8'h00;      memory[52073] <=  8'h00;      memory[52074] <=  8'h00;      memory[52075] <=  8'h00;      memory[52076] <=  8'h00;      memory[52077] <=  8'h00;      memory[52078] <=  8'h00;      memory[52079] <=  8'h00;      memory[52080] <=  8'h00;      memory[52081] <=  8'h00;      memory[52082] <=  8'h00;      memory[52083] <=  8'h00;      memory[52084] <=  8'h00;      memory[52085] <=  8'h00;      memory[52086] <=  8'h00;      memory[52087] <=  8'h00;      memory[52088] <=  8'h00;      memory[52089] <=  8'h00;      memory[52090] <=  8'h00;      memory[52091] <=  8'h00;      memory[52092] <=  8'h00;      memory[52093] <=  8'h00;      memory[52094] <=  8'h00;      memory[52095] <=  8'h00;      memory[52096] <=  8'h00;      memory[52097] <=  8'h00;      memory[52098] <=  8'h00;      memory[52099] <=  8'h00;      memory[52100] <=  8'h00;      memory[52101] <=  8'h00;      memory[52102] <=  8'h00;      memory[52103] <=  8'h00;      memory[52104] <=  8'h00;      memory[52105] <=  8'h00;      memory[52106] <=  8'h00;      memory[52107] <=  8'h00;      memory[52108] <=  8'h00;      memory[52109] <=  8'h00;      memory[52110] <=  8'h00;      memory[52111] <=  8'h00;      memory[52112] <=  8'h00;      memory[52113] <=  8'h00;      memory[52114] <=  8'h00;      memory[52115] <=  8'h00;      memory[52116] <=  8'h00;      memory[52117] <=  8'h00;      memory[52118] <=  8'h00;      memory[52119] <=  8'h00;      memory[52120] <=  8'h00;      memory[52121] <=  8'h00;      memory[52122] <=  8'h00;      memory[52123] <=  8'h00;      memory[52124] <=  8'h00;      memory[52125] <=  8'h00;      memory[52126] <=  8'h00;      memory[52127] <=  8'h00;      memory[52128] <=  8'h00;      memory[52129] <=  8'h00;      memory[52130] <=  8'h00;      memory[52131] <=  8'h00;      memory[52132] <=  8'h00;      memory[52133] <=  8'h00;      memory[52134] <=  8'h00;      memory[52135] <=  8'h00;      memory[52136] <=  8'h00;      memory[52137] <=  8'h00;      memory[52138] <=  8'h00;      memory[52139] <=  8'h00;      memory[52140] <=  8'h00;      memory[52141] <=  8'h00;      memory[52142] <=  8'h00;      memory[52143] <=  8'h00;      memory[52144] <=  8'h00;      memory[52145] <=  8'h00;      memory[52146] <=  8'h00;      memory[52147] <=  8'h00;      memory[52148] <=  8'h00;      memory[52149] <=  8'h00;      memory[52150] <=  8'h00;      memory[52151] <=  8'h00;      memory[52152] <=  8'h00;      memory[52153] <=  8'h00;      memory[52154] <=  8'h00;      memory[52155] <=  8'h00;      memory[52156] <=  8'h00;      memory[52157] <=  8'h00;      memory[52158] <=  8'h00;      memory[52159] <=  8'h00;      memory[52160] <=  8'h00;      memory[52161] <=  8'h00;      memory[52162] <=  8'h00;      memory[52163] <=  8'h00;      memory[52164] <=  8'h00;      memory[52165] <=  8'h00;      memory[52166] <=  8'h00;      memory[52167] <=  8'h00;      memory[52168] <=  8'h00;      memory[52169] <=  8'h00;      memory[52170] <=  8'h00;      memory[52171] <=  8'h00;      memory[52172] <=  8'h00;      memory[52173] <=  8'h00;      memory[52174] <=  8'h00;      memory[52175] <=  8'h00;      memory[52176] <=  8'h00;      memory[52177] <=  8'h00;      memory[52178] <=  8'h00;      memory[52179] <=  8'h00;      memory[52180] <=  8'h00;      memory[52181] <=  8'h00;      memory[52182] <=  8'h00;      memory[52183] <=  8'h00;      memory[52184] <=  8'h00;      memory[52185] <=  8'h00;      memory[52186] <=  8'h00;      memory[52187] <=  8'h00;      memory[52188] <=  8'h00;      memory[52189] <=  8'h00;      memory[52190] <=  8'h00;      memory[52191] <=  8'h00;      memory[52192] <=  8'h00;      memory[52193] <=  8'h00;      memory[52194] <=  8'h00;      memory[52195] <=  8'h00;      memory[52196] <=  8'h00;      memory[52197] <=  8'h00;      memory[52198] <=  8'h00;      memory[52199] <=  8'h00;      memory[52200] <=  8'h00;      memory[52201] <=  8'h00;      memory[52202] <=  8'h00;      memory[52203] <=  8'h00;      memory[52204] <=  8'h00;      memory[52205] <=  8'h00;      memory[52206] <=  8'h00;      memory[52207] <=  8'h00;      memory[52208] <=  8'h00;      memory[52209] <=  8'h00;      memory[52210] <=  8'h00;      memory[52211] <=  8'h00;      memory[52212] <=  8'h00;      memory[52213] <=  8'h00;      memory[52214] <=  8'h00;      memory[52215] <=  8'h00;      memory[52216] <=  8'h00;      memory[52217] <=  8'h00;      memory[52218] <=  8'h00;      memory[52219] <=  8'h00;      memory[52220] <=  8'h00;      memory[52221] <=  8'h00;      memory[52222] <=  8'h00;      memory[52223] <=  8'h00;      memory[52224] <=  8'h00;      memory[52225] <=  8'h00;      memory[52226] <=  8'h00;      memory[52227] <=  8'h00;      memory[52228] <=  8'h00;      memory[52229] <=  8'h00;      memory[52230] <=  8'h00;      memory[52231] <=  8'h00;      memory[52232] <=  8'h00;      memory[52233] <=  8'h00;      memory[52234] <=  8'h00;      memory[52235] <=  8'h00;      memory[52236] <=  8'h00;      memory[52237] <=  8'h00;      memory[52238] <=  8'h00;      memory[52239] <=  8'h00;      memory[52240] <=  8'h00;      memory[52241] <=  8'h00;      memory[52242] <=  8'h00;      memory[52243] <=  8'h00;      memory[52244] <=  8'h00;      memory[52245] <=  8'h00;      memory[52246] <=  8'h00;      memory[52247] <=  8'h00;      memory[52248] <=  8'h00;      memory[52249] <=  8'h00;      memory[52250] <=  8'h00;      memory[52251] <=  8'h00;      memory[52252] <=  8'h00;      memory[52253] <=  8'h00;      memory[52254] <=  8'h00;      memory[52255] <=  8'h00;      memory[52256] <=  8'h00;      memory[52257] <=  8'h00;      memory[52258] <=  8'h00;      memory[52259] <=  8'h00;      memory[52260] <=  8'h00;      memory[52261] <=  8'h00;      memory[52262] <=  8'h00;      memory[52263] <=  8'h00;      memory[52264] <=  8'h00;      memory[52265] <=  8'h00;      memory[52266] <=  8'h00;      memory[52267] <=  8'h00;      memory[52268] <=  8'h00;      memory[52269] <=  8'h00;      memory[52270] <=  8'h00;      memory[52271] <=  8'h00;      memory[52272] <=  8'h00;      memory[52273] <=  8'h00;      memory[52274] <=  8'h00;      memory[52275] <=  8'h00;      memory[52276] <=  8'h00;      memory[52277] <=  8'h00;      memory[52278] <=  8'h00;      memory[52279] <=  8'h00;      memory[52280] <=  8'h00;      memory[52281] <=  8'h00;      memory[52282] <=  8'h00;      memory[52283] <=  8'h00;      memory[52284] <=  8'h00;      memory[52285] <=  8'h00;      memory[52286] <=  8'h00;      memory[52287] <=  8'h00;      memory[52288] <=  8'h00;      memory[52289] <=  8'h00;      memory[52290] <=  8'h00;      memory[52291] <=  8'h00;      memory[52292] <=  8'h00;      memory[52293] <=  8'h00;      memory[52294] <=  8'h00;      memory[52295] <=  8'h00;      memory[52296] <=  8'h00;      memory[52297] <=  8'h00;      memory[52298] <=  8'h00;      memory[52299] <=  8'h00;      memory[52300] <=  8'h00;      memory[52301] <=  8'h00;      memory[52302] <=  8'h00;      memory[52303] <=  8'h00;      memory[52304] <=  8'h00;      memory[52305] <=  8'h00;      memory[52306] <=  8'h00;      memory[52307] <=  8'h00;      memory[52308] <=  8'h00;      memory[52309] <=  8'h00;      memory[52310] <=  8'h00;      memory[52311] <=  8'h00;      memory[52312] <=  8'h00;      memory[52313] <=  8'h00;      memory[52314] <=  8'h00;      memory[52315] <=  8'h00;      memory[52316] <=  8'h00;      memory[52317] <=  8'h00;      memory[52318] <=  8'h00;      memory[52319] <=  8'h00;      memory[52320] <=  8'h00;      memory[52321] <=  8'h00;      memory[52322] <=  8'h00;      memory[52323] <=  8'h00;      memory[52324] <=  8'h00;      memory[52325] <=  8'h00;      memory[52326] <=  8'h00;      memory[52327] <=  8'h00;      memory[52328] <=  8'h00;      memory[52329] <=  8'h00;      memory[52330] <=  8'h00;      memory[52331] <=  8'h00;      memory[52332] <=  8'h00;      memory[52333] <=  8'h00;      memory[52334] <=  8'h00;      memory[52335] <=  8'h00;      memory[52336] <=  8'h00;      memory[52337] <=  8'h00;      memory[52338] <=  8'h00;      memory[52339] <=  8'h00;      memory[52340] <=  8'h00;      memory[52341] <=  8'h00;      memory[52342] <=  8'h00;      memory[52343] <=  8'h00;      memory[52344] <=  8'h00;      memory[52345] <=  8'h00;      memory[52346] <=  8'h00;      memory[52347] <=  8'h00;      memory[52348] <=  8'h00;      memory[52349] <=  8'h00;      memory[52350] <=  8'h00;      memory[52351] <=  8'h00;      memory[52352] <=  8'h00;      memory[52353] <=  8'h00;      memory[52354] <=  8'h00;      memory[52355] <=  8'h00;      memory[52356] <=  8'h00;      memory[52357] <=  8'h00;      memory[52358] <=  8'h00;      memory[52359] <=  8'h00;      memory[52360] <=  8'h00;      memory[52361] <=  8'h00;      memory[52362] <=  8'h00;      memory[52363] <=  8'h00;      memory[52364] <=  8'h00;      memory[52365] <=  8'h00;      memory[52366] <=  8'h00;      memory[52367] <=  8'h00;      memory[52368] <=  8'h00;      memory[52369] <=  8'h00;      memory[52370] <=  8'h00;      memory[52371] <=  8'h00;      memory[52372] <=  8'h00;      memory[52373] <=  8'h00;      memory[52374] <=  8'h00;      memory[52375] <=  8'h00;      memory[52376] <=  8'h00;      memory[52377] <=  8'h00;      memory[52378] <=  8'h00;      memory[52379] <=  8'h00;      memory[52380] <=  8'h00;      memory[52381] <=  8'h00;      memory[52382] <=  8'h00;      memory[52383] <=  8'h00;      memory[52384] <=  8'h00;      memory[52385] <=  8'h00;      memory[52386] <=  8'h00;      memory[52387] <=  8'h00;      memory[52388] <=  8'h00;      memory[52389] <=  8'h00;      memory[52390] <=  8'h00;      memory[52391] <=  8'h00;      memory[52392] <=  8'h00;      memory[52393] <=  8'h00;      memory[52394] <=  8'h00;      memory[52395] <=  8'h00;      memory[52396] <=  8'h00;      memory[52397] <=  8'h00;      memory[52398] <=  8'h00;      memory[52399] <=  8'h00;      memory[52400] <=  8'h00;      memory[52401] <=  8'h00;      memory[52402] <=  8'h00;      memory[52403] <=  8'h00;      memory[52404] <=  8'h00;      memory[52405] <=  8'h00;      memory[52406] <=  8'h00;      memory[52407] <=  8'h00;      memory[52408] <=  8'h00;      memory[52409] <=  8'h00;      memory[52410] <=  8'h00;      memory[52411] <=  8'h00;      memory[52412] <=  8'h00;      memory[52413] <=  8'h00;      memory[52414] <=  8'h00;      memory[52415] <=  8'h00;      memory[52416] <=  8'h00;      memory[52417] <=  8'h00;      memory[52418] <=  8'h00;      memory[52419] <=  8'h00;      memory[52420] <=  8'h00;      memory[52421] <=  8'h00;      memory[52422] <=  8'h00;      memory[52423] <=  8'h00;      memory[52424] <=  8'h00;      memory[52425] <=  8'h00;      memory[52426] <=  8'h00;      memory[52427] <=  8'h00;      memory[52428] <=  8'h00;      memory[52429] <=  8'h00;      memory[52430] <=  8'h00;      memory[52431] <=  8'h00;      memory[52432] <=  8'h00;      memory[52433] <=  8'h00;      memory[52434] <=  8'h00;      memory[52435] <=  8'h00;      memory[52436] <=  8'h00;      memory[52437] <=  8'h00;      memory[52438] <=  8'h00;      memory[52439] <=  8'h00;      memory[52440] <=  8'h00;      memory[52441] <=  8'h00;      memory[52442] <=  8'h00;      memory[52443] <=  8'h00;      memory[52444] <=  8'h00;      memory[52445] <=  8'h00;      memory[52446] <=  8'h00;      memory[52447] <=  8'h00;      memory[52448] <=  8'h00;      memory[52449] <=  8'h00;      memory[52450] <=  8'h00;      memory[52451] <=  8'h00;      memory[52452] <=  8'h00;      memory[52453] <=  8'h00;      memory[52454] <=  8'h00;      memory[52455] <=  8'h00;      memory[52456] <=  8'h00;      memory[52457] <=  8'h00;      memory[52458] <=  8'h00;      memory[52459] <=  8'h00;      memory[52460] <=  8'h00;      memory[52461] <=  8'h00;      memory[52462] <=  8'h00;      memory[52463] <=  8'h00;      memory[52464] <=  8'h00;      memory[52465] <=  8'h00;      memory[52466] <=  8'h00;      memory[52467] <=  8'h00;      memory[52468] <=  8'h00;      memory[52469] <=  8'h00;      memory[52470] <=  8'h00;      memory[52471] <=  8'h00;      memory[52472] <=  8'h00;      memory[52473] <=  8'h00;      memory[52474] <=  8'h00;      memory[52475] <=  8'h00;      memory[52476] <=  8'h00;      memory[52477] <=  8'h00;      memory[52478] <=  8'h00;      memory[52479] <=  8'h00;      memory[52480] <=  8'h00;      memory[52481] <=  8'h00;      memory[52482] <=  8'h00;      memory[52483] <=  8'h00;      memory[52484] <=  8'h00;      memory[52485] <=  8'h00;      memory[52486] <=  8'h00;      memory[52487] <=  8'h00;      memory[52488] <=  8'h00;      memory[52489] <=  8'h00;      memory[52490] <=  8'h00;      memory[52491] <=  8'h00;      memory[52492] <=  8'h00;      memory[52493] <=  8'h00;      memory[52494] <=  8'h00;      memory[52495] <=  8'h00;      memory[52496] <=  8'h00;      memory[52497] <=  8'h00;      memory[52498] <=  8'h00;      memory[52499] <=  8'h00;      memory[52500] <=  8'h00;      memory[52501] <=  8'h00;      memory[52502] <=  8'h00;      memory[52503] <=  8'h00;      memory[52504] <=  8'h00;      memory[52505] <=  8'h00;      memory[52506] <=  8'h00;      memory[52507] <=  8'h00;      memory[52508] <=  8'h00;      memory[52509] <=  8'h00;      memory[52510] <=  8'h00;      memory[52511] <=  8'h00;      memory[52512] <=  8'h00;      memory[52513] <=  8'h00;      memory[52514] <=  8'h00;      memory[52515] <=  8'h00;      memory[52516] <=  8'h00;      memory[52517] <=  8'h00;      memory[52518] <=  8'h00;      memory[52519] <=  8'h00;      memory[52520] <=  8'h00;      memory[52521] <=  8'h00;      memory[52522] <=  8'h00;      memory[52523] <=  8'h00;      memory[52524] <=  8'h00;      memory[52525] <=  8'h00;      memory[52526] <=  8'h00;      memory[52527] <=  8'h00;      memory[52528] <=  8'h00;      memory[52529] <=  8'h00;      memory[52530] <=  8'h00;      memory[52531] <=  8'h00;      memory[52532] <=  8'h00;      memory[52533] <=  8'h00;      memory[52534] <=  8'h00;      memory[52535] <=  8'h00;      memory[52536] <=  8'h00;      memory[52537] <=  8'h00;      memory[52538] <=  8'h00;      memory[52539] <=  8'h00;      memory[52540] <=  8'h00;      memory[52541] <=  8'h00;      memory[52542] <=  8'h00;      memory[52543] <=  8'h00;      memory[52544] <=  8'h00;      memory[52545] <=  8'h00;      memory[52546] <=  8'h00;      memory[52547] <=  8'h00;      memory[52548] <=  8'h00;      memory[52549] <=  8'h00;      memory[52550] <=  8'h00;      memory[52551] <=  8'h00;      memory[52552] <=  8'h00;      memory[52553] <=  8'h00;      memory[52554] <=  8'h00;      memory[52555] <=  8'h00;      memory[52556] <=  8'h00;      memory[52557] <=  8'h00;      memory[52558] <=  8'h00;      memory[52559] <=  8'h00;      memory[52560] <=  8'h00;      memory[52561] <=  8'h00;      memory[52562] <=  8'h00;      memory[52563] <=  8'h00;      memory[52564] <=  8'h00;      memory[52565] <=  8'h00;      memory[52566] <=  8'h00;      memory[52567] <=  8'h00;      memory[52568] <=  8'h00;      memory[52569] <=  8'h00;      memory[52570] <=  8'h00;      memory[52571] <=  8'h00;      memory[52572] <=  8'h00;      memory[52573] <=  8'h00;      memory[52574] <=  8'h00;      memory[52575] <=  8'h00;      memory[52576] <=  8'h00;      memory[52577] <=  8'h00;      memory[52578] <=  8'h00;      memory[52579] <=  8'h00;      memory[52580] <=  8'h00;      memory[52581] <=  8'h00;      memory[52582] <=  8'h00;      memory[52583] <=  8'h00;      memory[52584] <=  8'h00;      memory[52585] <=  8'h00;      memory[52586] <=  8'h00;      memory[52587] <=  8'h00;      memory[52588] <=  8'h00;      memory[52589] <=  8'h00;      memory[52590] <=  8'h00;      memory[52591] <=  8'h00;      memory[52592] <=  8'h00;      memory[52593] <=  8'h00;      memory[52594] <=  8'h00;      memory[52595] <=  8'h00;      memory[52596] <=  8'h00;      memory[52597] <=  8'h00;      memory[52598] <=  8'h00;      memory[52599] <=  8'h00;      memory[52600] <=  8'h00;      memory[52601] <=  8'h00;      memory[52602] <=  8'h00;      memory[52603] <=  8'h00;      memory[52604] <=  8'h00;      memory[52605] <=  8'h00;      memory[52606] <=  8'h00;      memory[52607] <=  8'h00;      memory[52608] <=  8'h00;      memory[52609] <=  8'h00;      memory[52610] <=  8'h00;      memory[52611] <=  8'h00;      memory[52612] <=  8'h00;      memory[52613] <=  8'h00;      memory[52614] <=  8'h00;      memory[52615] <=  8'h00;      memory[52616] <=  8'h00;      memory[52617] <=  8'h00;      memory[52618] <=  8'h00;      memory[52619] <=  8'h00;      memory[52620] <=  8'h00;      memory[52621] <=  8'h00;      memory[52622] <=  8'h00;      memory[52623] <=  8'h00;      memory[52624] <=  8'h00;      memory[52625] <=  8'h00;      memory[52626] <=  8'h00;      memory[52627] <=  8'h00;      memory[52628] <=  8'h00;      memory[52629] <=  8'h00;      memory[52630] <=  8'h00;      memory[52631] <=  8'h00;      memory[52632] <=  8'h00;      memory[52633] <=  8'h00;      memory[52634] <=  8'h00;      memory[52635] <=  8'h00;      memory[52636] <=  8'h00;      memory[52637] <=  8'h00;      memory[52638] <=  8'h00;      memory[52639] <=  8'h00;      memory[52640] <=  8'h00;      memory[52641] <=  8'h00;      memory[52642] <=  8'h00;      memory[52643] <=  8'h00;      memory[52644] <=  8'h00;      memory[52645] <=  8'h00;      memory[52646] <=  8'h00;      memory[52647] <=  8'h00;      memory[52648] <=  8'h00;      memory[52649] <=  8'h00;      memory[52650] <=  8'h00;      memory[52651] <=  8'h00;      memory[52652] <=  8'h00;      memory[52653] <=  8'h00;      memory[52654] <=  8'h00;      memory[52655] <=  8'h00;      memory[52656] <=  8'h00;      memory[52657] <=  8'h00;      memory[52658] <=  8'h00;      memory[52659] <=  8'h00;      memory[52660] <=  8'h00;      memory[52661] <=  8'h00;      memory[52662] <=  8'h00;      memory[52663] <=  8'h00;      memory[52664] <=  8'h00;      memory[52665] <=  8'h00;      memory[52666] <=  8'h00;      memory[52667] <=  8'h00;      memory[52668] <=  8'h00;      memory[52669] <=  8'h00;      memory[52670] <=  8'h00;      memory[52671] <=  8'h00;      memory[52672] <=  8'h00;      memory[52673] <=  8'h00;      memory[52674] <=  8'h00;      memory[52675] <=  8'h00;      memory[52676] <=  8'h00;      memory[52677] <=  8'h00;      memory[52678] <=  8'h00;      memory[52679] <=  8'h00;      memory[52680] <=  8'h00;      memory[52681] <=  8'h00;      memory[52682] <=  8'h00;      memory[52683] <=  8'h00;      memory[52684] <=  8'h00;      memory[52685] <=  8'h00;      memory[52686] <=  8'h00;      memory[52687] <=  8'h00;      memory[52688] <=  8'h00;      memory[52689] <=  8'h00;      memory[52690] <=  8'h00;      memory[52691] <=  8'h00;      memory[52692] <=  8'h00;      memory[52693] <=  8'h00;      memory[52694] <=  8'h00;      memory[52695] <=  8'h00;      memory[52696] <=  8'h00;      memory[52697] <=  8'h00;      memory[52698] <=  8'h00;      memory[52699] <=  8'h00;      memory[52700] <=  8'h00;      memory[52701] <=  8'h00;      memory[52702] <=  8'h00;      memory[52703] <=  8'h00;      memory[52704] <=  8'h00;      memory[52705] <=  8'h00;      memory[52706] <=  8'h00;      memory[52707] <=  8'h00;      memory[52708] <=  8'h00;      memory[52709] <=  8'h00;      memory[52710] <=  8'h00;      memory[52711] <=  8'h00;      memory[52712] <=  8'h00;      memory[52713] <=  8'h00;      memory[52714] <=  8'h00;      memory[52715] <=  8'h00;      memory[52716] <=  8'h00;      memory[52717] <=  8'h00;      memory[52718] <=  8'h00;      memory[52719] <=  8'h00;      memory[52720] <=  8'h00;      memory[52721] <=  8'h00;      memory[52722] <=  8'h00;      memory[52723] <=  8'h00;      memory[52724] <=  8'h00;      memory[52725] <=  8'h00;      memory[52726] <=  8'h00;      memory[52727] <=  8'h00;      memory[52728] <=  8'h00;      memory[52729] <=  8'h00;      memory[52730] <=  8'h00;      memory[52731] <=  8'h00;      memory[52732] <=  8'h00;      memory[52733] <=  8'h00;      memory[52734] <=  8'h00;      memory[52735] <=  8'h00;      memory[52736] <=  8'h00;      memory[52737] <=  8'h00;      memory[52738] <=  8'h00;      memory[52739] <=  8'h00;      memory[52740] <=  8'h00;      memory[52741] <=  8'h00;      memory[52742] <=  8'h00;      memory[52743] <=  8'h00;      memory[52744] <=  8'h00;      memory[52745] <=  8'h00;      memory[52746] <=  8'h00;      memory[52747] <=  8'h00;      memory[52748] <=  8'h00;      memory[52749] <=  8'h00;      memory[52750] <=  8'h00;      memory[52751] <=  8'h00;      memory[52752] <=  8'h00;      memory[52753] <=  8'h00;      memory[52754] <=  8'h00;      memory[52755] <=  8'h00;      memory[52756] <=  8'h00;      memory[52757] <=  8'h00;      memory[52758] <=  8'h00;      memory[52759] <=  8'h00;      memory[52760] <=  8'h00;      memory[52761] <=  8'h00;      memory[52762] <=  8'h00;      memory[52763] <=  8'h00;      memory[52764] <=  8'h00;      memory[52765] <=  8'h00;      memory[52766] <=  8'h00;      memory[52767] <=  8'h00;      memory[52768] <=  8'h00;      memory[52769] <=  8'h00;      memory[52770] <=  8'h00;      memory[52771] <=  8'h00;      memory[52772] <=  8'h00;      memory[52773] <=  8'h00;      memory[52774] <=  8'h00;      memory[52775] <=  8'h00;      memory[52776] <=  8'h00;      memory[52777] <=  8'h00;      memory[52778] <=  8'h00;      memory[52779] <=  8'h00;      memory[52780] <=  8'h00;      memory[52781] <=  8'h00;      memory[52782] <=  8'h00;      memory[52783] <=  8'h00;      memory[52784] <=  8'h00;      memory[52785] <=  8'h00;      memory[52786] <=  8'h00;      memory[52787] <=  8'h00;      memory[52788] <=  8'h00;      memory[52789] <=  8'h00;      memory[52790] <=  8'h00;      memory[52791] <=  8'h00;      memory[52792] <=  8'h00;      memory[52793] <=  8'h00;      memory[52794] <=  8'h00;      memory[52795] <=  8'h00;      memory[52796] <=  8'h00;      memory[52797] <=  8'h00;      memory[52798] <=  8'h00;      memory[52799] <=  8'h00;      memory[52800] <=  8'h00;      memory[52801] <=  8'h00;      memory[52802] <=  8'h00;      memory[52803] <=  8'h00;      memory[52804] <=  8'h00;      memory[52805] <=  8'h00;      memory[52806] <=  8'h00;      memory[52807] <=  8'h00;      memory[52808] <=  8'h00;      memory[52809] <=  8'h00;      memory[52810] <=  8'h00;      memory[52811] <=  8'h00;      memory[52812] <=  8'h00;      memory[52813] <=  8'h00;      memory[52814] <=  8'h00;      memory[52815] <=  8'h00;      memory[52816] <=  8'h00;      memory[52817] <=  8'h00;      memory[52818] <=  8'h00;      memory[52819] <=  8'h00;      memory[52820] <=  8'h00;      memory[52821] <=  8'h00;      memory[52822] <=  8'h00;      memory[52823] <=  8'h00;      memory[52824] <=  8'h00;      memory[52825] <=  8'h00;      memory[52826] <=  8'h00;      memory[52827] <=  8'h00;      memory[52828] <=  8'h00;      memory[52829] <=  8'h00;      memory[52830] <=  8'h00;      memory[52831] <=  8'h00;      memory[52832] <=  8'h00;      memory[52833] <=  8'h00;      memory[52834] <=  8'h00;      memory[52835] <=  8'h00;      memory[52836] <=  8'h00;      memory[52837] <=  8'h00;      memory[52838] <=  8'h00;      memory[52839] <=  8'h00;      memory[52840] <=  8'h00;      memory[52841] <=  8'h00;      memory[52842] <=  8'h00;      memory[52843] <=  8'h00;      memory[52844] <=  8'h00;      memory[52845] <=  8'h00;      memory[52846] <=  8'h00;      memory[52847] <=  8'h00;      memory[52848] <=  8'h00;      memory[52849] <=  8'h00;      memory[52850] <=  8'h00;      memory[52851] <=  8'h00;      memory[52852] <=  8'h00;      memory[52853] <=  8'h00;      memory[52854] <=  8'h00;      memory[52855] <=  8'h00;      memory[52856] <=  8'h00;      memory[52857] <=  8'h00;      memory[52858] <=  8'h00;      memory[52859] <=  8'h00;      memory[52860] <=  8'h00;      memory[52861] <=  8'h00;      memory[52862] <=  8'h00;      memory[52863] <=  8'h00;      memory[52864] <=  8'h00;      memory[52865] <=  8'h00;      memory[52866] <=  8'h00;      memory[52867] <=  8'h00;      memory[52868] <=  8'h00;      memory[52869] <=  8'h00;      memory[52870] <=  8'h00;      memory[52871] <=  8'h00;      memory[52872] <=  8'h00;      memory[52873] <=  8'h00;      memory[52874] <=  8'h00;      memory[52875] <=  8'h00;      memory[52876] <=  8'h00;      memory[52877] <=  8'h00;      memory[52878] <=  8'h00;      memory[52879] <=  8'h00;      memory[52880] <=  8'h00;      memory[52881] <=  8'h00;      memory[52882] <=  8'h00;      memory[52883] <=  8'h00;      memory[52884] <=  8'h00;      memory[52885] <=  8'h00;      memory[52886] <=  8'h00;      memory[52887] <=  8'h00;      memory[52888] <=  8'h00;      memory[52889] <=  8'h00;      memory[52890] <=  8'h00;      memory[52891] <=  8'h00;      memory[52892] <=  8'h00;      memory[52893] <=  8'h00;      memory[52894] <=  8'h00;      memory[52895] <=  8'h00;      memory[52896] <=  8'h00;      memory[52897] <=  8'h00;      memory[52898] <=  8'h00;      memory[52899] <=  8'h00;      memory[52900] <=  8'h00;      memory[52901] <=  8'h00;      memory[52902] <=  8'h00;      memory[52903] <=  8'h00;      memory[52904] <=  8'h00;      memory[52905] <=  8'h00;      memory[52906] <=  8'h00;      memory[52907] <=  8'h00;      memory[52908] <=  8'h00;      memory[52909] <=  8'h00;      memory[52910] <=  8'h00;      memory[52911] <=  8'h00;      memory[52912] <=  8'h00;      memory[52913] <=  8'h00;      memory[52914] <=  8'h00;      memory[52915] <=  8'h00;      memory[52916] <=  8'h00;      memory[52917] <=  8'h00;      memory[52918] <=  8'h00;      memory[52919] <=  8'h00;      memory[52920] <=  8'h00;      memory[52921] <=  8'h00;      memory[52922] <=  8'h00;      memory[52923] <=  8'h00;      memory[52924] <=  8'h00;      memory[52925] <=  8'h00;      memory[52926] <=  8'h00;      memory[52927] <=  8'h00;      memory[52928] <=  8'h00;      memory[52929] <=  8'h00;      memory[52930] <=  8'h00;      memory[52931] <=  8'h00;      memory[52932] <=  8'h00;      memory[52933] <=  8'h00;      memory[52934] <=  8'h00;      memory[52935] <=  8'h00;      memory[52936] <=  8'h00;      memory[52937] <=  8'h00;      memory[52938] <=  8'h00;      memory[52939] <=  8'h00;      memory[52940] <=  8'h00;      memory[52941] <=  8'h00;      memory[52942] <=  8'h00;      memory[52943] <=  8'h00;      memory[52944] <=  8'h00;      memory[52945] <=  8'h00;      memory[52946] <=  8'h00;      memory[52947] <=  8'h00;      memory[52948] <=  8'h00;      memory[52949] <=  8'h00;      memory[52950] <=  8'h00;      memory[52951] <=  8'h00;      memory[52952] <=  8'h00;      memory[52953] <=  8'h00;      memory[52954] <=  8'h00;      memory[52955] <=  8'h00;      memory[52956] <=  8'h00;      memory[52957] <=  8'h00;      memory[52958] <=  8'h00;      memory[52959] <=  8'h00;      memory[52960] <=  8'h00;      memory[52961] <=  8'h00;      memory[52962] <=  8'h00;      memory[52963] <=  8'h00;      memory[52964] <=  8'h00;      memory[52965] <=  8'h00;      memory[52966] <=  8'h00;      memory[52967] <=  8'h00;      memory[52968] <=  8'h00;      memory[52969] <=  8'h00;      memory[52970] <=  8'h00;      memory[52971] <=  8'h00;      memory[52972] <=  8'h00;      memory[52973] <=  8'h00;      memory[52974] <=  8'h00;      memory[52975] <=  8'h00;      memory[52976] <=  8'h00;      memory[52977] <=  8'h00;      memory[52978] <=  8'h00;      memory[52979] <=  8'h00;      memory[52980] <=  8'h00;      memory[52981] <=  8'h00;      memory[52982] <=  8'h00;      memory[52983] <=  8'h00;      memory[52984] <=  8'h00;      memory[52985] <=  8'h00;      memory[52986] <=  8'h00;      memory[52987] <=  8'h00;      memory[52988] <=  8'h00;      memory[52989] <=  8'h00;      memory[52990] <=  8'h00;      memory[52991] <=  8'h00;      memory[52992] <=  8'h00;      memory[52993] <=  8'h00;      memory[52994] <=  8'h00;      memory[52995] <=  8'h00;      memory[52996] <=  8'h00;      memory[52997] <=  8'h00;      memory[52998] <=  8'h00;      memory[52999] <=  8'h00;      memory[53000] <=  8'h00;      memory[53001] <=  8'h00;      memory[53002] <=  8'h00;      memory[53003] <=  8'h00;      memory[53004] <=  8'h00;      memory[53005] <=  8'h00;      memory[53006] <=  8'h00;      memory[53007] <=  8'h00;      memory[53008] <=  8'h00;      memory[53009] <=  8'h00;      memory[53010] <=  8'h00;      memory[53011] <=  8'h00;      memory[53012] <=  8'h00;      memory[53013] <=  8'h00;      memory[53014] <=  8'h00;      memory[53015] <=  8'h00;      memory[53016] <=  8'h00;      memory[53017] <=  8'h00;      memory[53018] <=  8'h00;      memory[53019] <=  8'h00;      memory[53020] <=  8'h00;      memory[53021] <=  8'h00;      memory[53022] <=  8'h00;      memory[53023] <=  8'h00;      memory[53024] <=  8'h00;      memory[53025] <=  8'h00;      memory[53026] <=  8'h00;      memory[53027] <=  8'h00;      memory[53028] <=  8'h00;      memory[53029] <=  8'h00;      memory[53030] <=  8'h00;      memory[53031] <=  8'h00;      memory[53032] <=  8'h00;      memory[53033] <=  8'h00;      memory[53034] <=  8'h00;      memory[53035] <=  8'h00;      memory[53036] <=  8'h00;      memory[53037] <=  8'h00;      memory[53038] <=  8'h00;      memory[53039] <=  8'h00;      memory[53040] <=  8'h00;      memory[53041] <=  8'h00;      memory[53042] <=  8'h00;      memory[53043] <=  8'h00;      memory[53044] <=  8'h00;      memory[53045] <=  8'h00;      memory[53046] <=  8'h00;      memory[53047] <=  8'h00;      memory[53048] <=  8'h00;      memory[53049] <=  8'h00;      memory[53050] <=  8'h00;      memory[53051] <=  8'h00;      memory[53052] <=  8'h00;      memory[53053] <=  8'h00;      memory[53054] <=  8'h00;      memory[53055] <=  8'h00;      memory[53056] <=  8'h00;      memory[53057] <=  8'h00;      memory[53058] <=  8'h00;      memory[53059] <=  8'h00;      memory[53060] <=  8'h00;      memory[53061] <=  8'h00;      memory[53062] <=  8'h00;      memory[53063] <=  8'h00;      memory[53064] <=  8'h00;      memory[53065] <=  8'h00;      memory[53066] <=  8'h00;      memory[53067] <=  8'h00;      memory[53068] <=  8'h00;      memory[53069] <=  8'h00;      memory[53070] <=  8'h00;      memory[53071] <=  8'h00;      memory[53072] <=  8'h00;      memory[53073] <=  8'h00;      memory[53074] <=  8'h00;      memory[53075] <=  8'h00;      memory[53076] <=  8'h00;      memory[53077] <=  8'h00;      memory[53078] <=  8'h00;      memory[53079] <=  8'h00;      memory[53080] <=  8'h00;      memory[53081] <=  8'h00;      memory[53082] <=  8'h00;      memory[53083] <=  8'h00;      memory[53084] <=  8'h00;      memory[53085] <=  8'h00;      memory[53086] <=  8'h00;      memory[53087] <=  8'h00;      memory[53088] <=  8'h00;      memory[53089] <=  8'h00;      memory[53090] <=  8'h00;      memory[53091] <=  8'h00;      memory[53092] <=  8'h00;      memory[53093] <=  8'h00;      memory[53094] <=  8'h00;      memory[53095] <=  8'h00;      memory[53096] <=  8'h00;      memory[53097] <=  8'h00;      memory[53098] <=  8'h00;      memory[53099] <=  8'h00;      memory[53100] <=  8'h00;      memory[53101] <=  8'h00;      memory[53102] <=  8'h00;      memory[53103] <=  8'h00;      memory[53104] <=  8'h00;      memory[53105] <=  8'h00;      memory[53106] <=  8'h00;      memory[53107] <=  8'h00;      memory[53108] <=  8'h00;      memory[53109] <=  8'h00;      memory[53110] <=  8'h00;      memory[53111] <=  8'h00;      memory[53112] <=  8'h00;      memory[53113] <=  8'h00;      memory[53114] <=  8'h00;      memory[53115] <=  8'h00;      memory[53116] <=  8'h00;      memory[53117] <=  8'h00;      memory[53118] <=  8'h00;      memory[53119] <=  8'h00;      memory[53120] <=  8'h00;      memory[53121] <=  8'h00;      memory[53122] <=  8'h00;      memory[53123] <=  8'h00;      memory[53124] <=  8'h00;      memory[53125] <=  8'h00;      memory[53126] <=  8'h00;      memory[53127] <=  8'h00;      memory[53128] <=  8'h00;      memory[53129] <=  8'h00;      memory[53130] <=  8'h00;      memory[53131] <=  8'h00;      memory[53132] <=  8'h00;      memory[53133] <=  8'h00;      memory[53134] <=  8'h00;      memory[53135] <=  8'h00;      memory[53136] <=  8'h00;      memory[53137] <=  8'h00;      memory[53138] <=  8'h00;      memory[53139] <=  8'h00;      memory[53140] <=  8'h00;      memory[53141] <=  8'h00;      memory[53142] <=  8'h00;      memory[53143] <=  8'h00;      memory[53144] <=  8'h00;      memory[53145] <=  8'h00;      memory[53146] <=  8'h00;      memory[53147] <=  8'h00;      memory[53148] <=  8'h00;      memory[53149] <=  8'h00;      memory[53150] <=  8'h00;      memory[53151] <=  8'h00;      memory[53152] <=  8'h00;      memory[53153] <=  8'h00;      memory[53154] <=  8'h00;      memory[53155] <=  8'h00;      memory[53156] <=  8'h00;      memory[53157] <=  8'h00;      memory[53158] <=  8'h00;      memory[53159] <=  8'h00;      memory[53160] <=  8'h00;      memory[53161] <=  8'h00;      memory[53162] <=  8'h00;      memory[53163] <=  8'h00;      memory[53164] <=  8'h00;      memory[53165] <=  8'h00;      memory[53166] <=  8'h00;      memory[53167] <=  8'h00;      memory[53168] <=  8'h00;      memory[53169] <=  8'h00;      memory[53170] <=  8'h00;      memory[53171] <=  8'h00;      memory[53172] <=  8'h00;      memory[53173] <=  8'h00;      memory[53174] <=  8'h00;      memory[53175] <=  8'h00;      memory[53176] <=  8'h00;      memory[53177] <=  8'h00;      memory[53178] <=  8'h00;      memory[53179] <=  8'h00;      memory[53180] <=  8'h00;      memory[53181] <=  8'h00;      memory[53182] <=  8'h00;      memory[53183] <=  8'h00;      memory[53184] <=  8'h00;      memory[53185] <=  8'h00;      memory[53186] <=  8'h00;      memory[53187] <=  8'h00;      memory[53188] <=  8'h00;      memory[53189] <=  8'h00;      memory[53190] <=  8'h00;      memory[53191] <=  8'h00;      memory[53192] <=  8'h00;      memory[53193] <=  8'h00;      memory[53194] <=  8'h00;      memory[53195] <=  8'h00;      memory[53196] <=  8'h00;      memory[53197] <=  8'h00;      memory[53198] <=  8'h00;      memory[53199] <=  8'h00;      memory[53200] <=  8'h00;      memory[53201] <=  8'h00;      memory[53202] <=  8'h00;      memory[53203] <=  8'h00;      memory[53204] <=  8'h00;      memory[53205] <=  8'h00;      memory[53206] <=  8'h00;      memory[53207] <=  8'h00;      memory[53208] <=  8'h00;      memory[53209] <=  8'h00;      memory[53210] <=  8'h00;      memory[53211] <=  8'h00;      memory[53212] <=  8'h00;      memory[53213] <=  8'h00;      memory[53214] <=  8'h00;      memory[53215] <=  8'h00;      memory[53216] <=  8'h00;      memory[53217] <=  8'h00;      memory[53218] <=  8'h00;      memory[53219] <=  8'h00;      memory[53220] <=  8'h00;      memory[53221] <=  8'h00;      memory[53222] <=  8'h00;      memory[53223] <=  8'h00;      memory[53224] <=  8'h00;      memory[53225] <=  8'h00;      memory[53226] <=  8'h00;      memory[53227] <=  8'h00;      memory[53228] <=  8'h00;      memory[53229] <=  8'h00;      memory[53230] <=  8'h00;      memory[53231] <=  8'h00;      memory[53232] <=  8'h00;      memory[53233] <=  8'h00;      memory[53234] <=  8'h00;      memory[53235] <=  8'h00;      memory[53236] <=  8'h00;      memory[53237] <=  8'h00;      memory[53238] <=  8'h00;      memory[53239] <=  8'h00;      memory[53240] <=  8'h00;      memory[53241] <=  8'h00;      memory[53242] <=  8'h00;      memory[53243] <=  8'h00;      memory[53244] <=  8'h00;      memory[53245] <=  8'h00;      memory[53246] <=  8'h00;      memory[53247] <=  8'h00;      memory[53248] <=  8'h00;      memory[53249] <=  8'h00;      memory[53250] <=  8'h00;      memory[53251] <=  8'h00;      memory[53252] <=  8'h00;      memory[53253] <=  8'h00;      memory[53254] <=  8'h00;      memory[53255] <=  8'h00;      memory[53256] <=  8'h00;      memory[53257] <=  8'h00;      memory[53258] <=  8'h00;      memory[53259] <=  8'h00;      memory[53260] <=  8'h00;      memory[53261] <=  8'h00;      memory[53262] <=  8'h00;      memory[53263] <=  8'h00;      memory[53264] <=  8'h00;      memory[53265] <=  8'h00;      memory[53266] <=  8'h00;      memory[53267] <=  8'h00;      memory[53268] <=  8'h00;      memory[53269] <=  8'h00;      memory[53270] <=  8'h00;      memory[53271] <=  8'h00;      memory[53272] <=  8'h00;      memory[53273] <=  8'h00;      memory[53274] <=  8'h00;      memory[53275] <=  8'h00;      memory[53276] <=  8'h00;      memory[53277] <=  8'h00;      memory[53278] <=  8'h00;      memory[53279] <=  8'h00;      memory[53280] <=  8'h00;      memory[53281] <=  8'h00;      memory[53282] <=  8'h00;      memory[53283] <=  8'h00;      memory[53284] <=  8'h00;      memory[53285] <=  8'h00;      memory[53286] <=  8'h00;      memory[53287] <=  8'h00;      memory[53288] <=  8'h00;      memory[53289] <=  8'h00;      memory[53290] <=  8'h00;      memory[53291] <=  8'h00;      memory[53292] <=  8'h00;      memory[53293] <=  8'h00;      memory[53294] <=  8'h00;      memory[53295] <=  8'h00;      memory[53296] <=  8'h00;      memory[53297] <=  8'h00;      memory[53298] <=  8'h00;      memory[53299] <=  8'h00;      memory[53300] <=  8'h00;      memory[53301] <=  8'h00;      memory[53302] <=  8'h00;      memory[53303] <=  8'h00;      memory[53304] <=  8'h00;      memory[53305] <=  8'h00;      memory[53306] <=  8'h00;      memory[53307] <=  8'h00;      memory[53308] <=  8'h00;      memory[53309] <=  8'h00;      memory[53310] <=  8'h00;      memory[53311] <=  8'h00;      memory[53312] <=  8'h00;      memory[53313] <=  8'h00;      memory[53314] <=  8'h00;      memory[53315] <=  8'h00;      memory[53316] <=  8'h00;      memory[53317] <=  8'h00;      memory[53318] <=  8'h00;      memory[53319] <=  8'h00;      memory[53320] <=  8'h00;      memory[53321] <=  8'h00;      memory[53322] <=  8'h00;      memory[53323] <=  8'h00;      memory[53324] <=  8'h00;      memory[53325] <=  8'h00;      memory[53326] <=  8'h00;      memory[53327] <=  8'h00;      memory[53328] <=  8'h00;      memory[53329] <=  8'h00;      memory[53330] <=  8'h00;      memory[53331] <=  8'h00;      memory[53332] <=  8'h00;      memory[53333] <=  8'h00;      memory[53334] <=  8'h00;      memory[53335] <=  8'h00;      memory[53336] <=  8'h00;      memory[53337] <=  8'h00;      memory[53338] <=  8'h00;      memory[53339] <=  8'h00;      memory[53340] <=  8'h00;      memory[53341] <=  8'h00;      memory[53342] <=  8'h00;      memory[53343] <=  8'h00;      memory[53344] <=  8'h00;      memory[53345] <=  8'h00;      memory[53346] <=  8'h00;      memory[53347] <=  8'h00;      memory[53348] <=  8'h00;      memory[53349] <=  8'h00;      memory[53350] <=  8'h00;      memory[53351] <=  8'h00;      memory[53352] <=  8'h00;      memory[53353] <=  8'h00;      memory[53354] <=  8'h00;      memory[53355] <=  8'h00;      memory[53356] <=  8'h00;      memory[53357] <=  8'h00;      memory[53358] <=  8'h00;      memory[53359] <=  8'h00;      memory[53360] <=  8'h00;      memory[53361] <=  8'h00;      memory[53362] <=  8'h00;      memory[53363] <=  8'h00;      memory[53364] <=  8'h00;      memory[53365] <=  8'h00;      memory[53366] <=  8'h00;      memory[53367] <=  8'h00;      memory[53368] <=  8'h00;      memory[53369] <=  8'h00;      memory[53370] <=  8'h00;      memory[53371] <=  8'h00;      memory[53372] <=  8'h00;      memory[53373] <=  8'h00;      memory[53374] <=  8'h00;      memory[53375] <=  8'h00;      memory[53376] <=  8'h00;      memory[53377] <=  8'h00;      memory[53378] <=  8'h00;      memory[53379] <=  8'h00;      memory[53380] <=  8'h00;      memory[53381] <=  8'h00;      memory[53382] <=  8'h00;      memory[53383] <=  8'h00;      memory[53384] <=  8'h00;      memory[53385] <=  8'h00;      memory[53386] <=  8'h00;      memory[53387] <=  8'h00;      memory[53388] <=  8'h00;      memory[53389] <=  8'h00;      memory[53390] <=  8'h00;      memory[53391] <=  8'h00;      memory[53392] <=  8'h00;      memory[53393] <=  8'h00;      memory[53394] <=  8'h00;      memory[53395] <=  8'h00;      memory[53396] <=  8'h00;      memory[53397] <=  8'h00;      memory[53398] <=  8'h00;      memory[53399] <=  8'h00;      memory[53400] <=  8'h00;      memory[53401] <=  8'h00;      memory[53402] <=  8'h00;      memory[53403] <=  8'h00;      memory[53404] <=  8'h00;      memory[53405] <=  8'h00;      memory[53406] <=  8'h00;      memory[53407] <=  8'h00;      memory[53408] <=  8'h00;      memory[53409] <=  8'h00;      memory[53410] <=  8'h00;      memory[53411] <=  8'h00;      memory[53412] <=  8'h00;      memory[53413] <=  8'h00;      memory[53414] <=  8'h00;      memory[53415] <=  8'h00;      memory[53416] <=  8'h00;      memory[53417] <=  8'h00;      memory[53418] <=  8'h00;      memory[53419] <=  8'h00;      memory[53420] <=  8'h00;      memory[53421] <=  8'h00;      memory[53422] <=  8'h00;      memory[53423] <=  8'h00;      memory[53424] <=  8'h00;      memory[53425] <=  8'h00;      memory[53426] <=  8'h00;      memory[53427] <=  8'h00;      memory[53428] <=  8'h00;      memory[53429] <=  8'h00;      memory[53430] <=  8'h00;      memory[53431] <=  8'h00;      memory[53432] <=  8'h00;      memory[53433] <=  8'h00;      memory[53434] <=  8'h00;      memory[53435] <=  8'h00;      memory[53436] <=  8'h00;      memory[53437] <=  8'h00;      memory[53438] <=  8'h00;      memory[53439] <=  8'h00;      memory[53440] <=  8'h00;      memory[53441] <=  8'h00;      memory[53442] <=  8'h00;      memory[53443] <=  8'h00;      memory[53444] <=  8'h00;      memory[53445] <=  8'h00;      memory[53446] <=  8'h00;      memory[53447] <=  8'h00;      memory[53448] <=  8'h00;      memory[53449] <=  8'h00;      memory[53450] <=  8'h00;      memory[53451] <=  8'h00;      memory[53452] <=  8'h00;      memory[53453] <=  8'h00;      memory[53454] <=  8'h00;      memory[53455] <=  8'h00;      memory[53456] <=  8'h00;      memory[53457] <=  8'h00;      memory[53458] <=  8'h00;      memory[53459] <=  8'h00;      memory[53460] <=  8'h00;      memory[53461] <=  8'h00;      memory[53462] <=  8'h00;      memory[53463] <=  8'h00;      memory[53464] <=  8'h00;      memory[53465] <=  8'h00;      memory[53466] <=  8'h00;      memory[53467] <=  8'h00;      memory[53468] <=  8'h00;      memory[53469] <=  8'h00;      memory[53470] <=  8'h00;      memory[53471] <=  8'h00;      memory[53472] <=  8'h00;      memory[53473] <=  8'h00;      memory[53474] <=  8'h00;      memory[53475] <=  8'h00;      memory[53476] <=  8'h00;      memory[53477] <=  8'h00;      memory[53478] <=  8'h00;      memory[53479] <=  8'h00;      memory[53480] <=  8'h00;      memory[53481] <=  8'h00;      memory[53482] <=  8'h00;      memory[53483] <=  8'h00;      memory[53484] <=  8'h00;      memory[53485] <=  8'h00;      memory[53486] <=  8'h00;      memory[53487] <=  8'h00;      memory[53488] <=  8'h00;      memory[53489] <=  8'h00;      memory[53490] <=  8'h00;      memory[53491] <=  8'h00;      memory[53492] <=  8'h00;      memory[53493] <=  8'h00;      memory[53494] <=  8'h00;      memory[53495] <=  8'h00;      memory[53496] <=  8'h00;      memory[53497] <=  8'h00;      memory[53498] <=  8'h00;      memory[53499] <=  8'h00;      memory[53500] <=  8'h00;      memory[53501] <=  8'h00;      memory[53502] <=  8'h00;      memory[53503] <=  8'h00;      memory[53504] <=  8'h00;      memory[53505] <=  8'h00;      memory[53506] <=  8'h00;      memory[53507] <=  8'h00;      memory[53508] <=  8'h00;      memory[53509] <=  8'h00;      memory[53510] <=  8'h00;      memory[53511] <=  8'h00;      memory[53512] <=  8'h00;      memory[53513] <=  8'h00;      memory[53514] <=  8'h00;      memory[53515] <=  8'h00;      memory[53516] <=  8'h00;      memory[53517] <=  8'h00;      memory[53518] <=  8'h00;      memory[53519] <=  8'h00;      memory[53520] <=  8'h00;      memory[53521] <=  8'h00;      memory[53522] <=  8'h00;      memory[53523] <=  8'h00;      memory[53524] <=  8'h00;      memory[53525] <=  8'h00;      memory[53526] <=  8'h00;      memory[53527] <=  8'h00;      memory[53528] <=  8'h00;      memory[53529] <=  8'h00;      memory[53530] <=  8'h00;      memory[53531] <=  8'h00;      memory[53532] <=  8'h00;      memory[53533] <=  8'h00;      memory[53534] <=  8'h00;      memory[53535] <=  8'h00;      memory[53536] <=  8'h00;      memory[53537] <=  8'h00;      memory[53538] <=  8'h00;      memory[53539] <=  8'h00;      memory[53540] <=  8'h00;      memory[53541] <=  8'h00;      memory[53542] <=  8'h00;      memory[53543] <=  8'h00;      memory[53544] <=  8'h00;      memory[53545] <=  8'h00;      memory[53546] <=  8'h00;      memory[53547] <=  8'h00;      memory[53548] <=  8'h00;      memory[53549] <=  8'h00;      memory[53550] <=  8'h00;      memory[53551] <=  8'h00;      memory[53552] <=  8'h00;      memory[53553] <=  8'h00;      memory[53554] <=  8'h00;      memory[53555] <=  8'h00;      memory[53556] <=  8'h00;      memory[53557] <=  8'h00;      memory[53558] <=  8'h00;      memory[53559] <=  8'h00;      memory[53560] <=  8'h00;      memory[53561] <=  8'h00;      memory[53562] <=  8'h00;      memory[53563] <=  8'h00;      memory[53564] <=  8'h00;      memory[53565] <=  8'h00;      memory[53566] <=  8'h00;      memory[53567] <=  8'h00;      memory[53568] <=  8'h00;      memory[53569] <=  8'h00;      memory[53570] <=  8'h00;      memory[53571] <=  8'h00;      memory[53572] <=  8'h00;      memory[53573] <=  8'h00;      memory[53574] <=  8'h00;      memory[53575] <=  8'h00;      memory[53576] <=  8'h00;      memory[53577] <=  8'h00;      memory[53578] <=  8'h00;      memory[53579] <=  8'h00;      memory[53580] <=  8'h00;      memory[53581] <=  8'h00;      memory[53582] <=  8'h00;      memory[53583] <=  8'h00;      memory[53584] <=  8'h00;      memory[53585] <=  8'h00;      memory[53586] <=  8'h00;      memory[53587] <=  8'h00;      memory[53588] <=  8'h00;      memory[53589] <=  8'h00;      memory[53590] <=  8'h00;      memory[53591] <=  8'h00;      memory[53592] <=  8'h00;      memory[53593] <=  8'h00;      memory[53594] <=  8'h00;      memory[53595] <=  8'h00;      memory[53596] <=  8'h00;      memory[53597] <=  8'h00;      memory[53598] <=  8'h00;      memory[53599] <=  8'h00;      memory[53600] <=  8'h00;      memory[53601] <=  8'h00;      memory[53602] <=  8'h00;      memory[53603] <=  8'h00;      memory[53604] <=  8'h00;      memory[53605] <=  8'h00;      memory[53606] <=  8'h00;      memory[53607] <=  8'h00;      memory[53608] <=  8'h00;      memory[53609] <=  8'h00;      memory[53610] <=  8'h00;      memory[53611] <=  8'h00;      memory[53612] <=  8'h00;      memory[53613] <=  8'h00;      memory[53614] <=  8'h00;      memory[53615] <=  8'h00;      memory[53616] <=  8'h00;      memory[53617] <=  8'h00;      memory[53618] <=  8'h00;      memory[53619] <=  8'h00;      memory[53620] <=  8'h00;      memory[53621] <=  8'h00;      memory[53622] <=  8'h00;      memory[53623] <=  8'h00;      memory[53624] <=  8'h00;      memory[53625] <=  8'h00;      memory[53626] <=  8'h00;      memory[53627] <=  8'h00;      memory[53628] <=  8'h00;      memory[53629] <=  8'h00;      memory[53630] <=  8'h00;      memory[53631] <=  8'h00;      memory[53632] <=  8'h00;      memory[53633] <=  8'h00;      memory[53634] <=  8'h00;      memory[53635] <=  8'h00;      memory[53636] <=  8'h00;      memory[53637] <=  8'h00;      memory[53638] <=  8'h00;      memory[53639] <=  8'h00;      memory[53640] <=  8'h00;      memory[53641] <=  8'h00;      memory[53642] <=  8'h00;      memory[53643] <=  8'h00;      memory[53644] <=  8'h00;      memory[53645] <=  8'h00;      memory[53646] <=  8'h00;      memory[53647] <=  8'h00;      memory[53648] <=  8'h00;      memory[53649] <=  8'h00;      memory[53650] <=  8'h00;      memory[53651] <=  8'h00;      memory[53652] <=  8'h00;      memory[53653] <=  8'h00;      memory[53654] <=  8'h00;      memory[53655] <=  8'h00;      memory[53656] <=  8'h00;      memory[53657] <=  8'h00;      memory[53658] <=  8'h00;      memory[53659] <=  8'h00;      memory[53660] <=  8'h00;      memory[53661] <=  8'h00;      memory[53662] <=  8'h00;      memory[53663] <=  8'h00;      memory[53664] <=  8'h00;      memory[53665] <=  8'h00;      memory[53666] <=  8'h00;      memory[53667] <=  8'h00;      memory[53668] <=  8'h00;      memory[53669] <=  8'h00;      memory[53670] <=  8'h00;      memory[53671] <=  8'h00;      memory[53672] <=  8'h00;      memory[53673] <=  8'h00;      memory[53674] <=  8'h00;      memory[53675] <=  8'h00;      memory[53676] <=  8'h00;      memory[53677] <=  8'h00;      memory[53678] <=  8'h00;      memory[53679] <=  8'h00;      memory[53680] <=  8'h00;      memory[53681] <=  8'h00;      memory[53682] <=  8'h00;      memory[53683] <=  8'h00;      memory[53684] <=  8'h00;      memory[53685] <=  8'h00;      memory[53686] <=  8'h00;      memory[53687] <=  8'h00;      memory[53688] <=  8'h00;      memory[53689] <=  8'h00;      memory[53690] <=  8'h00;      memory[53691] <=  8'h00;      memory[53692] <=  8'h00;      memory[53693] <=  8'h00;      memory[53694] <=  8'h00;      memory[53695] <=  8'h00;      memory[53696] <=  8'h00;      memory[53697] <=  8'h00;      memory[53698] <=  8'h00;      memory[53699] <=  8'h00;      memory[53700] <=  8'h00;      memory[53701] <=  8'h00;      memory[53702] <=  8'h00;      memory[53703] <=  8'h00;      memory[53704] <=  8'h00;      memory[53705] <=  8'h00;      memory[53706] <=  8'h00;      memory[53707] <=  8'h00;      memory[53708] <=  8'h00;      memory[53709] <=  8'h00;      memory[53710] <=  8'h00;      memory[53711] <=  8'h00;      memory[53712] <=  8'h00;      memory[53713] <=  8'h00;      memory[53714] <=  8'h00;      memory[53715] <=  8'h00;      memory[53716] <=  8'h00;      memory[53717] <=  8'h00;      memory[53718] <=  8'h00;      memory[53719] <=  8'h00;      memory[53720] <=  8'h00;      memory[53721] <=  8'h00;      memory[53722] <=  8'h00;      memory[53723] <=  8'h00;      memory[53724] <=  8'h00;      memory[53725] <=  8'h00;      memory[53726] <=  8'h00;      memory[53727] <=  8'h00;      memory[53728] <=  8'h00;      memory[53729] <=  8'h00;      memory[53730] <=  8'h00;      memory[53731] <=  8'h00;      memory[53732] <=  8'h00;      memory[53733] <=  8'h00;      memory[53734] <=  8'h00;      memory[53735] <=  8'h00;      memory[53736] <=  8'h00;      memory[53737] <=  8'h00;      memory[53738] <=  8'h00;      memory[53739] <=  8'h00;      memory[53740] <=  8'h00;      memory[53741] <=  8'h00;      memory[53742] <=  8'h00;      memory[53743] <=  8'h00;      memory[53744] <=  8'h00;      memory[53745] <=  8'h00;      memory[53746] <=  8'h00;      memory[53747] <=  8'h00;      memory[53748] <=  8'h00;      memory[53749] <=  8'h00;      memory[53750] <=  8'h00;      memory[53751] <=  8'h00;      memory[53752] <=  8'h00;      memory[53753] <=  8'h00;      memory[53754] <=  8'h00;      memory[53755] <=  8'h00;      memory[53756] <=  8'h00;      memory[53757] <=  8'h00;      memory[53758] <=  8'h00;      memory[53759] <=  8'h00;      memory[53760] <=  8'h00;      memory[53761] <=  8'h00;      memory[53762] <=  8'h00;      memory[53763] <=  8'h00;      memory[53764] <=  8'h00;      memory[53765] <=  8'h00;      memory[53766] <=  8'h00;      memory[53767] <=  8'h00;      memory[53768] <=  8'h00;      memory[53769] <=  8'h00;      memory[53770] <=  8'h00;      memory[53771] <=  8'h00;      memory[53772] <=  8'h00;      memory[53773] <=  8'h00;      memory[53774] <=  8'h00;      memory[53775] <=  8'h00;      memory[53776] <=  8'h00;      memory[53777] <=  8'h00;      memory[53778] <=  8'h00;      memory[53779] <=  8'h00;      memory[53780] <=  8'h00;      memory[53781] <=  8'h00;      memory[53782] <=  8'h00;      memory[53783] <=  8'h00;      memory[53784] <=  8'h00;      memory[53785] <=  8'h00;      memory[53786] <=  8'h00;      memory[53787] <=  8'h00;      memory[53788] <=  8'h00;      memory[53789] <=  8'h00;      memory[53790] <=  8'h00;      memory[53791] <=  8'h00;      memory[53792] <=  8'h00;      memory[53793] <=  8'h00;      memory[53794] <=  8'h00;      memory[53795] <=  8'h00;      memory[53796] <=  8'h00;      memory[53797] <=  8'h00;      memory[53798] <=  8'h00;      memory[53799] <=  8'h00;      memory[53800] <=  8'h00;      memory[53801] <=  8'h00;      memory[53802] <=  8'h00;      memory[53803] <=  8'h00;      memory[53804] <=  8'h00;      memory[53805] <=  8'h00;      memory[53806] <=  8'h00;      memory[53807] <=  8'h00;      memory[53808] <=  8'h00;      memory[53809] <=  8'h00;      memory[53810] <=  8'h00;      memory[53811] <=  8'h00;      memory[53812] <=  8'h00;      memory[53813] <=  8'h00;      memory[53814] <=  8'h00;      memory[53815] <=  8'h00;      memory[53816] <=  8'h00;      memory[53817] <=  8'h00;      memory[53818] <=  8'h00;      memory[53819] <=  8'h00;      memory[53820] <=  8'h00;      memory[53821] <=  8'h00;      memory[53822] <=  8'h00;      memory[53823] <=  8'h00;      memory[53824] <=  8'h00;      memory[53825] <=  8'h00;      memory[53826] <=  8'h00;      memory[53827] <=  8'h00;      memory[53828] <=  8'h00;      memory[53829] <=  8'h00;      memory[53830] <=  8'h00;      memory[53831] <=  8'h00;      memory[53832] <=  8'h00;      memory[53833] <=  8'h00;      memory[53834] <=  8'h00;      memory[53835] <=  8'h00;      memory[53836] <=  8'h00;      memory[53837] <=  8'h00;      memory[53838] <=  8'h00;      memory[53839] <=  8'h00;      memory[53840] <=  8'h00;      memory[53841] <=  8'h00;      memory[53842] <=  8'h00;      memory[53843] <=  8'h00;      memory[53844] <=  8'h00;      memory[53845] <=  8'h00;      memory[53846] <=  8'h00;      memory[53847] <=  8'h00;      memory[53848] <=  8'h00;      memory[53849] <=  8'h00;      memory[53850] <=  8'h00;      memory[53851] <=  8'h00;      memory[53852] <=  8'h00;      memory[53853] <=  8'h00;      memory[53854] <=  8'h00;      memory[53855] <=  8'h00;      memory[53856] <=  8'h00;      memory[53857] <=  8'h00;      memory[53858] <=  8'h00;      memory[53859] <=  8'h00;      memory[53860] <=  8'h00;      memory[53861] <=  8'h00;      memory[53862] <=  8'h00;      memory[53863] <=  8'h00;      memory[53864] <=  8'h00;      memory[53865] <=  8'h00;      memory[53866] <=  8'h00;      memory[53867] <=  8'h00;      memory[53868] <=  8'h00;      memory[53869] <=  8'h00;      memory[53870] <=  8'h00;      memory[53871] <=  8'h00;      memory[53872] <=  8'h00;      memory[53873] <=  8'h00;      memory[53874] <=  8'h00;      memory[53875] <=  8'h00;      memory[53876] <=  8'h00;      memory[53877] <=  8'h00;      memory[53878] <=  8'h00;      memory[53879] <=  8'h00;      memory[53880] <=  8'h00;      memory[53881] <=  8'h00;      memory[53882] <=  8'h00;      memory[53883] <=  8'h00;      memory[53884] <=  8'h00;      memory[53885] <=  8'h00;      memory[53886] <=  8'h00;      memory[53887] <=  8'h00;      memory[53888] <=  8'h00;      memory[53889] <=  8'h00;      memory[53890] <=  8'h00;      memory[53891] <=  8'h00;      memory[53892] <=  8'h00;      memory[53893] <=  8'h00;      memory[53894] <=  8'h00;      memory[53895] <=  8'h00;      memory[53896] <=  8'h00;      memory[53897] <=  8'h00;      memory[53898] <=  8'h00;      memory[53899] <=  8'h00;      memory[53900] <=  8'h00;      memory[53901] <=  8'h00;      memory[53902] <=  8'h00;      memory[53903] <=  8'h00;      memory[53904] <=  8'h00;      memory[53905] <=  8'h00;      memory[53906] <=  8'h00;      memory[53907] <=  8'h00;      memory[53908] <=  8'h00;      memory[53909] <=  8'h00;      memory[53910] <=  8'h00;      memory[53911] <=  8'h00;      memory[53912] <=  8'h00;      memory[53913] <=  8'h00;      memory[53914] <=  8'h00;      memory[53915] <=  8'h00;      memory[53916] <=  8'h00;      memory[53917] <=  8'h00;      memory[53918] <=  8'h00;      memory[53919] <=  8'h00;      memory[53920] <=  8'h00;      memory[53921] <=  8'h00;      memory[53922] <=  8'h00;      memory[53923] <=  8'h00;      memory[53924] <=  8'h00;      memory[53925] <=  8'h00;      memory[53926] <=  8'h00;      memory[53927] <=  8'h00;      memory[53928] <=  8'h00;      memory[53929] <=  8'h00;      memory[53930] <=  8'h00;      memory[53931] <=  8'h00;      memory[53932] <=  8'h00;      memory[53933] <=  8'h00;      memory[53934] <=  8'h00;      memory[53935] <=  8'h00;      memory[53936] <=  8'h00;      memory[53937] <=  8'h00;      memory[53938] <=  8'h00;      memory[53939] <=  8'h00;      memory[53940] <=  8'h00;      memory[53941] <=  8'h00;      memory[53942] <=  8'h00;      memory[53943] <=  8'h00;      memory[53944] <=  8'h00;      memory[53945] <=  8'h00;      memory[53946] <=  8'h00;      memory[53947] <=  8'h00;      memory[53948] <=  8'h00;      memory[53949] <=  8'h00;      memory[53950] <=  8'h00;      memory[53951] <=  8'h00;      memory[53952] <=  8'h00;      memory[53953] <=  8'h00;      memory[53954] <=  8'h00;      memory[53955] <=  8'h00;      memory[53956] <=  8'h00;      memory[53957] <=  8'h00;      memory[53958] <=  8'h00;      memory[53959] <=  8'h00;      memory[53960] <=  8'h00;      memory[53961] <=  8'h00;      memory[53962] <=  8'h00;      memory[53963] <=  8'h00;      memory[53964] <=  8'h00;      memory[53965] <=  8'h00;      memory[53966] <=  8'h00;      memory[53967] <=  8'h00;      memory[53968] <=  8'h00;      memory[53969] <=  8'h00;      memory[53970] <=  8'h00;      memory[53971] <=  8'h00;      memory[53972] <=  8'h00;      memory[53973] <=  8'h00;      memory[53974] <=  8'h00;      memory[53975] <=  8'h00;      memory[53976] <=  8'h00;      memory[53977] <=  8'h00;      memory[53978] <=  8'h00;      memory[53979] <=  8'h00;      memory[53980] <=  8'h00;      memory[53981] <=  8'h00;      memory[53982] <=  8'h00;      memory[53983] <=  8'h00;      memory[53984] <=  8'h00;      memory[53985] <=  8'h00;      memory[53986] <=  8'h00;      memory[53987] <=  8'h00;      memory[53988] <=  8'h00;      memory[53989] <=  8'h00;      memory[53990] <=  8'h00;      memory[53991] <=  8'h00;      memory[53992] <=  8'h00;      memory[53993] <=  8'h00;      memory[53994] <=  8'h00;      memory[53995] <=  8'h00;      memory[53996] <=  8'h00;      memory[53997] <=  8'h00;      memory[53998] <=  8'h00;      memory[53999] <=  8'h00;      memory[54000] <=  8'h00;      memory[54001] <=  8'h00;      memory[54002] <=  8'h00;      memory[54003] <=  8'h00;      memory[54004] <=  8'h00;      memory[54005] <=  8'h00;      memory[54006] <=  8'h00;      memory[54007] <=  8'h00;      memory[54008] <=  8'h00;      memory[54009] <=  8'h00;      memory[54010] <=  8'h00;      memory[54011] <=  8'h00;      memory[54012] <=  8'h00;      memory[54013] <=  8'h00;      memory[54014] <=  8'h00;      memory[54015] <=  8'h00;      memory[54016] <=  8'h00;      memory[54017] <=  8'h00;      memory[54018] <=  8'h00;      memory[54019] <=  8'h00;      memory[54020] <=  8'h00;      memory[54021] <=  8'h00;      memory[54022] <=  8'h00;      memory[54023] <=  8'h00;      memory[54024] <=  8'h00;      memory[54025] <=  8'h00;      memory[54026] <=  8'h00;      memory[54027] <=  8'h00;      memory[54028] <=  8'h00;      memory[54029] <=  8'h00;      memory[54030] <=  8'h00;      memory[54031] <=  8'h00;      memory[54032] <=  8'h00;      memory[54033] <=  8'h00;      memory[54034] <=  8'h00;      memory[54035] <=  8'h00;      memory[54036] <=  8'h00;      memory[54037] <=  8'h00;      memory[54038] <=  8'h00;      memory[54039] <=  8'h00;      memory[54040] <=  8'h00;      memory[54041] <=  8'h00;      memory[54042] <=  8'h00;      memory[54043] <=  8'h00;      memory[54044] <=  8'h00;      memory[54045] <=  8'h00;      memory[54046] <=  8'h00;      memory[54047] <=  8'h00;      memory[54048] <=  8'h00;      memory[54049] <=  8'h00;      memory[54050] <=  8'h00;      memory[54051] <=  8'h00;      memory[54052] <=  8'h00;      memory[54053] <=  8'h00;      memory[54054] <=  8'h00;      memory[54055] <=  8'h00;      memory[54056] <=  8'h00;      memory[54057] <=  8'h00;      memory[54058] <=  8'h00;      memory[54059] <=  8'h00;      memory[54060] <=  8'h00;      memory[54061] <=  8'h00;      memory[54062] <=  8'h00;      memory[54063] <=  8'h00;      memory[54064] <=  8'h00;      memory[54065] <=  8'h00;      memory[54066] <=  8'h00;      memory[54067] <=  8'h00;      memory[54068] <=  8'h00;      memory[54069] <=  8'h00;      memory[54070] <=  8'h00;      memory[54071] <=  8'h00;      memory[54072] <=  8'h00;      memory[54073] <=  8'h00;      memory[54074] <=  8'h00;      memory[54075] <=  8'h00;      memory[54076] <=  8'h00;      memory[54077] <=  8'h00;      memory[54078] <=  8'h00;      memory[54079] <=  8'h00;      memory[54080] <=  8'h00;      memory[54081] <=  8'h00;      memory[54082] <=  8'h00;      memory[54083] <=  8'h00;      memory[54084] <=  8'h00;      memory[54085] <=  8'h00;      memory[54086] <=  8'h00;      memory[54087] <=  8'h00;      memory[54088] <=  8'h00;      memory[54089] <=  8'h00;      memory[54090] <=  8'h00;      memory[54091] <=  8'h00;      memory[54092] <=  8'h00;      memory[54093] <=  8'h00;      memory[54094] <=  8'h00;      memory[54095] <=  8'h00;      memory[54096] <=  8'h00;      memory[54097] <=  8'h00;      memory[54098] <=  8'h00;      memory[54099] <=  8'h00;      memory[54100] <=  8'h00;      memory[54101] <=  8'h00;      memory[54102] <=  8'h00;      memory[54103] <=  8'h00;      memory[54104] <=  8'h00;      memory[54105] <=  8'h00;      memory[54106] <=  8'h00;      memory[54107] <=  8'h00;      memory[54108] <=  8'h00;      memory[54109] <=  8'h00;      memory[54110] <=  8'h00;      memory[54111] <=  8'h00;      memory[54112] <=  8'h00;      memory[54113] <=  8'h00;      memory[54114] <=  8'h00;      memory[54115] <=  8'h00;      memory[54116] <=  8'h00;      memory[54117] <=  8'h00;      memory[54118] <=  8'h00;      memory[54119] <=  8'h00;      memory[54120] <=  8'h00;      memory[54121] <=  8'h00;      memory[54122] <=  8'h00;      memory[54123] <=  8'h00;      memory[54124] <=  8'h00;      memory[54125] <=  8'h00;      memory[54126] <=  8'h00;      memory[54127] <=  8'h00;      memory[54128] <=  8'h00;      memory[54129] <=  8'h00;      memory[54130] <=  8'h00;      memory[54131] <=  8'h00;      memory[54132] <=  8'h00;      memory[54133] <=  8'h00;      memory[54134] <=  8'h00;      memory[54135] <=  8'h00;      memory[54136] <=  8'h00;      memory[54137] <=  8'h00;      memory[54138] <=  8'h00;      memory[54139] <=  8'h00;      memory[54140] <=  8'h00;      memory[54141] <=  8'h00;      memory[54142] <=  8'h00;      memory[54143] <=  8'h00;      memory[54144] <=  8'h00;      memory[54145] <=  8'h00;      memory[54146] <=  8'h00;      memory[54147] <=  8'h00;      memory[54148] <=  8'h00;      memory[54149] <=  8'h00;      memory[54150] <=  8'h00;      memory[54151] <=  8'h00;      memory[54152] <=  8'h00;      memory[54153] <=  8'h00;      memory[54154] <=  8'h00;      memory[54155] <=  8'h00;      memory[54156] <=  8'h00;      memory[54157] <=  8'h00;      memory[54158] <=  8'h00;      memory[54159] <=  8'h00;      memory[54160] <=  8'h00;      memory[54161] <=  8'h00;      memory[54162] <=  8'h00;      memory[54163] <=  8'h00;      memory[54164] <=  8'h00;      memory[54165] <=  8'h00;      memory[54166] <=  8'h00;      memory[54167] <=  8'h00;      memory[54168] <=  8'h00;      memory[54169] <=  8'h00;      memory[54170] <=  8'h00;      memory[54171] <=  8'h00;      memory[54172] <=  8'h00;      memory[54173] <=  8'h00;      memory[54174] <=  8'h00;      memory[54175] <=  8'h00;      memory[54176] <=  8'h00;      memory[54177] <=  8'h00;      memory[54178] <=  8'h00;      memory[54179] <=  8'h00;      memory[54180] <=  8'h00;      memory[54181] <=  8'h00;      memory[54182] <=  8'h00;      memory[54183] <=  8'h00;      memory[54184] <=  8'h00;      memory[54185] <=  8'h00;      memory[54186] <=  8'h00;      memory[54187] <=  8'h00;      memory[54188] <=  8'h00;      memory[54189] <=  8'h00;      memory[54190] <=  8'h00;      memory[54191] <=  8'h00;      memory[54192] <=  8'h00;      memory[54193] <=  8'h00;      memory[54194] <=  8'h00;      memory[54195] <=  8'h00;      memory[54196] <=  8'h00;      memory[54197] <=  8'h00;      memory[54198] <=  8'h00;      memory[54199] <=  8'h00;      memory[54200] <=  8'h00;      memory[54201] <=  8'h00;      memory[54202] <=  8'h00;      memory[54203] <=  8'h00;      memory[54204] <=  8'h00;      memory[54205] <=  8'h00;      memory[54206] <=  8'h00;      memory[54207] <=  8'h00;      memory[54208] <=  8'h00;      memory[54209] <=  8'h00;      memory[54210] <=  8'h00;      memory[54211] <=  8'h00;      memory[54212] <=  8'h00;      memory[54213] <=  8'h00;      memory[54214] <=  8'h00;      memory[54215] <=  8'h00;      memory[54216] <=  8'h00;      memory[54217] <=  8'h00;      memory[54218] <=  8'h00;      memory[54219] <=  8'h00;      memory[54220] <=  8'h00;      memory[54221] <=  8'h00;      memory[54222] <=  8'h00;      memory[54223] <=  8'h00;      memory[54224] <=  8'h00;      memory[54225] <=  8'h00;      memory[54226] <=  8'h00;      memory[54227] <=  8'h00;      memory[54228] <=  8'h00;      memory[54229] <=  8'h00;      memory[54230] <=  8'h00;      memory[54231] <=  8'h00;      memory[54232] <=  8'h00;      memory[54233] <=  8'h00;      memory[54234] <=  8'h00;      memory[54235] <=  8'h00;      memory[54236] <=  8'h00;      memory[54237] <=  8'h00;      memory[54238] <=  8'h00;      memory[54239] <=  8'h00;      memory[54240] <=  8'h00;      memory[54241] <=  8'h00;      memory[54242] <=  8'h00;      memory[54243] <=  8'h00;      memory[54244] <=  8'h00;      memory[54245] <=  8'h00;      memory[54246] <=  8'h00;      memory[54247] <=  8'h00;      memory[54248] <=  8'h00;      memory[54249] <=  8'h00;      memory[54250] <=  8'h00;      memory[54251] <=  8'h00;      memory[54252] <=  8'h00;      memory[54253] <=  8'h00;      memory[54254] <=  8'h00;      memory[54255] <=  8'h00;      memory[54256] <=  8'h00;      memory[54257] <=  8'h00;      memory[54258] <=  8'h00;      memory[54259] <=  8'h00;      memory[54260] <=  8'h00;      memory[54261] <=  8'h00;      memory[54262] <=  8'h00;      memory[54263] <=  8'h00;      memory[54264] <=  8'h00;      memory[54265] <=  8'h00;      memory[54266] <=  8'h00;      memory[54267] <=  8'h00;      memory[54268] <=  8'h00;      memory[54269] <=  8'h00;      memory[54270] <=  8'h00;      memory[54271] <=  8'h00;      memory[54272] <=  8'h00;      memory[54273] <=  8'h00;      memory[54274] <=  8'h00;      memory[54275] <=  8'h00;      memory[54276] <=  8'h00;      memory[54277] <=  8'h00;      memory[54278] <=  8'h00;      memory[54279] <=  8'h00;      memory[54280] <=  8'h00;      memory[54281] <=  8'h00;      memory[54282] <=  8'h00;      memory[54283] <=  8'h00;      memory[54284] <=  8'h00;      memory[54285] <=  8'h00;      memory[54286] <=  8'h00;      memory[54287] <=  8'h00;      memory[54288] <=  8'h00;      memory[54289] <=  8'h00;      memory[54290] <=  8'h00;      memory[54291] <=  8'h00;      memory[54292] <=  8'h00;      memory[54293] <=  8'h00;      memory[54294] <=  8'h00;      memory[54295] <=  8'h00;      memory[54296] <=  8'h00;      memory[54297] <=  8'h00;      memory[54298] <=  8'h00;      memory[54299] <=  8'h00;      memory[54300] <=  8'h00;      memory[54301] <=  8'h00;      memory[54302] <=  8'h00;      memory[54303] <=  8'h00;      memory[54304] <=  8'h00;      memory[54305] <=  8'h00;      memory[54306] <=  8'h00;      memory[54307] <=  8'h00;      memory[54308] <=  8'h00;      memory[54309] <=  8'h00;      memory[54310] <=  8'h00;      memory[54311] <=  8'h00;      memory[54312] <=  8'h00;      memory[54313] <=  8'h00;      memory[54314] <=  8'h00;      memory[54315] <=  8'h00;      memory[54316] <=  8'h00;      memory[54317] <=  8'h00;      memory[54318] <=  8'h00;      memory[54319] <=  8'h00;      memory[54320] <=  8'h00;      memory[54321] <=  8'h00;      memory[54322] <=  8'h00;      memory[54323] <=  8'h00;      memory[54324] <=  8'h00;      memory[54325] <=  8'h00;      memory[54326] <=  8'h00;      memory[54327] <=  8'h00;      memory[54328] <=  8'h00;      memory[54329] <=  8'h00;      memory[54330] <=  8'h00;      memory[54331] <=  8'h00;      memory[54332] <=  8'h00;      memory[54333] <=  8'h00;      memory[54334] <=  8'h00;      memory[54335] <=  8'h00;      memory[54336] <=  8'h00;      memory[54337] <=  8'h00;      memory[54338] <=  8'h00;      memory[54339] <=  8'h00;      memory[54340] <=  8'h00;      memory[54341] <=  8'h00;      memory[54342] <=  8'h00;      memory[54343] <=  8'h00;      memory[54344] <=  8'h00;      memory[54345] <=  8'h00;      memory[54346] <=  8'h00;      memory[54347] <=  8'h00;      memory[54348] <=  8'h00;      memory[54349] <=  8'h00;      memory[54350] <=  8'h00;      memory[54351] <=  8'h00;      memory[54352] <=  8'h00;      memory[54353] <=  8'h00;      memory[54354] <=  8'h00;      memory[54355] <=  8'h00;      memory[54356] <=  8'h00;      memory[54357] <=  8'h00;      memory[54358] <=  8'h00;      memory[54359] <=  8'h00;      memory[54360] <=  8'h00;      memory[54361] <=  8'h00;      memory[54362] <=  8'h00;      memory[54363] <=  8'h00;      memory[54364] <=  8'h00;      memory[54365] <=  8'h00;      memory[54366] <=  8'h00;      memory[54367] <=  8'h00;      memory[54368] <=  8'h00;      memory[54369] <=  8'h00;      memory[54370] <=  8'h00;      memory[54371] <=  8'h00;      memory[54372] <=  8'h00;      memory[54373] <=  8'h00;      memory[54374] <=  8'h00;      memory[54375] <=  8'h00;      memory[54376] <=  8'h00;      memory[54377] <=  8'h00;      memory[54378] <=  8'h00;      memory[54379] <=  8'h00;      memory[54380] <=  8'h00;      memory[54381] <=  8'h00;      memory[54382] <=  8'h00;      memory[54383] <=  8'h00;      memory[54384] <=  8'h00;      memory[54385] <=  8'h00;      memory[54386] <=  8'h00;      memory[54387] <=  8'h00;      memory[54388] <=  8'h00;      memory[54389] <=  8'h00;      memory[54390] <=  8'h00;      memory[54391] <=  8'h00;      memory[54392] <=  8'h00;      memory[54393] <=  8'h00;      memory[54394] <=  8'h00;      memory[54395] <=  8'h00;      memory[54396] <=  8'h00;      memory[54397] <=  8'h00;      memory[54398] <=  8'h00;      memory[54399] <=  8'h00;      memory[54400] <=  8'h00;      memory[54401] <=  8'h00;      memory[54402] <=  8'h00;      memory[54403] <=  8'h00;      memory[54404] <=  8'h00;      memory[54405] <=  8'h00;      memory[54406] <=  8'h00;      memory[54407] <=  8'h00;      memory[54408] <=  8'h00;      memory[54409] <=  8'h00;      memory[54410] <=  8'h00;      memory[54411] <=  8'h00;      memory[54412] <=  8'h00;      memory[54413] <=  8'h00;      memory[54414] <=  8'h00;      memory[54415] <=  8'h00;      memory[54416] <=  8'h00;      memory[54417] <=  8'h00;      memory[54418] <=  8'h00;      memory[54419] <=  8'h00;      memory[54420] <=  8'h00;      memory[54421] <=  8'h00;      memory[54422] <=  8'h00;      memory[54423] <=  8'h00;      memory[54424] <=  8'h00;      memory[54425] <=  8'h00;      memory[54426] <=  8'h00;      memory[54427] <=  8'h00;      memory[54428] <=  8'h00;      memory[54429] <=  8'h00;      memory[54430] <=  8'h00;      memory[54431] <=  8'h00;      memory[54432] <=  8'h00;      memory[54433] <=  8'h00;      memory[54434] <=  8'h00;      memory[54435] <=  8'h00;      memory[54436] <=  8'h00;      memory[54437] <=  8'h00;      memory[54438] <=  8'h00;      memory[54439] <=  8'h00;      memory[54440] <=  8'h00;      memory[54441] <=  8'h00;      memory[54442] <=  8'h00;      memory[54443] <=  8'h00;      memory[54444] <=  8'h00;      memory[54445] <=  8'h00;      memory[54446] <=  8'h00;      memory[54447] <=  8'h00;      memory[54448] <=  8'h00;      memory[54449] <=  8'h00;      memory[54450] <=  8'h00;      memory[54451] <=  8'h00;      memory[54452] <=  8'h00;      memory[54453] <=  8'h00;      memory[54454] <=  8'h00;      memory[54455] <=  8'h00;      memory[54456] <=  8'h00;      memory[54457] <=  8'h00;      memory[54458] <=  8'h00;      memory[54459] <=  8'h00;      memory[54460] <=  8'h00;      memory[54461] <=  8'h00;      memory[54462] <=  8'h00;      memory[54463] <=  8'h00;      memory[54464] <=  8'h00;      memory[54465] <=  8'h00;      memory[54466] <=  8'h00;      memory[54467] <=  8'h00;      memory[54468] <=  8'h00;      memory[54469] <=  8'h00;      memory[54470] <=  8'h00;      memory[54471] <=  8'h00;      memory[54472] <=  8'h00;      memory[54473] <=  8'h00;      memory[54474] <=  8'h00;      memory[54475] <=  8'h00;      memory[54476] <=  8'h00;      memory[54477] <=  8'h00;      memory[54478] <=  8'h00;      memory[54479] <=  8'h00;      memory[54480] <=  8'h00;      memory[54481] <=  8'h00;      memory[54482] <=  8'h00;      memory[54483] <=  8'h00;      memory[54484] <=  8'h00;      memory[54485] <=  8'h00;      memory[54486] <=  8'h00;      memory[54487] <=  8'h00;      memory[54488] <=  8'h00;      memory[54489] <=  8'h00;      memory[54490] <=  8'h00;      memory[54491] <=  8'h00;      memory[54492] <=  8'h00;      memory[54493] <=  8'h00;      memory[54494] <=  8'h00;      memory[54495] <=  8'h00;      memory[54496] <=  8'h00;      memory[54497] <=  8'h00;      memory[54498] <=  8'h00;      memory[54499] <=  8'h00;      memory[54500] <=  8'h00;      memory[54501] <=  8'h00;      memory[54502] <=  8'h00;      memory[54503] <=  8'h00;      memory[54504] <=  8'h00;      memory[54505] <=  8'h00;      memory[54506] <=  8'h00;      memory[54507] <=  8'h00;      memory[54508] <=  8'h00;      memory[54509] <=  8'h00;      memory[54510] <=  8'h00;      memory[54511] <=  8'h00;      memory[54512] <=  8'h00;      memory[54513] <=  8'h00;      memory[54514] <=  8'h00;      memory[54515] <=  8'h00;      memory[54516] <=  8'h00;      memory[54517] <=  8'h00;      memory[54518] <=  8'h00;      memory[54519] <=  8'h00;      memory[54520] <=  8'h00;      memory[54521] <=  8'h00;      memory[54522] <=  8'h00;      memory[54523] <=  8'h00;      memory[54524] <=  8'h00;      memory[54525] <=  8'h00;      memory[54526] <=  8'h00;      memory[54527] <=  8'h00;      memory[54528] <=  8'h00;      memory[54529] <=  8'h00;      memory[54530] <=  8'h00;      memory[54531] <=  8'h00;      memory[54532] <=  8'h00;      memory[54533] <=  8'h00;      memory[54534] <=  8'h00;      memory[54535] <=  8'h00;      memory[54536] <=  8'h00;      memory[54537] <=  8'h00;      memory[54538] <=  8'h00;      memory[54539] <=  8'h00;      memory[54540] <=  8'h00;      memory[54541] <=  8'h00;      memory[54542] <=  8'h00;      memory[54543] <=  8'h00;      memory[54544] <=  8'h00;      memory[54545] <=  8'h00;      memory[54546] <=  8'h00;      memory[54547] <=  8'h00;      memory[54548] <=  8'h00;      memory[54549] <=  8'h00;      memory[54550] <=  8'h00;      memory[54551] <=  8'h00;      memory[54552] <=  8'h00;      memory[54553] <=  8'h00;      memory[54554] <=  8'h00;      memory[54555] <=  8'h00;      memory[54556] <=  8'h00;      memory[54557] <=  8'h00;      memory[54558] <=  8'h00;      memory[54559] <=  8'h00;      memory[54560] <=  8'h00;      memory[54561] <=  8'h00;      memory[54562] <=  8'h00;      memory[54563] <=  8'h00;      memory[54564] <=  8'h00;      memory[54565] <=  8'h00;      memory[54566] <=  8'h00;      memory[54567] <=  8'h00;      memory[54568] <=  8'h00;      memory[54569] <=  8'h00;      memory[54570] <=  8'h00;      memory[54571] <=  8'h00;      memory[54572] <=  8'h00;      memory[54573] <=  8'h00;      memory[54574] <=  8'h00;      memory[54575] <=  8'h00;      memory[54576] <=  8'h00;      memory[54577] <=  8'h00;      memory[54578] <=  8'h00;      memory[54579] <=  8'h00;      memory[54580] <=  8'h00;      memory[54581] <=  8'h00;      memory[54582] <=  8'h00;      memory[54583] <=  8'h00;      memory[54584] <=  8'h00;      memory[54585] <=  8'h00;      memory[54586] <=  8'h00;      memory[54587] <=  8'h00;      memory[54588] <=  8'h00;      memory[54589] <=  8'h00;      memory[54590] <=  8'h00;      memory[54591] <=  8'h00;      memory[54592] <=  8'h00;      memory[54593] <=  8'h00;      memory[54594] <=  8'h00;      memory[54595] <=  8'h00;      memory[54596] <=  8'h00;      memory[54597] <=  8'h00;      memory[54598] <=  8'h00;      memory[54599] <=  8'h00;      memory[54600] <=  8'h00;      memory[54601] <=  8'h00;      memory[54602] <=  8'h00;      memory[54603] <=  8'h00;      memory[54604] <=  8'h00;      memory[54605] <=  8'h00;      memory[54606] <=  8'h00;      memory[54607] <=  8'h00;      memory[54608] <=  8'h00;      memory[54609] <=  8'h00;      memory[54610] <=  8'h00;      memory[54611] <=  8'h00;      memory[54612] <=  8'h00;      memory[54613] <=  8'h00;      memory[54614] <=  8'h00;      memory[54615] <=  8'h00;      memory[54616] <=  8'h00;      memory[54617] <=  8'h00;      memory[54618] <=  8'h00;      memory[54619] <=  8'h00;      memory[54620] <=  8'h00;      memory[54621] <=  8'h00;      memory[54622] <=  8'h00;      memory[54623] <=  8'h00;      memory[54624] <=  8'h00;      memory[54625] <=  8'h00;      memory[54626] <=  8'h00;      memory[54627] <=  8'h00;      memory[54628] <=  8'h00;      memory[54629] <=  8'h00;      memory[54630] <=  8'h00;      memory[54631] <=  8'h00;      memory[54632] <=  8'h00;      memory[54633] <=  8'h00;      memory[54634] <=  8'h00;      memory[54635] <=  8'h00;      memory[54636] <=  8'h00;      memory[54637] <=  8'h00;      memory[54638] <=  8'h00;      memory[54639] <=  8'h00;      memory[54640] <=  8'h00;      memory[54641] <=  8'h00;      memory[54642] <=  8'h00;      memory[54643] <=  8'h00;      memory[54644] <=  8'h00;      memory[54645] <=  8'h00;      memory[54646] <=  8'h00;      memory[54647] <=  8'h00;      memory[54648] <=  8'h00;      memory[54649] <=  8'h00;      memory[54650] <=  8'h00;      memory[54651] <=  8'h00;      memory[54652] <=  8'h00;      memory[54653] <=  8'h00;      memory[54654] <=  8'h00;      memory[54655] <=  8'h00;      memory[54656] <=  8'h00;      memory[54657] <=  8'h00;      memory[54658] <=  8'h00;      memory[54659] <=  8'h00;      memory[54660] <=  8'h00;      memory[54661] <=  8'h00;      memory[54662] <=  8'h00;      memory[54663] <=  8'h00;      memory[54664] <=  8'h00;      memory[54665] <=  8'h00;      memory[54666] <=  8'h00;      memory[54667] <=  8'h00;      memory[54668] <=  8'h00;      memory[54669] <=  8'h00;      memory[54670] <=  8'h00;      memory[54671] <=  8'h00;      memory[54672] <=  8'h00;      memory[54673] <=  8'h00;      memory[54674] <=  8'h00;      memory[54675] <=  8'h00;      memory[54676] <=  8'h00;      memory[54677] <=  8'h00;      memory[54678] <=  8'h00;      memory[54679] <=  8'h00;      memory[54680] <=  8'h00;      memory[54681] <=  8'h00;      memory[54682] <=  8'h00;      memory[54683] <=  8'h00;      memory[54684] <=  8'h00;      memory[54685] <=  8'h00;      memory[54686] <=  8'h00;      memory[54687] <=  8'h00;      memory[54688] <=  8'h00;      memory[54689] <=  8'h00;      memory[54690] <=  8'h00;      memory[54691] <=  8'h00;      memory[54692] <=  8'h00;      memory[54693] <=  8'h00;      memory[54694] <=  8'h00;      memory[54695] <=  8'h00;      memory[54696] <=  8'h00;      memory[54697] <=  8'h00;      memory[54698] <=  8'h00;      memory[54699] <=  8'h00;      memory[54700] <=  8'h00;      memory[54701] <=  8'h00;      memory[54702] <=  8'h00;      memory[54703] <=  8'h00;      memory[54704] <=  8'h00;      memory[54705] <=  8'h00;      memory[54706] <=  8'h00;      memory[54707] <=  8'h00;      memory[54708] <=  8'h00;      memory[54709] <=  8'h00;      memory[54710] <=  8'h00;      memory[54711] <=  8'h00;      memory[54712] <=  8'h00;      memory[54713] <=  8'h00;      memory[54714] <=  8'h00;      memory[54715] <=  8'h00;      memory[54716] <=  8'h00;      memory[54717] <=  8'h00;      memory[54718] <=  8'h00;      memory[54719] <=  8'h00;      memory[54720] <=  8'h00;      memory[54721] <=  8'h00;      memory[54722] <=  8'h00;      memory[54723] <=  8'h00;      memory[54724] <=  8'h00;      memory[54725] <=  8'h00;      memory[54726] <=  8'h00;      memory[54727] <=  8'h00;      memory[54728] <=  8'h00;      memory[54729] <=  8'h00;      memory[54730] <=  8'h00;      memory[54731] <=  8'h00;      memory[54732] <=  8'h00;      memory[54733] <=  8'h00;      memory[54734] <=  8'h00;      memory[54735] <=  8'h00;      memory[54736] <=  8'h00;      memory[54737] <=  8'h00;      memory[54738] <=  8'h00;      memory[54739] <=  8'h00;      memory[54740] <=  8'h00;      memory[54741] <=  8'h00;      memory[54742] <=  8'h00;      memory[54743] <=  8'h00;      memory[54744] <=  8'h00;      memory[54745] <=  8'h00;      memory[54746] <=  8'h00;      memory[54747] <=  8'h00;      memory[54748] <=  8'h00;      memory[54749] <=  8'h00;      memory[54750] <=  8'h00;      memory[54751] <=  8'h00;      memory[54752] <=  8'h00;      memory[54753] <=  8'h00;      memory[54754] <=  8'h00;      memory[54755] <=  8'h00;      memory[54756] <=  8'h00;      memory[54757] <=  8'h00;      memory[54758] <=  8'h00;      memory[54759] <=  8'h00;      memory[54760] <=  8'h00;      memory[54761] <=  8'h00;      memory[54762] <=  8'h00;      memory[54763] <=  8'h00;      memory[54764] <=  8'h00;      memory[54765] <=  8'h00;      memory[54766] <=  8'h00;      memory[54767] <=  8'h00;      memory[54768] <=  8'h00;      memory[54769] <=  8'h00;      memory[54770] <=  8'h00;      memory[54771] <=  8'h00;      memory[54772] <=  8'h00;      memory[54773] <=  8'h00;      memory[54774] <=  8'h00;      memory[54775] <=  8'h00;      memory[54776] <=  8'h00;      memory[54777] <=  8'h00;      memory[54778] <=  8'h00;      memory[54779] <=  8'h00;      memory[54780] <=  8'h00;      memory[54781] <=  8'h00;      memory[54782] <=  8'h00;      memory[54783] <=  8'h00;      memory[54784] <=  8'h00;      memory[54785] <=  8'h00;      memory[54786] <=  8'h00;      memory[54787] <=  8'h00;      memory[54788] <=  8'h00;      memory[54789] <=  8'h00;      memory[54790] <=  8'h00;      memory[54791] <=  8'h00;      memory[54792] <=  8'h00;      memory[54793] <=  8'h00;      memory[54794] <=  8'h00;      memory[54795] <=  8'h00;      memory[54796] <=  8'h00;      memory[54797] <=  8'h00;      memory[54798] <=  8'h00;      memory[54799] <=  8'h00;      memory[54800] <=  8'h00;      memory[54801] <=  8'h00;      memory[54802] <=  8'h00;      memory[54803] <=  8'h00;      memory[54804] <=  8'h00;      memory[54805] <=  8'h00;      memory[54806] <=  8'h00;      memory[54807] <=  8'h00;      memory[54808] <=  8'h00;      memory[54809] <=  8'h00;      memory[54810] <=  8'h00;      memory[54811] <=  8'h00;      memory[54812] <=  8'h00;      memory[54813] <=  8'h00;      memory[54814] <=  8'h00;      memory[54815] <=  8'h00;      memory[54816] <=  8'h00;      memory[54817] <=  8'h00;      memory[54818] <=  8'h00;      memory[54819] <=  8'h00;      memory[54820] <=  8'h00;      memory[54821] <=  8'h00;      memory[54822] <=  8'h00;      memory[54823] <=  8'h00;      memory[54824] <=  8'h00;      memory[54825] <=  8'h00;      memory[54826] <=  8'h00;      memory[54827] <=  8'h00;      memory[54828] <=  8'h00;      memory[54829] <=  8'h00;      memory[54830] <=  8'h00;      memory[54831] <=  8'h00;      memory[54832] <=  8'h00;      memory[54833] <=  8'h00;      memory[54834] <=  8'h00;      memory[54835] <=  8'h00;      memory[54836] <=  8'h00;      memory[54837] <=  8'h00;      memory[54838] <=  8'h00;      memory[54839] <=  8'h00;      memory[54840] <=  8'h00;      memory[54841] <=  8'h00;      memory[54842] <=  8'h00;      memory[54843] <=  8'h00;      memory[54844] <=  8'h00;      memory[54845] <=  8'h00;      memory[54846] <=  8'h00;      memory[54847] <=  8'h00;      memory[54848] <=  8'h00;      memory[54849] <=  8'h00;      memory[54850] <=  8'h00;      memory[54851] <=  8'h00;      memory[54852] <=  8'h00;      memory[54853] <=  8'h00;      memory[54854] <=  8'h00;      memory[54855] <=  8'h00;      memory[54856] <=  8'h00;      memory[54857] <=  8'h00;      memory[54858] <=  8'h00;      memory[54859] <=  8'h00;      memory[54860] <=  8'h00;      memory[54861] <=  8'h00;      memory[54862] <=  8'h00;      memory[54863] <=  8'h00;      memory[54864] <=  8'h00;      memory[54865] <=  8'h00;      memory[54866] <=  8'h00;      memory[54867] <=  8'h00;      memory[54868] <=  8'h00;      memory[54869] <=  8'h00;      memory[54870] <=  8'h00;      memory[54871] <=  8'h00;      memory[54872] <=  8'h00;      memory[54873] <=  8'h00;      memory[54874] <=  8'h00;      memory[54875] <=  8'h00;      memory[54876] <=  8'h00;      memory[54877] <=  8'h00;      memory[54878] <=  8'h00;      memory[54879] <=  8'h00;      memory[54880] <=  8'h00;      memory[54881] <=  8'h00;      memory[54882] <=  8'h00;      memory[54883] <=  8'h00;      memory[54884] <=  8'h00;      memory[54885] <=  8'h00;      memory[54886] <=  8'h00;      memory[54887] <=  8'h00;      memory[54888] <=  8'h00;      memory[54889] <=  8'h00;      memory[54890] <=  8'h00;      memory[54891] <=  8'h00;      memory[54892] <=  8'h00;      memory[54893] <=  8'h00;      memory[54894] <=  8'h00;      memory[54895] <=  8'h00;      memory[54896] <=  8'h00;      memory[54897] <=  8'h00;      memory[54898] <=  8'h00;      memory[54899] <=  8'h00;      memory[54900] <=  8'h00;      memory[54901] <=  8'h00;      memory[54902] <=  8'h00;      memory[54903] <=  8'h00;      memory[54904] <=  8'h00;      memory[54905] <=  8'h00;      memory[54906] <=  8'h00;      memory[54907] <=  8'h00;      memory[54908] <=  8'h00;      memory[54909] <=  8'h00;      memory[54910] <=  8'h00;      memory[54911] <=  8'h00;      memory[54912] <=  8'h00;      memory[54913] <=  8'h00;      memory[54914] <=  8'h00;      memory[54915] <=  8'h00;      memory[54916] <=  8'h00;      memory[54917] <=  8'h00;      memory[54918] <=  8'h00;      memory[54919] <=  8'h00;      memory[54920] <=  8'h00;      memory[54921] <=  8'h00;      memory[54922] <=  8'h00;      memory[54923] <=  8'h00;      memory[54924] <=  8'h00;      memory[54925] <=  8'h00;      memory[54926] <=  8'h00;      memory[54927] <=  8'h00;      memory[54928] <=  8'h00;      memory[54929] <=  8'h00;      memory[54930] <=  8'h00;      memory[54931] <=  8'h00;      memory[54932] <=  8'h00;      memory[54933] <=  8'h00;      memory[54934] <=  8'h00;      memory[54935] <=  8'h00;      memory[54936] <=  8'h00;      memory[54937] <=  8'h00;      memory[54938] <=  8'h00;      memory[54939] <=  8'h00;      memory[54940] <=  8'h00;      memory[54941] <=  8'h00;      memory[54942] <=  8'h00;      memory[54943] <=  8'h00;      memory[54944] <=  8'h00;      memory[54945] <=  8'h00;      memory[54946] <=  8'h00;      memory[54947] <=  8'h00;      memory[54948] <=  8'h00;      memory[54949] <=  8'h00;      memory[54950] <=  8'h00;      memory[54951] <=  8'h00;      memory[54952] <=  8'h00;      memory[54953] <=  8'h00;      memory[54954] <=  8'h00;      memory[54955] <=  8'h00;      memory[54956] <=  8'h00;      memory[54957] <=  8'h00;      memory[54958] <=  8'h00;      memory[54959] <=  8'h00;      memory[54960] <=  8'h00;      memory[54961] <=  8'h00;      memory[54962] <=  8'h00;      memory[54963] <=  8'h00;      memory[54964] <=  8'h00;      memory[54965] <=  8'h00;      memory[54966] <=  8'h00;      memory[54967] <=  8'h00;      memory[54968] <=  8'h00;      memory[54969] <=  8'h00;      memory[54970] <=  8'h00;      memory[54971] <=  8'h00;      memory[54972] <=  8'h00;      memory[54973] <=  8'h00;      memory[54974] <=  8'h00;      memory[54975] <=  8'h00;      memory[54976] <=  8'h00;      memory[54977] <=  8'h00;      memory[54978] <=  8'h00;      memory[54979] <=  8'h00;      memory[54980] <=  8'h00;      memory[54981] <=  8'h00;      memory[54982] <=  8'h00;      memory[54983] <=  8'h00;      memory[54984] <=  8'h00;      memory[54985] <=  8'h00;      memory[54986] <=  8'h00;      memory[54987] <=  8'h00;      memory[54988] <=  8'h00;      memory[54989] <=  8'h00;      memory[54990] <=  8'h00;      memory[54991] <=  8'h00;      memory[54992] <=  8'h00;      memory[54993] <=  8'h00;      memory[54994] <=  8'h00;      memory[54995] <=  8'h00;      memory[54996] <=  8'h00;      memory[54997] <=  8'h00;      memory[54998] <=  8'h00;      memory[54999] <=  8'h00;      memory[55000] <=  8'h00;      memory[55001] <=  8'h00;      memory[55002] <=  8'h00;      memory[55003] <=  8'h00;      memory[55004] <=  8'h00;      memory[55005] <=  8'h00;      memory[55006] <=  8'h00;      memory[55007] <=  8'h00;      memory[55008] <=  8'h00;      memory[55009] <=  8'h00;      memory[55010] <=  8'h00;      memory[55011] <=  8'h00;      memory[55012] <=  8'h00;      memory[55013] <=  8'h00;      memory[55014] <=  8'h00;      memory[55015] <=  8'h00;      memory[55016] <=  8'h00;      memory[55017] <=  8'h00;      memory[55018] <=  8'h00;      memory[55019] <=  8'h00;      memory[55020] <=  8'h00;      memory[55021] <=  8'h00;      memory[55022] <=  8'h00;      memory[55023] <=  8'h00;      memory[55024] <=  8'h00;      memory[55025] <=  8'h00;      memory[55026] <=  8'h00;      memory[55027] <=  8'h00;      memory[55028] <=  8'h00;      memory[55029] <=  8'h00;      memory[55030] <=  8'h00;      memory[55031] <=  8'h00;      memory[55032] <=  8'h00;      memory[55033] <=  8'h00;      memory[55034] <=  8'h00;      memory[55035] <=  8'h00;      memory[55036] <=  8'h00;      memory[55037] <=  8'h00;      memory[55038] <=  8'h00;      memory[55039] <=  8'h00;      memory[55040] <=  8'h00;      memory[55041] <=  8'h00;      memory[55042] <=  8'h00;      memory[55043] <=  8'h00;      memory[55044] <=  8'h00;      memory[55045] <=  8'h00;      memory[55046] <=  8'h00;      memory[55047] <=  8'h00;      memory[55048] <=  8'h00;      memory[55049] <=  8'h00;      memory[55050] <=  8'h00;      memory[55051] <=  8'h00;      memory[55052] <=  8'h00;      memory[55053] <=  8'h00;      memory[55054] <=  8'h00;      memory[55055] <=  8'h00;      memory[55056] <=  8'h00;      memory[55057] <=  8'h00;      memory[55058] <=  8'h00;      memory[55059] <=  8'h00;      memory[55060] <=  8'h00;      memory[55061] <=  8'h00;      memory[55062] <=  8'h00;      memory[55063] <=  8'h00;      memory[55064] <=  8'h00;      memory[55065] <=  8'h00;      memory[55066] <=  8'h00;      memory[55067] <=  8'h00;      memory[55068] <=  8'h00;      memory[55069] <=  8'h00;      memory[55070] <=  8'h00;      memory[55071] <=  8'h00;      memory[55072] <=  8'h00;      memory[55073] <=  8'h00;      memory[55074] <=  8'h00;      memory[55075] <=  8'h00;      memory[55076] <=  8'h00;      memory[55077] <=  8'h00;      memory[55078] <=  8'h00;      memory[55079] <=  8'h00;      memory[55080] <=  8'h00;      memory[55081] <=  8'h00;      memory[55082] <=  8'h00;      memory[55083] <=  8'h00;      memory[55084] <=  8'h00;      memory[55085] <=  8'h00;      memory[55086] <=  8'h00;      memory[55087] <=  8'h00;      memory[55088] <=  8'h00;      memory[55089] <=  8'h00;      memory[55090] <=  8'h00;      memory[55091] <=  8'h00;      memory[55092] <=  8'h00;      memory[55093] <=  8'h00;      memory[55094] <=  8'h00;      memory[55095] <=  8'h00;      memory[55096] <=  8'h00;      memory[55097] <=  8'h00;      memory[55098] <=  8'h00;      memory[55099] <=  8'h00;      memory[55100] <=  8'h00;      memory[55101] <=  8'h00;      memory[55102] <=  8'h00;      memory[55103] <=  8'h00;      memory[55104] <=  8'h00;      memory[55105] <=  8'h00;      memory[55106] <=  8'h00;      memory[55107] <=  8'h00;      memory[55108] <=  8'h00;      memory[55109] <=  8'h00;      memory[55110] <=  8'h00;      memory[55111] <=  8'h00;      memory[55112] <=  8'h00;      memory[55113] <=  8'h00;      memory[55114] <=  8'h00;      memory[55115] <=  8'h00;      memory[55116] <=  8'h00;      memory[55117] <=  8'h00;      memory[55118] <=  8'h00;      memory[55119] <=  8'h00;      memory[55120] <=  8'h00;      memory[55121] <=  8'h00;      memory[55122] <=  8'h00;      memory[55123] <=  8'h00;      memory[55124] <=  8'h00;      memory[55125] <=  8'h00;      memory[55126] <=  8'h00;      memory[55127] <=  8'h00;      memory[55128] <=  8'h00;      memory[55129] <=  8'h00;      memory[55130] <=  8'h00;      memory[55131] <=  8'h00;      memory[55132] <=  8'h00;      memory[55133] <=  8'h00;      memory[55134] <=  8'h00;      memory[55135] <=  8'h00;      memory[55136] <=  8'h00;      memory[55137] <=  8'h00;      memory[55138] <=  8'h00;      memory[55139] <=  8'h00;      memory[55140] <=  8'h00;      memory[55141] <=  8'h00;      memory[55142] <=  8'h00;      memory[55143] <=  8'h00;      memory[55144] <=  8'h00;      memory[55145] <=  8'h00;      memory[55146] <=  8'h00;      memory[55147] <=  8'h00;      memory[55148] <=  8'h00;      memory[55149] <=  8'h00;      memory[55150] <=  8'h00;      memory[55151] <=  8'h00;      memory[55152] <=  8'h00;      memory[55153] <=  8'h00;      memory[55154] <=  8'h00;      memory[55155] <=  8'h00;      memory[55156] <=  8'h00;      memory[55157] <=  8'h00;      memory[55158] <=  8'h00;      memory[55159] <=  8'h00;      memory[55160] <=  8'h00;      memory[55161] <=  8'h00;      memory[55162] <=  8'h00;      memory[55163] <=  8'h00;      memory[55164] <=  8'h00;      memory[55165] <=  8'h00;      memory[55166] <=  8'h00;      memory[55167] <=  8'h00;      memory[55168] <=  8'h00;      memory[55169] <=  8'h00;      memory[55170] <=  8'h00;      memory[55171] <=  8'h00;      memory[55172] <=  8'h00;      memory[55173] <=  8'h00;      memory[55174] <=  8'h00;      memory[55175] <=  8'h00;      memory[55176] <=  8'h00;      memory[55177] <=  8'h00;      memory[55178] <=  8'h00;      memory[55179] <=  8'h00;      memory[55180] <=  8'h00;      memory[55181] <=  8'h00;      memory[55182] <=  8'h00;      memory[55183] <=  8'h00;      memory[55184] <=  8'h00;      memory[55185] <=  8'h00;      memory[55186] <=  8'h00;      memory[55187] <=  8'h00;      memory[55188] <=  8'h00;      memory[55189] <=  8'h00;      memory[55190] <=  8'h00;      memory[55191] <=  8'h00;      memory[55192] <=  8'h00;      memory[55193] <=  8'h00;      memory[55194] <=  8'h00;      memory[55195] <=  8'h00;      memory[55196] <=  8'h00;      memory[55197] <=  8'h00;      memory[55198] <=  8'h00;      memory[55199] <=  8'h00;      memory[55200] <=  8'h00;      memory[55201] <=  8'h00;      memory[55202] <=  8'h00;      memory[55203] <=  8'h00;      memory[55204] <=  8'h00;      memory[55205] <=  8'h00;      memory[55206] <=  8'h00;      memory[55207] <=  8'h00;      memory[55208] <=  8'h00;      memory[55209] <=  8'h00;      memory[55210] <=  8'h00;      memory[55211] <=  8'h00;      memory[55212] <=  8'h00;      memory[55213] <=  8'h00;      memory[55214] <=  8'h00;      memory[55215] <=  8'h00;      memory[55216] <=  8'h00;      memory[55217] <=  8'h00;      memory[55218] <=  8'h00;      memory[55219] <=  8'h00;      memory[55220] <=  8'h00;      memory[55221] <=  8'h00;      memory[55222] <=  8'h00;      memory[55223] <=  8'h00;      memory[55224] <=  8'h00;      memory[55225] <=  8'h00;      memory[55226] <=  8'h00;      memory[55227] <=  8'h00;      memory[55228] <=  8'h00;      memory[55229] <=  8'h00;      memory[55230] <=  8'h00;      memory[55231] <=  8'h00;      memory[55232] <=  8'h00;      memory[55233] <=  8'h00;      memory[55234] <=  8'h00;      memory[55235] <=  8'h00;      memory[55236] <=  8'h00;      memory[55237] <=  8'h00;      memory[55238] <=  8'h00;      memory[55239] <=  8'h00;      memory[55240] <=  8'h00;      memory[55241] <=  8'h00;      memory[55242] <=  8'h00;      memory[55243] <=  8'h00;      memory[55244] <=  8'h00;      memory[55245] <=  8'h00;      memory[55246] <=  8'h00;      memory[55247] <=  8'h00;      memory[55248] <=  8'h00;      memory[55249] <=  8'h00;      memory[55250] <=  8'h00;      memory[55251] <=  8'h00;      memory[55252] <=  8'h00;      memory[55253] <=  8'h00;      memory[55254] <=  8'h00;      memory[55255] <=  8'h00;      memory[55256] <=  8'h00;      memory[55257] <=  8'h00;      memory[55258] <=  8'h00;      memory[55259] <=  8'h00;      memory[55260] <=  8'h00;      memory[55261] <=  8'h00;      memory[55262] <=  8'h00;      memory[55263] <=  8'h00;      memory[55264] <=  8'h00;      memory[55265] <=  8'h00;      memory[55266] <=  8'h00;      memory[55267] <=  8'h00;      memory[55268] <=  8'h00;      memory[55269] <=  8'h00;      memory[55270] <=  8'h00;      memory[55271] <=  8'h00;      memory[55272] <=  8'h00;      memory[55273] <=  8'h00;      memory[55274] <=  8'h00;      memory[55275] <=  8'h00;      memory[55276] <=  8'h00;      memory[55277] <=  8'h00;      memory[55278] <=  8'h00;      memory[55279] <=  8'h00;      memory[55280] <=  8'h00;      memory[55281] <=  8'h00;      memory[55282] <=  8'h00;      memory[55283] <=  8'h00;      memory[55284] <=  8'h00;      memory[55285] <=  8'h00;      memory[55286] <=  8'h00;      memory[55287] <=  8'h00;      memory[55288] <=  8'h00;      memory[55289] <=  8'h00;      memory[55290] <=  8'h00;      memory[55291] <=  8'h00;      memory[55292] <=  8'h00;      memory[55293] <=  8'h00;      memory[55294] <=  8'h00;      memory[55295] <=  8'h00;      memory[55296] <=  8'h00;      memory[55297] <=  8'h00;      memory[55298] <=  8'h00;      memory[55299] <=  8'h00;      memory[55300] <=  8'h00;      memory[55301] <=  8'h00;      memory[55302] <=  8'h00;      memory[55303] <=  8'h00;      memory[55304] <=  8'h00;      memory[55305] <=  8'h00;      memory[55306] <=  8'h00;      memory[55307] <=  8'h00;      memory[55308] <=  8'h00;      memory[55309] <=  8'h00;      memory[55310] <=  8'h00;      memory[55311] <=  8'h00;      memory[55312] <=  8'h00;      memory[55313] <=  8'h00;      memory[55314] <=  8'h00;      memory[55315] <=  8'h00;      memory[55316] <=  8'h00;      memory[55317] <=  8'h00;      memory[55318] <=  8'h00;      memory[55319] <=  8'h00;      memory[55320] <=  8'h00;      memory[55321] <=  8'h00;      memory[55322] <=  8'h00;      memory[55323] <=  8'h00;      memory[55324] <=  8'h00;      memory[55325] <=  8'h00;      memory[55326] <=  8'h00;      memory[55327] <=  8'h00;      memory[55328] <=  8'h00;      memory[55329] <=  8'h00;      memory[55330] <=  8'h00;      memory[55331] <=  8'h00;      memory[55332] <=  8'h00;      memory[55333] <=  8'h00;      memory[55334] <=  8'h00;      memory[55335] <=  8'h00;      memory[55336] <=  8'h00;      memory[55337] <=  8'h00;      memory[55338] <=  8'h00;      memory[55339] <=  8'h00;      memory[55340] <=  8'h00;      memory[55341] <=  8'h00;      memory[55342] <=  8'h00;      memory[55343] <=  8'h00;      memory[55344] <=  8'h00;      memory[55345] <=  8'h00;      memory[55346] <=  8'h00;      memory[55347] <=  8'h00;      memory[55348] <=  8'h00;      memory[55349] <=  8'h00;      memory[55350] <=  8'h00;      memory[55351] <=  8'h00;      memory[55352] <=  8'h00;      memory[55353] <=  8'h00;      memory[55354] <=  8'h00;      memory[55355] <=  8'h00;      memory[55356] <=  8'h00;      memory[55357] <=  8'h00;      memory[55358] <=  8'h00;      memory[55359] <=  8'h00;      memory[55360] <=  8'h00;      memory[55361] <=  8'h00;      memory[55362] <=  8'h00;      memory[55363] <=  8'h00;      memory[55364] <=  8'h00;      memory[55365] <=  8'h00;      memory[55366] <=  8'h00;      memory[55367] <=  8'h00;      memory[55368] <=  8'h00;      memory[55369] <=  8'h00;      memory[55370] <=  8'h00;      memory[55371] <=  8'h00;      memory[55372] <=  8'h00;      memory[55373] <=  8'h00;      memory[55374] <=  8'h00;      memory[55375] <=  8'h00;      memory[55376] <=  8'h00;      memory[55377] <=  8'h00;      memory[55378] <=  8'h00;      memory[55379] <=  8'h00;      memory[55380] <=  8'h00;      memory[55381] <=  8'h00;      memory[55382] <=  8'h00;      memory[55383] <=  8'h00;      memory[55384] <=  8'h00;      memory[55385] <=  8'h00;      memory[55386] <=  8'h00;      memory[55387] <=  8'h00;      memory[55388] <=  8'h00;      memory[55389] <=  8'h00;      memory[55390] <=  8'h00;      memory[55391] <=  8'h00;      memory[55392] <=  8'h00;      memory[55393] <=  8'h00;      memory[55394] <=  8'h00;      memory[55395] <=  8'h00;      memory[55396] <=  8'h00;      memory[55397] <=  8'h00;      memory[55398] <=  8'h00;      memory[55399] <=  8'h00;      memory[55400] <=  8'h00;      memory[55401] <=  8'h00;      memory[55402] <=  8'h00;      memory[55403] <=  8'h00;      memory[55404] <=  8'h00;      memory[55405] <=  8'h00;      memory[55406] <=  8'h00;      memory[55407] <=  8'h00;      memory[55408] <=  8'h00;      memory[55409] <=  8'h00;      memory[55410] <=  8'h00;      memory[55411] <=  8'h00;      memory[55412] <=  8'h00;      memory[55413] <=  8'h00;      memory[55414] <=  8'h00;      memory[55415] <=  8'h00;      memory[55416] <=  8'h00;      memory[55417] <=  8'h00;      memory[55418] <=  8'h00;      memory[55419] <=  8'h00;      memory[55420] <=  8'h00;      memory[55421] <=  8'h00;      memory[55422] <=  8'h00;      memory[55423] <=  8'h00;      memory[55424] <=  8'h00;      memory[55425] <=  8'h00;      memory[55426] <=  8'h00;      memory[55427] <=  8'h00;      memory[55428] <=  8'h00;      memory[55429] <=  8'h00;      memory[55430] <=  8'h00;      memory[55431] <=  8'h00;      memory[55432] <=  8'h00;      memory[55433] <=  8'h00;      memory[55434] <=  8'h00;      memory[55435] <=  8'h00;      memory[55436] <=  8'h00;      memory[55437] <=  8'h00;      memory[55438] <=  8'h00;      memory[55439] <=  8'h00;      memory[55440] <=  8'h00;      memory[55441] <=  8'h00;      memory[55442] <=  8'h00;      memory[55443] <=  8'h00;      memory[55444] <=  8'h00;      memory[55445] <=  8'h00;      memory[55446] <=  8'h00;      memory[55447] <=  8'h00;      memory[55448] <=  8'h00;      memory[55449] <=  8'h00;      memory[55450] <=  8'h00;      memory[55451] <=  8'h00;      memory[55452] <=  8'h00;      memory[55453] <=  8'h00;      memory[55454] <=  8'h00;      memory[55455] <=  8'h00;      memory[55456] <=  8'h00;      memory[55457] <=  8'h00;      memory[55458] <=  8'h00;      memory[55459] <=  8'h00;      memory[55460] <=  8'h00;      memory[55461] <=  8'h00;      memory[55462] <=  8'h00;      memory[55463] <=  8'h00;      memory[55464] <=  8'h00;      memory[55465] <=  8'h00;      memory[55466] <=  8'h00;      memory[55467] <=  8'h00;      memory[55468] <=  8'h00;      memory[55469] <=  8'h00;      memory[55470] <=  8'h00;      memory[55471] <=  8'h00;      memory[55472] <=  8'h00;      memory[55473] <=  8'h00;      memory[55474] <=  8'h00;      memory[55475] <=  8'h00;      memory[55476] <=  8'h00;      memory[55477] <=  8'h00;      memory[55478] <=  8'h00;      memory[55479] <=  8'h00;      memory[55480] <=  8'h00;      memory[55481] <=  8'h00;      memory[55482] <=  8'h00;      memory[55483] <=  8'h00;      memory[55484] <=  8'h00;      memory[55485] <=  8'h00;      memory[55486] <=  8'h00;      memory[55487] <=  8'h00;      memory[55488] <=  8'h00;      memory[55489] <=  8'h00;      memory[55490] <=  8'h00;      memory[55491] <=  8'h00;      memory[55492] <=  8'h00;      memory[55493] <=  8'h00;      memory[55494] <=  8'h00;      memory[55495] <=  8'h00;      memory[55496] <=  8'h00;      memory[55497] <=  8'h00;      memory[55498] <=  8'h00;      memory[55499] <=  8'h00;      memory[55500] <=  8'h00;      memory[55501] <=  8'h00;      memory[55502] <=  8'h00;      memory[55503] <=  8'h00;      memory[55504] <=  8'h00;      memory[55505] <=  8'h00;      memory[55506] <=  8'h00;      memory[55507] <=  8'h00;      memory[55508] <=  8'h00;      memory[55509] <=  8'h00;      memory[55510] <=  8'h00;      memory[55511] <=  8'h00;      memory[55512] <=  8'h00;      memory[55513] <=  8'h00;      memory[55514] <=  8'h00;      memory[55515] <=  8'h00;      memory[55516] <=  8'h00;      memory[55517] <=  8'h00;      memory[55518] <=  8'h00;      memory[55519] <=  8'h00;      memory[55520] <=  8'h00;      memory[55521] <=  8'h00;      memory[55522] <=  8'h00;      memory[55523] <=  8'h00;      memory[55524] <=  8'h00;      memory[55525] <=  8'h00;      memory[55526] <=  8'h00;      memory[55527] <=  8'h00;      memory[55528] <=  8'h00;      memory[55529] <=  8'h00;      memory[55530] <=  8'h00;      memory[55531] <=  8'h00;      memory[55532] <=  8'h00;      memory[55533] <=  8'h00;      memory[55534] <=  8'h00;      memory[55535] <=  8'h00;      memory[55536] <=  8'h00;      memory[55537] <=  8'h00;      memory[55538] <=  8'h00;      memory[55539] <=  8'h00;      memory[55540] <=  8'h00;      memory[55541] <=  8'h00;      memory[55542] <=  8'h00;      memory[55543] <=  8'h00;      memory[55544] <=  8'h00;      memory[55545] <=  8'h00;      memory[55546] <=  8'h00;      memory[55547] <=  8'h00;      memory[55548] <=  8'h00;      memory[55549] <=  8'h00;      memory[55550] <=  8'h00;      memory[55551] <=  8'h00;      memory[55552] <=  8'h00;      memory[55553] <=  8'h00;      memory[55554] <=  8'h00;      memory[55555] <=  8'h00;      memory[55556] <=  8'h00;      memory[55557] <=  8'h00;      memory[55558] <=  8'h00;      memory[55559] <=  8'h00;      memory[55560] <=  8'h00;      memory[55561] <=  8'h00;      memory[55562] <=  8'h00;      memory[55563] <=  8'h00;      memory[55564] <=  8'h00;      memory[55565] <=  8'h00;      memory[55566] <=  8'h00;      memory[55567] <=  8'h00;      memory[55568] <=  8'h00;      memory[55569] <=  8'h00;      memory[55570] <=  8'h00;      memory[55571] <=  8'h00;      memory[55572] <=  8'h00;      memory[55573] <=  8'h00;      memory[55574] <=  8'h00;      memory[55575] <=  8'h00;      memory[55576] <=  8'h00;      memory[55577] <=  8'h00;      memory[55578] <=  8'h00;      memory[55579] <=  8'h00;      memory[55580] <=  8'h00;      memory[55581] <=  8'h00;      memory[55582] <=  8'h00;      memory[55583] <=  8'h00;      memory[55584] <=  8'h00;      memory[55585] <=  8'h00;      memory[55586] <=  8'h00;      memory[55587] <=  8'h00;      memory[55588] <=  8'h00;      memory[55589] <=  8'h00;      memory[55590] <=  8'h00;      memory[55591] <=  8'h00;      memory[55592] <=  8'h00;      memory[55593] <=  8'h00;      memory[55594] <=  8'h00;      memory[55595] <=  8'h00;      memory[55596] <=  8'h00;      memory[55597] <=  8'h00;      memory[55598] <=  8'h00;      memory[55599] <=  8'h00;      memory[55600] <=  8'h00;      memory[55601] <=  8'h00;      memory[55602] <=  8'h00;      memory[55603] <=  8'h00;      memory[55604] <=  8'h00;      memory[55605] <=  8'h00;      memory[55606] <=  8'h00;      memory[55607] <=  8'h00;      memory[55608] <=  8'h00;      memory[55609] <=  8'h00;      memory[55610] <=  8'h00;      memory[55611] <=  8'h00;      memory[55612] <=  8'h00;      memory[55613] <=  8'h00;      memory[55614] <=  8'h00;      memory[55615] <=  8'h00;      memory[55616] <=  8'h00;      memory[55617] <=  8'h00;      memory[55618] <=  8'h00;      memory[55619] <=  8'h00;      memory[55620] <=  8'h00;      memory[55621] <=  8'h00;      memory[55622] <=  8'h00;      memory[55623] <=  8'h00;      memory[55624] <=  8'h00;      memory[55625] <=  8'h00;      memory[55626] <=  8'h00;      memory[55627] <=  8'h00;      memory[55628] <=  8'h00;      memory[55629] <=  8'h00;      memory[55630] <=  8'h00;      memory[55631] <=  8'h00;      memory[55632] <=  8'h00;      memory[55633] <=  8'h00;      memory[55634] <=  8'h00;      memory[55635] <=  8'h00;      memory[55636] <=  8'h00;      memory[55637] <=  8'h00;      memory[55638] <=  8'h00;      memory[55639] <=  8'h00;      memory[55640] <=  8'h00;      memory[55641] <=  8'h00;      memory[55642] <=  8'h00;      memory[55643] <=  8'h00;      memory[55644] <=  8'h00;      memory[55645] <=  8'h00;      memory[55646] <=  8'h00;      memory[55647] <=  8'h00;      memory[55648] <=  8'h00;      memory[55649] <=  8'h00;      memory[55650] <=  8'h00;      memory[55651] <=  8'h00;      memory[55652] <=  8'h00;      memory[55653] <=  8'h00;      memory[55654] <=  8'h00;      memory[55655] <=  8'h00;      memory[55656] <=  8'h00;      memory[55657] <=  8'h00;      memory[55658] <=  8'h00;      memory[55659] <=  8'h00;      memory[55660] <=  8'h00;      memory[55661] <=  8'h00;      memory[55662] <=  8'h00;      memory[55663] <=  8'h00;      memory[55664] <=  8'h00;      memory[55665] <=  8'h00;      memory[55666] <=  8'h00;      memory[55667] <=  8'h00;      memory[55668] <=  8'h00;      memory[55669] <=  8'h00;      memory[55670] <=  8'h00;      memory[55671] <=  8'h00;      memory[55672] <=  8'h00;      memory[55673] <=  8'h00;      memory[55674] <=  8'h00;      memory[55675] <=  8'h00;      memory[55676] <=  8'h00;      memory[55677] <=  8'h00;      memory[55678] <=  8'h00;      memory[55679] <=  8'h00;      memory[55680] <=  8'h00;      memory[55681] <=  8'h00;      memory[55682] <=  8'h00;      memory[55683] <=  8'h00;      memory[55684] <=  8'h00;      memory[55685] <=  8'h00;      memory[55686] <=  8'h00;      memory[55687] <=  8'h00;      memory[55688] <=  8'h00;      memory[55689] <=  8'h00;      memory[55690] <=  8'h00;      memory[55691] <=  8'h00;      memory[55692] <=  8'h00;      memory[55693] <=  8'h00;      memory[55694] <=  8'h00;      memory[55695] <=  8'h00;      memory[55696] <=  8'h00;      memory[55697] <=  8'h00;      memory[55698] <=  8'h00;      memory[55699] <=  8'h00;      memory[55700] <=  8'h00;      memory[55701] <=  8'h00;      memory[55702] <=  8'h00;      memory[55703] <=  8'h00;      memory[55704] <=  8'h00;      memory[55705] <=  8'h00;      memory[55706] <=  8'h00;      memory[55707] <=  8'h00;      memory[55708] <=  8'h00;      memory[55709] <=  8'h00;      memory[55710] <=  8'h00;      memory[55711] <=  8'h00;      memory[55712] <=  8'h00;      memory[55713] <=  8'h00;      memory[55714] <=  8'h00;      memory[55715] <=  8'h00;      memory[55716] <=  8'h00;      memory[55717] <=  8'h00;      memory[55718] <=  8'h00;      memory[55719] <=  8'h00;      memory[55720] <=  8'h00;      memory[55721] <=  8'h00;      memory[55722] <=  8'h00;      memory[55723] <=  8'h00;      memory[55724] <=  8'h00;      memory[55725] <=  8'h00;      memory[55726] <=  8'h00;      memory[55727] <=  8'h00;      memory[55728] <=  8'h00;      memory[55729] <=  8'h00;      memory[55730] <=  8'h00;      memory[55731] <=  8'h00;      memory[55732] <=  8'h00;      memory[55733] <=  8'h00;      memory[55734] <=  8'h00;      memory[55735] <=  8'h00;      memory[55736] <=  8'h00;      memory[55737] <=  8'h00;      memory[55738] <=  8'h00;      memory[55739] <=  8'h00;      memory[55740] <=  8'h00;      memory[55741] <=  8'h00;      memory[55742] <=  8'h00;      memory[55743] <=  8'h00;      memory[55744] <=  8'h00;      memory[55745] <=  8'h00;      memory[55746] <=  8'h00;      memory[55747] <=  8'h00;      memory[55748] <=  8'h00;      memory[55749] <=  8'h00;      memory[55750] <=  8'h00;      memory[55751] <=  8'h00;      memory[55752] <=  8'h00;      memory[55753] <=  8'h00;      memory[55754] <=  8'h00;      memory[55755] <=  8'h00;      memory[55756] <=  8'h00;      memory[55757] <=  8'h00;      memory[55758] <=  8'h00;      memory[55759] <=  8'h00;      memory[55760] <=  8'h00;      memory[55761] <=  8'h00;      memory[55762] <=  8'h00;      memory[55763] <=  8'h00;      memory[55764] <=  8'h00;      memory[55765] <=  8'h00;      memory[55766] <=  8'h00;      memory[55767] <=  8'h00;      memory[55768] <=  8'h00;      memory[55769] <=  8'h00;      memory[55770] <=  8'h00;      memory[55771] <=  8'h00;      memory[55772] <=  8'h00;      memory[55773] <=  8'h00;      memory[55774] <=  8'h00;      memory[55775] <=  8'h00;      memory[55776] <=  8'h00;      memory[55777] <=  8'h00;      memory[55778] <=  8'h00;      memory[55779] <=  8'h00;      memory[55780] <=  8'h00;      memory[55781] <=  8'h00;      memory[55782] <=  8'h00;      memory[55783] <=  8'h00;      memory[55784] <=  8'h00;      memory[55785] <=  8'h00;      memory[55786] <=  8'h00;      memory[55787] <=  8'h00;      memory[55788] <=  8'h00;      memory[55789] <=  8'h00;      memory[55790] <=  8'h00;      memory[55791] <=  8'h00;      memory[55792] <=  8'h00;      memory[55793] <=  8'h00;      memory[55794] <=  8'h00;      memory[55795] <=  8'h00;      memory[55796] <=  8'h00;      memory[55797] <=  8'h00;      memory[55798] <=  8'h00;      memory[55799] <=  8'h00;      memory[55800] <=  8'h00;      memory[55801] <=  8'h00;      memory[55802] <=  8'h00;      memory[55803] <=  8'h00;      memory[55804] <=  8'h00;      memory[55805] <=  8'h00;      memory[55806] <=  8'h00;      memory[55807] <=  8'h00;      memory[55808] <=  8'h00;      memory[55809] <=  8'h00;      memory[55810] <=  8'h00;      memory[55811] <=  8'h00;      memory[55812] <=  8'h00;      memory[55813] <=  8'h00;      memory[55814] <=  8'h00;      memory[55815] <=  8'h00;      memory[55816] <=  8'h00;      memory[55817] <=  8'h00;      memory[55818] <=  8'h00;      memory[55819] <=  8'h00;      memory[55820] <=  8'h00;      memory[55821] <=  8'h00;      memory[55822] <=  8'h00;      memory[55823] <=  8'h00;      memory[55824] <=  8'h00;      memory[55825] <=  8'h00;      memory[55826] <=  8'h00;      memory[55827] <=  8'h00;      memory[55828] <=  8'h00;      memory[55829] <=  8'h00;      memory[55830] <=  8'h00;      memory[55831] <=  8'h00;      memory[55832] <=  8'h00;      memory[55833] <=  8'h00;      memory[55834] <=  8'h00;      memory[55835] <=  8'h00;      memory[55836] <=  8'h00;      memory[55837] <=  8'h00;      memory[55838] <=  8'h00;      memory[55839] <=  8'h00;      memory[55840] <=  8'h00;      memory[55841] <=  8'h00;      memory[55842] <=  8'h00;      memory[55843] <=  8'h00;      memory[55844] <=  8'h00;      memory[55845] <=  8'h00;      memory[55846] <=  8'h00;      memory[55847] <=  8'h00;      memory[55848] <=  8'h00;      memory[55849] <=  8'h00;      memory[55850] <=  8'h00;      memory[55851] <=  8'h00;      memory[55852] <=  8'h00;      memory[55853] <=  8'h00;      memory[55854] <=  8'h00;      memory[55855] <=  8'h00;      memory[55856] <=  8'h00;      memory[55857] <=  8'h00;      memory[55858] <=  8'h00;      memory[55859] <=  8'h00;      memory[55860] <=  8'h00;      memory[55861] <=  8'h00;      memory[55862] <=  8'h00;      memory[55863] <=  8'h00;      memory[55864] <=  8'h00;      memory[55865] <=  8'h00;      memory[55866] <=  8'h00;      memory[55867] <=  8'h00;      memory[55868] <=  8'h00;      memory[55869] <=  8'h00;      memory[55870] <=  8'h00;      memory[55871] <=  8'h00;      memory[55872] <=  8'h00;      memory[55873] <=  8'h00;      memory[55874] <=  8'h00;      memory[55875] <=  8'h00;      memory[55876] <=  8'h00;      memory[55877] <=  8'h00;      memory[55878] <=  8'h00;      memory[55879] <=  8'h00;      memory[55880] <=  8'h00;      memory[55881] <=  8'h00;      memory[55882] <=  8'h00;      memory[55883] <=  8'h00;      memory[55884] <=  8'h00;      memory[55885] <=  8'h00;      memory[55886] <=  8'h00;      memory[55887] <=  8'h00;      memory[55888] <=  8'h00;      memory[55889] <=  8'h00;      memory[55890] <=  8'h00;      memory[55891] <=  8'h00;      memory[55892] <=  8'h00;      memory[55893] <=  8'h00;      memory[55894] <=  8'h00;      memory[55895] <=  8'h00;      memory[55896] <=  8'h00;      memory[55897] <=  8'h00;      memory[55898] <=  8'h00;      memory[55899] <=  8'h00;      memory[55900] <=  8'h00;      memory[55901] <=  8'h00;      memory[55902] <=  8'h00;      memory[55903] <=  8'h00;      memory[55904] <=  8'h00;      memory[55905] <=  8'h00;      memory[55906] <=  8'h00;      memory[55907] <=  8'h00;      memory[55908] <=  8'h00;      memory[55909] <=  8'h00;      memory[55910] <=  8'h00;      memory[55911] <=  8'h00;      memory[55912] <=  8'h00;      memory[55913] <=  8'h00;      memory[55914] <=  8'h00;      memory[55915] <=  8'h00;      memory[55916] <=  8'h00;      memory[55917] <=  8'h00;      memory[55918] <=  8'h00;      memory[55919] <=  8'h00;      memory[55920] <=  8'h00;      memory[55921] <=  8'h00;      memory[55922] <=  8'h00;      memory[55923] <=  8'h00;      memory[55924] <=  8'h00;      memory[55925] <=  8'h00;      memory[55926] <=  8'h00;      memory[55927] <=  8'h00;      memory[55928] <=  8'h00;      memory[55929] <=  8'h00;      memory[55930] <=  8'h00;      memory[55931] <=  8'h00;      memory[55932] <=  8'h00;      memory[55933] <=  8'h00;      memory[55934] <=  8'h00;      memory[55935] <=  8'h00;      memory[55936] <=  8'h00;      memory[55937] <=  8'h00;      memory[55938] <=  8'h00;      memory[55939] <=  8'h00;      memory[55940] <=  8'h00;      memory[55941] <=  8'h00;      memory[55942] <=  8'h00;      memory[55943] <=  8'h00;      memory[55944] <=  8'h00;      memory[55945] <=  8'h00;      memory[55946] <=  8'h00;      memory[55947] <=  8'h00;      memory[55948] <=  8'h00;      memory[55949] <=  8'h00;      memory[55950] <=  8'h00;      memory[55951] <=  8'h00;      memory[55952] <=  8'h00;      memory[55953] <=  8'h00;      memory[55954] <=  8'h00;      memory[55955] <=  8'h00;      memory[55956] <=  8'h00;      memory[55957] <=  8'h00;      memory[55958] <=  8'h00;      memory[55959] <=  8'h00;      memory[55960] <=  8'h00;      memory[55961] <=  8'h00;      memory[55962] <=  8'h00;      memory[55963] <=  8'h00;      memory[55964] <=  8'h00;      memory[55965] <=  8'h00;      memory[55966] <=  8'h00;      memory[55967] <=  8'h00;      memory[55968] <=  8'h00;      memory[55969] <=  8'h00;      memory[55970] <=  8'h00;      memory[55971] <=  8'h00;      memory[55972] <=  8'h00;      memory[55973] <=  8'h00;      memory[55974] <=  8'h00;      memory[55975] <=  8'h00;      memory[55976] <=  8'h00;      memory[55977] <=  8'h00;      memory[55978] <=  8'h00;      memory[55979] <=  8'h00;      memory[55980] <=  8'h00;      memory[55981] <=  8'h00;      memory[55982] <=  8'h00;      memory[55983] <=  8'h00;      memory[55984] <=  8'h00;      memory[55985] <=  8'h00;      memory[55986] <=  8'h00;      memory[55987] <=  8'h00;      memory[55988] <=  8'h00;      memory[55989] <=  8'h00;      memory[55990] <=  8'h00;      memory[55991] <=  8'h00;      memory[55992] <=  8'h00;      memory[55993] <=  8'h00;      memory[55994] <=  8'h00;      memory[55995] <=  8'h00;      memory[55996] <=  8'h00;      memory[55997] <=  8'h00;      memory[55998] <=  8'h00;      memory[55999] <=  8'h00;      memory[56000] <=  8'h00;      memory[56001] <=  8'h00;      memory[56002] <=  8'h00;      memory[56003] <=  8'h00;      memory[56004] <=  8'h00;      memory[56005] <=  8'h00;      memory[56006] <=  8'h00;      memory[56007] <=  8'h00;      memory[56008] <=  8'h00;      memory[56009] <=  8'h00;      memory[56010] <=  8'h00;      memory[56011] <=  8'h00;      memory[56012] <=  8'h00;      memory[56013] <=  8'h00;      memory[56014] <=  8'h00;      memory[56015] <=  8'h00;      memory[56016] <=  8'h00;      memory[56017] <=  8'h00;      memory[56018] <=  8'h00;      memory[56019] <=  8'h00;      memory[56020] <=  8'h00;      memory[56021] <=  8'h00;      memory[56022] <=  8'h00;      memory[56023] <=  8'h00;      memory[56024] <=  8'h00;      memory[56025] <=  8'h00;      memory[56026] <=  8'h00;      memory[56027] <=  8'h00;      memory[56028] <=  8'h00;      memory[56029] <=  8'h00;      memory[56030] <=  8'h00;      memory[56031] <=  8'h00;      memory[56032] <=  8'h00;      memory[56033] <=  8'h00;      memory[56034] <=  8'h00;      memory[56035] <=  8'h00;      memory[56036] <=  8'h00;      memory[56037] <=  8'h00;      memory[56038] <=  8'h00;      memory[56039] <=  8'h00;      memory[56040] <=  8'h00;      memory[56041] <=  8'h00;      memory[56042] <=  8'h00;      memory[56043] <=  8'h00;      memory[56044] <=  8'h00;      memory[56045] <=  8'h00;      memory[56046] <=  8'h00;      memory[56047] <=  8'h00;      memory[56048] <=  8'h00;      memory[56049] <=  8'h00;      memory[56050] <=  8'h00;      memory[56051] <=  8'h00;      memory[56052] <=  8'h00;      memory[56053] <=  8'h00;      memory[56054] <=  8'h00;      memory[56055] <=  8'h00;      memory[56056] <=  8'h00;      memory[56057] <=  8'h00;      memory[56058] <=  8'h00;      memory[56059] <=  8'h00;      memory[56060] <=  8'h00;      memory[56061] <=  8'h00;      memory[56062] <=  8'h00;      memory[56063] <=  8'h00;      memory[56064] <=  8'h00;      memory[56065] <=  8'h00;      memory[56066] <=  8'h00;      memory[56067] <=  8'h00;      memory[56068] <=  8'h00;      memory[56069] <=  8'h00;      memory[56070] <=  8'h00;      memory[56071] <=  8'h00;      memory[56072] <=  8'h00;      memory[56073] <=  8'h00;      memory[56074] <=  8'h00;      memory[56075] <=  8'h00;      memory[56076] <=  8'h00;      memory[56077] <=  8'h00;      memory[56078] <=  8'h00;      memory[56079] <=  8'h00;      memory[56080] <=  8'h00;      memory[56081] <=  8'h00;      memory[56082] <=  8'h00;      memory[56083] <=  8'h00;      memory[56084] <=  8'h00;      memory[56085] <=  8'h00;      memory[56086] <=  8'h00;      memory[56087] <=  8'h00;      memory[56088] <=  8'h00;      memory[56089] <=  8'h00;      memory[56090] <=  8'h00;      memory[56091] <=  8'h00;      memory[56092] <=  8'h00;      memory[56093] <=  8'h00;      memory[56094] <=  8'h00;      memory[56095] <=  8'h00;      memory[56096] <=  8'h00;      memory[56097] <=  8'h00;      memory[56098] <=  8'h00;      memory[56099] <=  8'h00;      memory[56100] <=  8'h00;      memory[56101] <=  8'h00;      memory[56102] <=  8'h00;      memory[56103] <=  8'h00;      memory[56104] <=  8'h00;      memory[56105] <=  8'h00;      memory[56106] <=  8'h00;      memory[56107] <=  8'h00;      memory[56108] <=  8'h00;      memory[56109] <=  8'h00;      memory[56110] <=  8'h00;      memory[56111] <=  8'h00;      memory[56112] <=  8'h00;      memory[56113] <=  8'h00;      memory[56114] <=  8'h00;      memory[56115] <=  8'h00;      memory[56116] <=  8'h00;      memory[56117] <=  8'h00;      memory[56118] <=  8'h00;      memory[56119] <=  8'h00;      memory[56120] <=  8'h00;      memory[56121] <=  8'h00;      memory[56122] <=  8'h00;      memory[56123] <=  8'h00;      memory[56124] <=  8'h00;      memory[56125] <=  8'h00;      memory[56126] <=  8'h00;      memory[56127] <=  8'h00;      memory[56128] <=  8'h00;      memory[56129] <=  8'h00;      memory[56130] <=  8'h00;      memory[56131] <=  8'h00;      memory[56132] <=  8'h00;      memory[56133] <=  8'h00;      memory[56134] <=  8'h00;      memory[56135] <=  8'h00;      memory[56136] <=  8'h00;      memory[56137] <=  8'h00;      memory[56138] <=  8'h00;      memory[56139] <=  8'h00;      memory[56140] <=  8'h00;      memory[56141] <=  8'h00;      memory[56142] <=  8'h00;      memory[56143] <=  8'h00;      memory[56144] <=  8'h00;      memory[56145] <=  8'h00;      memory[56146] <=  8'h00;      memory[56147] <=  8'h00;      memory[56148] <=  8'h00;      memory[56149] <=  8'h00;      memory[56150] <=  8'h00;      memory[56151] <=  8'h00;      memory[56152] <=  8'h00;      memory[56153] <=  8'h00;      memory[56154] <=  8'h00;      memory[56155] <=  8'h00;      memory[56156] <=  8'h00;      memory[56157] <=  8'h00;      memory[56158] <=  8'h00;      memory[56159] <=  8'h00;      memory[56160] <=  8'h00;      memory[56161] <=  8'h00;      memory[56162] <=  8'h00;      memory[56163] <=  8'h00;      memory[56164] <=  8'h00;      memory[56165] <=  8'h00;      memory[56166] <=  8'h00;      memory[56167] <=  8'h00;      memory[56168] <=  8'h00;      memory[56169] <=  8'h00;      memory[56170] <=  8'h00;      memory[56171] <=  8'h00;      memory[56172] <=  8'h00;      memory[56173] <=  8'h00;      memory[56174] <=  8'h00;      memory[56175] <=  8'h00;      memory[56176] <=  8'h00;      memory[56177] <=  8'h00;      memory[56178] <=  8'h00;      memory[56179] <=  8'h00;      memory[56180] <=  8'h00;      memory[56181] <=  8'h00;      memory[56182] <=  8'h00;      memory[56183] <=  8'h00;      memory[56184] <=  8'h00;      memory[56185] <=  8'h00;      memory[56186] <=  8'h00;      memory[56187] <=  8'h00;      memory[56188] <=  8'h00;      memory[56189] <=  8'h00;      memory[56190] <=  8'h00;      memory[56191] <=  8'h00;      memory[56192] <=  8'h00;      memory[56193] <=  8'h00;      memory[56194] <=  8'h00;      memory[56195] <=  8'h00;      memory[56196] <=  8'h00;      memory[56197] <=  8'h00;      memory[56198] <=  8'h00;      memory[56199] <=  8'h00;      memory[56200] <=  8'h00;      memory[56201] <=  8'h00;      memory[56202] <=  8'h00;      memory[56203] <=  8'h00;      memory[56204] <=  8'h00;      memory[56205] <=  8'h00;      memory[56206] <=  8'h00;      memory[56207] <=  8'h00;      memory[56208] <=  8'h00;      memory[56209] <=  8'h00;      memory[56210] <=  8'h00;      memory[56211] <=  8'h00;      memory[56212] <=  8'h00;      memory[56213] <=  8'h00;      memory[56214] <=  8'h00;      memory[56215] <=  8'h00;      memory[56216] <=  8'h00;      memory[56217] <=  8'h00;      memory[56218] <=  8'h00;      memory[56219] <=  8'h00;      memory[56220] <=  8'h00;      memory[56221] <=  8'h00;      memory[56222] <=  8'h00;      memory[56223] <=  8'h00;      memory[56224] <=  8'h00;      memory[56225] <=  8'h00;      memory[56226] <=  8'h00;      memory[56227] <=  8'h00;      memory[56228] <=  8'h00;      memory[56229] <=  8'h00;      memory[56230] <=  8'h00;      memory[56231] <=  8'h00;      memory[56232] <=  8'h00;      memory[56233] <=  8'h00;      memory[56234] <=  8'h00;      memory[56235] <=  8'h00;      memory[56236] <=  8'h00;      memory[56237] <=  8'h00;      memory[56238] <=  8'h00;      memory[56239] <=  8'h00;      memory[56240] <=  8'h00;      memory[56241] <=  8'h00;      memory[56242] <=  8'h00;      memory[56243] <=  8'h00;      memory[56244] <=  8'h00;      memory[56245] <=  8'h00;      memory[56246] <=  8'h00;      memory[56247] <=  8'h00;      memory[56248] <=  8'h00;      memory[56249] <=  8'h00;      memory[56250] <=  8'h00;      memory[56251] <=  8'h00;      memory[56252] <=  8'h00;      memory[56253] <=  8'h00;      memory[56254] <=  8'h00;      memory[56255] <=  8'h00;      memory[56256] <=  8'h00;      memory[56257] <=  8'h00;      memory[56258] <=  8'h00;      memory[56259] <=  8'h00;      memory[56260] <=  8'h00;      memory[56261] <=  8'h00;      memory[56262] <=  8'h00;      memory[56263] <=  8'h00;      memory[56264] <=  8'h00;      memory[56265] <=  8'h00;      memory[56266] <=  8'h00;      memory[56267] <=  8'h00;      memory[56268] <=  8'h00;      memory[56269] <=  8'h00;      memory[56270] <=  8'h00;      memory[56271] <=  8'h00;      memory[56272] <=  8'h00;      memory[56273] <=  8'h00;      memory[56274] <=  8'h00;      memory[56275] <=  8'h00;      memory[56276] <=  8'h00;      memory[56277] <=  8'h00;      memory[56278] <=  8'h00;      memory[56279] <=  8'h00;      memory[56280] <=  8'h00;      memory[56281] <=  8'h00;      memory[56282] <=  8'h00;      memory[56283] <=  8'h00;      memory[56284] <=  8'h00;      memory[56285] <=  8'h00;      memory[56286] <=  8'h00;      memory[56287] <=  8'h00;      memory[56288] <=  8'h00;      memory[56289] <=  8'h00;      memory[56290] <=  8'h00;      memory[56291] <=  8'h00;      memory[56292] <=  8'h00;      memory[56293] <=  8'h00;      memory[56294] <=  8'h00;      memory[56295] <=  8'h00;      memory[56296] <=  8'h00;      memory[56297] <=  8'h00;      memory[56298] <=  8'h00;      memory[56299] <=  8'h00;      memory[56300] <=  8'h00;      memory[56301] <=  8'h00;      memory[56302] <=  8'h00;      memory[56303] <=  8'h00;      memory[56304] <=  8'h00;      memory[56305] <=  8'h00;      memory[56306] <=  8'h00;      memory[56307] <=  8'h00;      memory[56308] <=  8'h00;      memory[56309] <=  8'h00;      memory[56310] <=  8'h00;      memory[56311] <=  8'h00;      memory[56312] <=  8'h00;      memory[56313] <=  8'h00;      memory[56314] <=  8'h00;      memory[56315] <=  8'h00;      memory[56316] <=  8'h00;      memory[56317] <=  8'h00;      memory[56318] <=  8'h00;      memory[56319] <=  8'h00;      memory[56320] <=  8'h00;      memory[56321] <=  8'h00;      memory[56322] <=  8'h00;      memory[56323] <=  8'h00;      memory[56324] <=  8'h00;      memory[56325] <=  8'h00;      memory[56326] <=  8'h00;      memory[56327] <=  8'h00;      memory[56328] <=  8'h00;      memory[56329] <=  8'h00;      memory[56330] <=  8'h00;      memory[56331] <=  8'h00;      memory[56332] <=  8'h00;      memory[56333] <=  8'h00;      memory[56334] <=  8'h00;      memory[56335] <=  8'h00;      memory[56336] <=  8'h00;      memory[56337] <=  8'h00;      memory[56338] <=  8'h00;      memory[56339] <=  8'h00;      memory[56340] <=  8'h00;      memory[56341] <=  8'h00;      memory[56342] <=  8'h00;      memory[56343] <=  8'h00;      memory[56344] <=  8'h00;      memory[56345] <=  8'h00;      memory[56346] <=  8'h00;      memory[56347] <=  8'h00;      memory[56348] <=  8'h00;      memory[56349] <=  8'h00;      memory[56350] <=  8'h00;      memory[56351] <=  8'h00;      memory[56352] <=  8'h00;      memory[56353] <=  8'h00;      memory[56354] <=  8'h00;      memory[56355] <=  8'h00;      memory[56356] <=  8'h00;      memory[56357] <=  8'h00;      memory[56358] <=  8'h00;      memory[56359] <=  8'h00;      memory[56360] <=  8'h00;      memory[56361] <=  8'h00;      memory[56362] <=  8'h00;      memory[56363] <=  8'h00;      memory[56364] <=  8'h00;      memory[56365] <=  8'h00;      memory[56366] <=  8'h00;      memory[56367] <=  8'h00;      memory[56368] <=  8'h00;      memory[56369] <=  8'h00;      memory[56370] <=  8'h00;      memory[56371] <=  8'h00;      memory[56372] <=  8'h00;      memory[56373] <=  8'h00;      memory[56374] <=  8'h00;      memory[56375] <=  8'h00;      memory[56376] <=  8'h00;      memory[56377] <=  8'h00;      memory[56378] <=  8'h00;      memory[56379] <=  8'h00;      memory[56380] <=  8'h00;      memory[56381] <=  8'h00;      memory[56382] <=  8'h00;      memory[56383] <=  8'h00;      memory[56384] <=  8'h00;      memory[56385] <=  8'h00;      memory[56386] <=  8'h00;      memory[56387] <=  8'h00;      memory[56388] <=  8'h00;      memory[56389] <=  8'h00;      memory[56390] <=  8'h00;      memory[56391] <=  8'h00;      memory[56392] <=  8'h00;      memory[56393] <=  8'h00;      memory[56394] <=  8'h00;      memory[56395] <=  8'h00;      memory[56396] <=  8'h00;      memory[56397] <=  8'h00;      memory[56398] <=  8'h00;      memory[56399] <=  8'h00;      memory[56400] <=  8'h00;      memory[56401] <=  8'h00;      memory[56402] <=  8'h00;      memory[56403] <=  8'h00;      memory[56404] <=  8'h00;      memory[56405] <=  8'h00;      memory[56406] <=  8'h00;      memory[56407] <=  8'h00;      memory[56408] <=  8'h00;      memory[56409] <=  8'h00;      memory[56410] <=  8'h00;      memory[56411] <=  8'h00;      memory[56412] <=  8'h00;      memory[56413] <=  8'h00;      memory[56414] <=  8'h00;      memory[56415] <=  8'h00;      memory[56416] <=  8'h00;      memory[56417] <=  8'h00;      memory[56418] <=  8'h00;      memory[56419] <=  8'h00;      memory[56420] <=  8'h00;      memory[56421] <=  8'h00;      memory[56422] <=  8'h00;      memory[56423] <=  8'h00;      memory[56424] <=  8'h00;      memory[56425] <=  8'h00;      memory[56426] <=  8'h00;      memory[56427] <=  8'h00;      memory[56428] <=  8'h00;      memory[56429] <=  8'h00;      memory[56430] <=  8'h00;      memory[56431] <=  8'h00;      memory[56432] <=  8'h00;      memory[56433] <=  8'h00;      memory[56434] <=  8'h00;      memory[56435] <=  8'h00;      memory[56436] <=  8'h00;      memory[56437] <=  8'h00;      memory[56438] <=  8'h00;      memory[56439] <=  8'h00;      memory[56440] <=  8'h00;      memory[56441] <=  8'h00;      memory[56442] <=  8'h00;      memory[56443] <=  8'h00;      memory[56444] <=  8'h00;      memory[56445] <=  8'h00;      memory[56446] <=  8'h00;      memory[56447] <=  8'h00;      memory[56448] <=  8'h00;      memory[56449] <=  8'h00;      memory[56450] <=  8'h00;      memory[56451] <=  8'h00;      memory[56452] <=  8'h00;      memory[56453] <=  8'h00;      memory[56454] <=  8'h00;      memory[56455] <=  8'h00;      memory[56456] <=  8'h00;      memory[56457] <=  8'h00;      memory[56458] <=  8'h00;      memory[56459] <=  8'h00;      memory[56460] <=  8'h00;      memory[56461] <=  8'h00;      memory[56462] <=  8'h00;      memory[56463] <=  8'h00;      memory[56464] <=  8'h00;      memory[56465] <=  8'h00;      memory[56466] <=  8'h00;      memory[56467] <=  8'h00;      memory[56468] <=  8'h00;      memory[56469] <=  8'h00;      memory[56470] <=  8'h00;      memory[56471] <=  8'h00;      memory[56472] <=  8'h00;      memory[56473] <=  8'h00;      memory[56474] <=  8'h00;      memory[56475] <=  8'h00;      memory[56476] <=  8'h00;      memory[56477] <=  8'h00;      memory[56478] <=  8'h00;      memory[56479] <=  8'h00;      memory[56480] <=  8'h00;      memory[56481] <=  8'h00;      memory[56482] <=  8'h00;      memory[56483] <=  8'h00;      memory[56484] <=  8'h00;      memory[56485] <=  8'h00;      memory[56486] <=  8'h00;      memory[56487] <=  8'h00;      memory[56488] <=  8'h00;      memory[56489] <=  8'h00;      memory[56490] <=  8'h00;      memory[56491] <=  8'h00;      memory[56492] <=  8'h00;      memory[56493] <=  8'h00;      memory[56494] <=  8'h00;      memory[56495] <=  8'h00;      memory[56496] <=  8'h00;      memory[56497] <=  8'h00;      memory[56498] <=  8'h00;      memory[56499] <=  8'h00;      memory[56500] <=  8'h00;      memory[56501] <=  8'h00;      memory[56502] <=  8'h00;      memory[56503] <=  8'h00;      memory[56504] <=  8'h00;      memory[56505] <=  8'h00;      memory[56506] <=  8'h00;      memory[56507] <=  8'h00;      memory[56508] <=  8'h00;      memory[56509] <=  8'h00;      memory[56510] <=  8'h00;      memory[56511] <=  8'h00;      memory[56512] <=  8'h00;      memory[56513] <=  8'h00;      memory[56514] <=  8'h00;      memory[56515] <=  8'h00;      memory[56516] <=  8'h00;      memory[56517] <=  8'h00;      memory[56518] <=  8'h00;      memory[56519] <=  8'h00;      memory[56520] <=  8'h00;      memory[56521] <=  8'h00;      memory[56522] <=  8'h00;      memory[56523] <=  8'h00;      memory[56524] <=  8'h00;      memory[56525] <=  8'h00;      memory[56526] <=  8'h00;      memory[56527] <=  8'h00;      memory[56528] <=  8'h00;      memory[56529] <=  8'h00;      memory[56530] <=  8'h00;      memory[56531] <=  8'h00;      memory[56532] <=  8'h00;      memory[56533] <=  8'h00;      memory[56534] <=  8'h00;      memory[56535] <=  8'h00;      memory[56536] <=  8'h00;      memory[56537] <=  8'h00;      memory[56538] <=  8'h00;      memory[56539] <=  8'h00;      memory[56540] <=  8'h00;      memory[56541] <=  8'h00;      memory[56542] <=  8'h00;      memory[56543] <=  8'h00;      memory[56544] <=  8'h00;      memory[56545] <=  8'h00;      memory[56546] <=  8'h00;      memory[56547] <=  8'h00;      memory[56548] <=  8'h00;      memory[56549] <=  8'h00;      memory[56550] <=  8'h00;      memory[56551] <=  8'h00;      memory[56552] <=  8'h00;      memory[56553] <=  8'h00;      memory[56554] <=  8'h00;      memory[56555] <=  8'h00;      memory[56556] <=  8'h00;      memory[56557] <=  8'h00;      memory[56558] <=  8'h00;      memory[56559] <=  8'h00;      memory[56560] <=  8'h00;      memory[56561] <=  8'h00;      memory[56562] <=  8'h00;      memory[56563] <=  8'h00;      memory[56564] <=  8'h00;      memory[56565] <=  8'h00;      memory[56566] <=  8'h00;      memory[56567] <=  8'h00;      memory[56568] <=  8'h00;      memory[56569] <=  8'h00;      memory[56570] <=  8'h00;      memory[56571] <=  8'h00;      memory[56572] <=  8'h00;      memory[56573] <=  8'h00;      memory[56574] <=  8'h00;      memory[56575] <=  8'h00;      memory[56576] <=  8'h00;      memory[56577] <=  8'h00;      memory[56578] <=  8'h00;      memory[56579] <=  8'h00;      memory[56580] <=  8'h00;      memory[56581] <=  8'h00;      memory[56582] <=  8'h00;      memory[56583] <=  8'h00;      memory[56584] <=  8'h00;      memory[56585] <=  8'h00;      memory[56586] <=  8'h00;      memory[56587] <=  8'h00;      memory[56588] <=  8'h00;      memory[56589] <=  8'h00;      memory[56590] <=  8'h00;      memory[56591] <=  8'h00;      memory[56592] <=  8'h00;      memory[56593] <=  8'h00;      memory[56594] <=  8'h00;      memory[56595] <=  8'h00;      memory[56596] <=  8'h00;      memory[56597] <=  8'h00;      memory[56598] <=  8'h00;      memory[56599] <=  8'h00;      memory[56600] <=  8'h00;      memory[56601] <=  8'h00;      memory[56602] <=  8'h00;      memory[56603] <=  8'h00;      memory[56604] <=  8'h00;      memory[56605] <=  8'h00;      memory[56606] <=  8'h00;      memory[56607] <=  8'h00;      memory[56608] <=  8'h00;      memory[56609] <=  8'h00;      memory[56610] <=  8'h00;      memory[56611] <=  8'h00;      memory[56612] <=  8'h00;      memory[56613] <=  8'h00;      memory[56614] <=  8'h00;      memory[56615] <=  8'h00;      memory[56616] <=  8'h00;      memory[56617] <=  8'h00;      memory[56618] <=  8'h00;      memory[56619] <=  8'h00;      memory[56620] <=  8'h00;      memory[56621] <=  8'h00;      memory[56622] <=  8'h00;      memory[56623] <=  8'h00;      memory[56624] <=  8'h00;      memory[56625] <=  8'h00;      memory[56626] <=  8'h00;      memory[56627] <=  8'h00;      memory[56628] <=  8'h00;      memory[56629] <=  8'h00;      memory[56630] <=  8'h00;      memory[56631] <=  8'h00;      memory[56632] <=  8'h00;      memory[56633] <=  8'h00;      memory[56634] <=  8'h00;      memory[56635] <=  8'h00;      memory[56636] <=  8'h00;      memory[56637] <=  8'h00;      memory[56638] <=  8'h00;      memory[56639] <=  8'h00;      memory[56640] <=  8'h00;      memory[56641] <=  8'h00;      memory[56642] <=  8'h00;      memory[56643] <=  8'h00;      memory[56644] <=  8'h00;      memory[56645] <=  8'h00;      memory[56646] <=  8'h00;      memory[56647] <=  8'h00;      memory[56648] <=  8'h00;      memory[56649] <=  8'h00;      memory[56650] <=  8'h00;      memory[56651] <=  8'h00;      memory[56652] <=  8'h00;      memory[56653] <=  8'h00;      memory[56654] <=  8'h00;      memory[56655] <=  8'h00;      memory[56656] <=  8'h00;      memory[56657] <=  8'h00;      memory[56658] <=  8'h00;      memory[56659] <=  8'h00;      memory[56660] <=  8'h00;      memory[56661] <=  8'h00;      memory[56662] <=  8'h00;      memory[56663] <=  8'h00;      memory[56664] <=  8'h00;      memory[56665] <=  8'h00;      memory[56666] <=  8'h00;      memory[56667] <=  8'h00;      memory[56668] <=  8'h00;      memory[56669] <=  8'h00;      memory[56670] <=  8'h00;      memory[56671] <=  8'h00;      memory[56672] <=  8'h00;      memory[56673] <=  8'h00;      memory[56674] <=  8'h00;      memory[56675] <=  8'h00;      memory[56676] <=  8'h00;      memory[56677] <=  8'h00;      memory[56678] <=  8'h00;      memory[56679] <=  8'h00;      memory[56680] <=  8'h00;      memory[56681] <=  8'h00;      memory[56682] <=  8'h00;      memory[56683] <=  8'h00;      memory[56684] <=  8'h00;      memory[56685] <=  8'h00;      memory[56686] <=  8'h00;      memory[56687] <=  8'h00;      memory[56688] <=  8'h00;      memory[56689] <=  8'h00;      memory[56690] <=  8'h00;      memory[56691] <=  8'h00;      memory[56692] <=  8'h00;      memory[56693] <=  8'h00;      memory[56694] <=  8'h00;      memory[56695] <=  8'h00;      memory[56696] <=  8'h00;      memory[56697] <=  8'h00;      memory[56698] <=  8'h00;      memory[56699] <=  8'h00;      memory[56700] <=  8'h00;      memory[56701] <=  8'h00;      memory[56702] <=  8'h00;      memory[56703] <=  8'h00;      memory[56704] <=  8'h00;      memory[56705] <=  8'h00;      memory[56706] <=  8'h00;      memory[56707] <=  8'h00;      memory[56708] <=  8'h00;      memory[56709] <=  8'h00;      memory[56710] <=  8'h00;      memory[56711] <=  8'h00;      memory[56712] <=  8'h00;      memory[56713] <=  8'h00;      memory[56714] <=  8'h00;      memory[56715] <=  8'h00;      memory[56716] <=  8'h00;      memory[56717] <=  8'h00;      memory[56718] <=  8'h00;      memory[56719] <=  8'h00;      memory[56720] <=  8'h00;      memory[56721] <=  8'h00;      memory[56722] <=  8'h00;      memory[56723] <=  8'h00;      memory[56724] <=  8'h00;      memory[56725] <=  8'h00;      memory[56726] <=  8'h00;      memory[56727] <=  8'h00;      memory[56728] <=  8'h00;      memory[56729] <=  8'h00;      memory[56730] <=  8'h00;      memory[56731] <=  8'h00;      memory[56732] <=  8'h00;      memory[56733] <=  8'h00;      memory[56734] <=  8'h00;      memory[56735] <=  8'h00;      memory[56736] <=  8'h00;      memory[56737] <=  8'h00;      memory[56738] <=  8'h00;      memory[56739] <=  8'h00;      memory[56740] <=  8'h00;      memory[56741] <=  8'h00;      memory[56742] <=  8'h00;      memory[56743] <=  8'h00;      memory[56744] <=  8'h00;      memory[56745] <=  8'h00;      memory[56746] <=  8'h00;      memory[56747] <=  8'h00;      memory[56748] <=  8'h00;      memory[56749] <=  8'h00;      memory[56750] <=  8'h00;      memory[56751] <=  8'h00;      memory[56752] <=  8'h00;      memory[56753] <=  8'h00;      memory[56754] <=  8'h00;      memory[56755] <=  8'h00;      memory[56756] <=  8'h00;      memory[56757] <=  8'h00;      memory[56758] <=  8'h00;      memory[56759] <=  8'h00;      memory[56760] <=  8'h00;      memory[56761] <=  8'h00;      memory[56762] <=  8'h00;      memory[56763] <=  8'h00;      memory[56764] <=  8'h00;      memory[56765] <=  8'h00;      memory[56766] <=  8'h00;      memory[56767] <=  8'h00;      memory[56768] <=  8'h00;      memory[56769] <=  8'h00;      memory[56770] <=  8'h00;      memory[56771] <=  8'h00;      memory[56772] <=  8'h00;      memory[56773] <=  8'h00;      memory[56774] <=  8'h00;      memory[56775] <=  8'h00;      memory[56776] <=  8'h00;      memory[56777] <=  8'h00;      memory[56778] <=  8'h00;      memory[56779] <=  8'h00;      memory[56780] <=  8'h00;      memory[56781] <=  8'h00;      memory[56782] <=  8'h00;      memory[56783] <=  8'h00;      memory[56784] <=  8'h00;      memory[56785] <=  8'h00;      memory[56786] <=  8'h00;      memory[56787] <=  8'h00;      memory[56788] <=  8'h00;      memory[56789] <=  8'h00;      memory[56790] <=  8'h00;      memory[56791] <=  8'h00;      memory[56792] <=  8'h00;      memory[56793] <=  8'h00;      memory[56794] <=  8'h00;      memory[56795] <=  8'h00;      memory[56796] <=  8'h00;      memory[56797] <=  8'h00;      memory[56798] <=  8'h00;      memory[56799] <=  8'h00;      memory[56800] <=  8'h00;      memory[56801] <=  8'h00;      memory[56802] <=  8'h00;      memory[56803] <=  8'h00;      memory[56804] <=  8'h00;      memory[56805] <=  8'h00;      memory[56806] <=  8'h00;      memory[56807] <=  8'h00;      memory[56808] <=  8'h00;      memory[56809] <=  8'h00;      memory[56810] <=  8'h00;      memory[56811] <=  8'h00;      memory[56812] <=  8'h00;      memory[56813] <=  8'h00;      memory[56814] <=  8'h00;      memory[56815] <=  8'h00;      memory[56816] <=  8'h00;      memory[56817] <=  8'h00;      memory[56818] <=  8'h00;      memory[56819] <=  8'h00;      memory[56820] <=  8'h00;      memory[56821] <=  8'h00;      memory[56822] <=  8'h00;      memory[56823] <=  8'h00;      memory[56824] <=  8'h00;      memory[56825] <=  8'h00;      memory[56826] <=  8'h00;      memory[56827] <=  8'h00;      memory[56828] <=  8'h00;      memory[56829] <=  8'h00;      memory[56830] <=  8'h00;      memory[56831] <=  8'h00;      memory[56832] <=  8'h00;      memory[56833] <=  8'h00;      memory[56834] <=  8'h00;      memory[56835] <=  8'h00;      memory[56836] <=  8'h00;      memory[56837] <=  8'h00;      memory[56838] <=  8'h00;      memory[56839] <=  8'h00;      memory[56840] <=  8'h00;      memory[56841] <=  8'h00;      memory[56842] <=  8'h00;      memory[56843] <=  8'h00;      memory[56844] <=  8'h00;      memory[56845] <=  8'h00;      memory[56846] <=  8'h00;      memory[56847] <=  8'h00;      memory[56848] <=  8'h00;      memory[56849] <=  8'h00;      memory[56850] <=  8'h00;      memory[56851] <=  8'h00;      memory[56852] <=  8'h00;      memory[56853] <=  8'h00;      memory[56854] <=  8'h00;      memory[56855] <=  8'h00;      memory[56856] <=  8'h00;      memory[56857] <=  8'h00;      memory[56858] <=  8'h00;      memory[56859] <=  8'h00;      memory[56860] <=  8'h00;      memory[56861] <=  8'h00;      memory[56862] <=  8'h00;      memory[56863] <=  8'h00;      memory[56864] <=  8'h00;      memory[56865] <=  8'h00;      memory[56866] <=  8'h00;      memory[56867] <=  8'h00;      memory[56868] <=  8'h00;      memory[56869] <=  8'h00;      memory[56870] <=  8'h00;      memory[56871] <=  8'h00;      memory[56872] <=  8'h00;      memory[56873] <=  8'h00;      memory[56874] <=  8'h00;      memory[56875] <=  8'h00;      memory[56876] <=  8'h00;      memory[56877] <=  8'h00;      memory[56878] <=  8'h00;      memory[56879] <=  8'h00;      memory[56880] <=  8'h00;      memory[56881] <=  8'h00;      memory[56882] <=  8'h00;      memory[56883] <=  8'h00;      memory[56884] <=  8'h00;      memory[56885] <=  8'h00;      memory[56886] <=  8'h00;      memory[56887] <=  8'h00;      memory[56888] <=  8'h00;      memory[56889] <=  8'h00;      memory[56890] <=  8'h00;      memory[56891] <=  8'h00;      memory[56892] <=  8'h00;      memory[56893] <=  8'h00;      memory[56894] <=  8'h00;      memory[56895] <=  8'h00;      memory[56896] <=  8'h00;      memory[56897] <=  8'h00;      memory[56898] <=  8'h00;      memory[56899] <=  8'h00;      memory[56900] <=  8'h00;      memory[56901] <=  8'h00;      memory[56902] <=  8'h00;      memory[56903] <=  8'h00;      memory[56904] <=  8'h00;      memory[56905] <=  8'h00;      memory[56906] <=  8'h00;      memory[56907] <=  8'h00;      memory[56908] <=  8'h00;      memory[56909] <=  8'h00;      memory[56910] <=  8'h00;      memory[56911] <=  8'h00;      memory[56912] <=  8'h00;      memory[56913] <=  8'h00;      memory[56914] <=  8'h00;      memory[56915] <=  8'h00;      memory[56916] <=  8'h00;      memory[56917] <=  8'h00;      memory[56918] <=  8'h00;      memory[56919] <=  8'h00;      memory[56920] <=  8'h00;      memory[56921] <=  8'h00;      memory[56922] <=  8'h00;      memory[56923] <=  8'h00;      memory[56924] <=  8'h00;      memory[56925] <=  8'h00;      memory[56926] <=  8'h00;      memory[56927] <=  8'h00;      memory[56928] <=  8'h00;      memory[56929] <=  8'h00;      memory[56930] <=  8'h00;      memory[56931] <=  8'h00;      memory[56932] <=  8'h00;      memory[56933] <=  8'h00;      memory[56934] <=  8'h00;      memory[56935] <=  8'h00;      memory[56936] <=  8'h00;      memory[56937] <=  8'h00;      memory[56938] <=  8'h00;      memory[56939] <=  8'h00;      memory[56940] <=  8'h00;      memory[56941] <=  8'h00;      memory[56942] <=  8'h00;      memory[56943] <=  8'h00;      memory[56944] <=  8'h00;      memory[56945] <=  8'h00;      memory[56946] <=  8'h00;      memory[56947] <=  8'h00;      memory[56948] <=  8'h00;      memory[56949] <=  8'h00;      memory[56950] <=  8'h00;      memory[56951] <=  8'h00;      memory[56952] <=  8'h00;      memory[56953] <=  8'h00;      memory[56954] <=  8'h00;      memory[56955] <=  8'h00;      memory[56956] <=  8'h00;      memory[56957] <=  8'h00;      memory[56958] <=  8'h00;      memory[56959] <=  8'h00;      memory[56960] <=  8'h00;      memory[56961] <=  8'h00;      memory[56962] <=  8'h00;      memory[56963] <=  8'h00;      memory[56964] <=  8'h00;      memory[56965] <=  8'h00;      memory[56966] <=  8'h00;      memory[56967] <=  8'h00;      memory[56968] <=  8'h00;      memory[56969] <=  8'h00;      memory[56970] <=  8'h00;      memory[56971] <=  8'h00;      memory[56972] <=  8'h00;      memory[56973] <=  8'h00;      memory[56974] <=  8'h00;      memory[56975] <=  8'h00;      memory[56976] <=  8'h00;      memory[56977] <=  8'h00;      memory[56978] <=  8'h00;      memory[56979] <=  8'h00;      memory[56980] <=  8'h00;      memory[56981] <=  8'h00;      memory[56982] <=  8'h00;      memory[56983] <=  8'h00;      memory[56984] <=  8'h00;      memory[56985] <=  8'h00;      memory[56986] <=  8'h00;      memory[56987] <=  8'h00;      memory[56988] <=  8'h00;      memory[56989] <=  8'h00;      memory[56990] <=  8'h00;      memory[56991] <=  8'h00;      memory[56992] <=  8'h00;      memory[56993] <=  8'h00;      memory[56994] <=  8'h00;      memory[56995] <=  8'h00;      memory[56996] <=  8'h00;      memory[56997] <=  8'h00;      memory[56998] <=  8'h00;      memory[56999] <=  8'h00;      memory[57000] <=  8'h00;      memory[57001] <=  8'h00;      memory[57002] <=  8'h00;      memory[57003] <=  8'h00;      memory[57004] <=  8'h00;      memory[57005] <=  8'h00;      memory[57006] <=  8'h00;      memory[57007] <=  8'h00;      memory[57008] <=  8'h00;      memory[57009] <=  8'h00;      memory[57010] <=  8'h00;      memory[57011] <=  8'h00;      memory[57012] <=  8'h00;      memory[57013] <=  8'h00;      memory[57014] <=  8'h00;      memory[57015] <=  8'h00;      memory[57016] <=  8'h00;      memory[57017] <=  8'h00;      memory[57018] <=  8'h00;      memory[57019] <=  8'h00;      memory[57020] <=  8'h00;      memory[57021] <=  8'h00;      memory[57022] <=  8'h00;      memory[57023] <=  8'h00;      memory[57024] <=  8'h00;      memory[57025] <=  8'h00;      memory[57026] <=  8'h00;      memory[57027] <=  8'h00;      memory[57028] <=  8'h00;      memory[57029] <=  8'h00;      memory[57030] <=  8'h00;      memory[57031] <=  8'h00;      memory[57032] <=  8'h00;      memory[57033] <=  8'h00;      memory[57034] <=  8'h00;      memory[57035] <=  8'h00;      memory[57036] <=  8'h00;      memory[57037] <=  8'h00;      memory[57038] <=  8'h00;      memory[57039] <=  8'h00;      memory[57040] <=  8'h00;      memory[57041] <=  8'h00;      memory[57042] <=  8'h00;      memory[57043] <=  8'h00;      memory[57044] <=  8'h00;      memory[57045] <=  8'h00;      memory[57046] <=  8'h00;      memory[57047] <=  8'h00;      memory[57048] <=  8'h00;      memory[57049] <=  8'h00;      memory[57050] <=  8'h00;      memory[57051] <=  8'h00;      memory[57052] <=  8'h00;      memory[57053] <=  8'h00;      memory[57054] <=  8'h00;      memory[57055] <=  8'h00;      memory[57056] <=  8'h00;      memory[57057] <=  8'h00;      memory[57058] <=  8'h00;      memory[57059] <=  8'h00;      memory[57060] <=  8'h00;      memory[57061] <=  8'h00;      memory[57062] <=  8'h00;      memory[57063] <=  8'h00;      memory[57064] <=  8'h00;      memory[57065] <=  8'h00;      memory[57066] <=  8'h00;      memory[57067] <=  8'h00;      memory[57068] <=  8'h00;      memory[57069] <=  8'h00;      memory[57070] <=  8'h00;      memory[57071] <=  8'h00;      memory[57072] <=  8'h00;      memory[57073] <=  8'h00;      memory[57074] <=  8'h00;      memory[57075] <=  8'h00;      memory[57076] <=  8'h00;      memory[57077] <=  8'h00;      memory[57078] <=  8'h00;      memory[57079] <=  8'h00;      memory[57080] <=  8'h00;      memory[57081] <=  8'h00;      memory[57082] <=  8'h00;      memory[57083] <=  8'h00;      memory[57084] <=  8'h00;      memory[57085] <=  8'h00;      memory[57086] <=  8'h00;      memory[57087] <=  8'h00;      memory[57088] <=  8'h00;      memory[57089] <=  8'h00;      memory[57090] <=  8'h00;      memory[57091] <=  8'h00;      memory[57092] <=  8'h00;      memory[57093] <=  8'h00;      memory[57094] <=  8'h00;      memory[57095] <=  8'h00;      memory[57096] <=  8'h00;      memory[57097] <=  8'h00;      memory[57098] <=  8'h00;      memory[57099] <=  8'h00;      memory[57100] <=  8'h00;      memory[57101] <=  8'h00;      memory[57102] <=  8'h00;      memory[57103] <=  8'h00;      memory[57104] <=  8'h00;      memory[57105] <=  8'h00;      memory[57106] <=  8'h00;      memory[57107] <=  8'h00;      memory[57108] <=  8'h00;      memory[57109] <=  8'h00;      memory[57110] <=  8'h00;      memory[57111] <=  8'h00;      memory[57112] <=  8'h00;      memory[57113] <=  8'h00;      memory[57114] <=  8'h00;      memory[57115] <=  8'h00;      memory[57116] <=  8'h00;      memory[57117] <=  8'h00;      memory[57118] <=  8'h00;      memory[57119] <=  8'h00;      memory[57120] <=  8'h00;      memory[57121] <=  8'h00;      memory[57122] <=  8'h00;      memory[57123] <=  8'h00;      memory[57124] <=  8'h00;      memory[57125] <=  8'h00;      memory[57126] <=  8'h00;      memory[57127] <=  8'h00;      memory[57128] <=  8'h00;      memory[57129] <=  8'h00;      memory[57130] <=  8'h00;      memory[57131] <=  8'h00;      memory[57132] <=  8'h00;      memory[57133] <=  8'h00;      memory[57134] <=  8'h00;      memory[57135] <=  8'h00;      memory[57136] <=  8'h00;      memory[57137] <=  8'h00;      memory[57138] <=  8'h00;      memory[57139] <=  8'h00;      memory[57140] <=  8'h00;      memory[57141] <=  8'h00;      memory[57142] <=  8'h00;      memory[57143] <=  8'h00;      memory[57144] <=  8'h00;      memory[57145] <=  8'h00;      memory[57146] <=  8'h00;      memory[57147] <=  8'h00;      memory[57148] <=  8'h00;      memory[57149] <=  8'h00;      memory[57150] <=  8'h00;      memory[57151] <=  8'h00;      memory[57152] <=  8'h00;      memory[57153] <=  8'h00;      memory[57154] <=  8'h00;      memory[57155] <=  8'h00;      memory[57156] <=  8'h00;      memory[57157] <=  8'h00;      memory[57158] <=  8'h00;      memory[57159] <=  8'h00;      memory[57160] <=  8'h00;      memory[57161] <=  8'h00;      memory[57162] <=  8'h00;      memory[57163] <=  8'h00;      memory[57164] <=  8'h00;      memory[57165] <=  8'h00;      memory[57166] <=  8'h00;      memory[57167] <=  8'h00;      memory[57168] <=  8'h00;      memory[57169] <=  8'h00;      memory[57170] <=  8'h00;      memory[57171] <=  8'h00;      memory[57172] <=  8'h00;      memory[57173] <=  8'h00;      memory[57174] <=  8'h00;      memory[57175] <=  8'h00;      memory[57176] <=  8'h00;      memory[57177] <=  8'h00;      memory[57178] <=  8'h00;      memory[57179] <=  8'h00;      memory[57180] <=  8'h00;      memory[57181] <=  8'h00;      memory[57182] <=  8'h00;      memory[57183] <=  8'h00;      memory[57184] <=  8'h00;      memory[57185] <=  8'h00;      memory[57186] <=  8'h00;      memory[57187] <=  8'h00;      memory[57188] <=  8'h00;      memory[57189] <=  8'h00;      memory[57190] <=  8'h00;      memory[57191] <=  8'h00;      memory[57192] <=  8'h00;      memory[57193] <=  8'h00;      memory[57194] <=  8'h00;      memory[57195] <=  8'h00;      memory[57196] <=  8'h00;      memory[57197] <=  8'h00;      memory[57198] <=  8'h00;      memory[57199] <=  8'h00;      memory[57200] <=  8'h00;      memory[57201] <=  8'h00;      memory[57202] <=  8'h00;      memory[57203] <=  8'h00;      memory[57204] <=  8'h00;      memory[57205] <=  8'h00;      memory[57206] <=  8'h00;      memory[57207] <=  8'h00;      memory[57208] <=  8'h00;      memory[57209] <=  8'h00;      memory[57210] <=  8'h00;      memory[57211] <=  8'h00;      memory[57212] <=  8'h00;      memory[57213] <=  8'h00;      memory[57214] <=  8'h00;      memory[57215] <=  8'h00;      memory[57216] <=  8'h00;      memory[57217] <=  8'h00;      memory[57218] <=  8'h00;      memory[57219] <=  8'h00;      memory[57220] <=  8'h00;      memory[57221] <=  8'h00;      memory[57222] <=  8'h00;      memory[57223] <=  8'h00;      memory[57224] <=  8'h00;      memory[57225] <=  8'h00;      memory[57226] <=  8'h00;      memory[57227] <=  8'h00;      memory[57228] <=  8'h00;      memory[57229] <=  8'h00;      memory[57230] <=  8'h00;      memory[57231] <=  8'h00;      memory[57232] <=  8'h00;      memory[57233] <=  8'h00;      memory[57234] <=  8'h00;      memory[57235] <=  8'h00;      memory[57236] <=  8'h00;      memory[57237] <=  8'h00;      memory[57238] <=  8'h00;      memory[57239] <=  8'h00;      memory[57240] <=  8'h00;      memory[57241] <=  8'h00;      memory[57242] <=  8'h00;      memory[57243] <=  8'h00;      memory[57244] <=  8'h00;      memory[57245] <=  8'h00;      memory[57246] <=  8'h00;      memory[57247] <=  8'h00;      memory[57248] <=  8'h00;      memory[57249] <=  8'h00;      memory[57250] <=  8'h00;      memory[57251] <=  8'h00;      memory[57252] <=  8'h00;      memory[57253] <=  8'h00;      memory[57254] <=  8'h00;      memory[57255] <=  8'h00;      memory[57256] <=  8'h00;      memory[57257] <=  8'h00;      memory[57258] <=  8'h00;      memory[57259] <=  8'h00;      memory[57260] <=  8'h00;      memory[57261] <=  8'h00;      memory[57262] <=  8'h00;      memory[57263] <=  8'h00;      memory[57264] <=  8'h00;      memory[57265] <=  8'h00;      memory[57266] <=  8'h00;      memory[57267] <=  8'h00;      memory[57268] <=  8'h00;      memory[57269] <=  8'h00;      memory[57270] <=  8'h00;      memory[57271] <=  8'h00;      memory[57272] <=  8'h00;      memory[57273] <=  8'h00;      memory[57274] <=  8'h00;      memory[57275] <=  8'h00;      memory[57276] <=  8'h00;      memory[57277] <=  8'h00;      memory[57278] <=  8'h00;      memory[57279] <=  8'h00;      memory[57280] <=  8'h00;      memory[57281] <=  8'h00;      memory[57282] <=  8'h00;      memory[57283] <=  8'h00;      memory[57284] <=  8'h00;      memory[57285] <=  8'h00;      memory[57286] <=  8'h00;      memory[57287] <=  8'h00;      memory[57288] <=  8'h00;      memory[57289] <=  8'h00;      memory[57290] <=  8'h00;      memory[57291] <=  8'h00;      memory[57292] <=  8'h00;      memory[57293] <=  8'h00;      memory[57294] <=  8'h00;      memory[57295] <=  8'h00;      memory[57296] <=  8'h00;      memory[57297] <=  8'h00;      memory[57298] <=  8'h00;      memory[57299] <=  8'h00;      memory[57300] <=  8'h00;      memory[57301] <=  8'h00;      memory[57302] <=  8'h00;      memory[57303] <=  8'h00;      memory[57304] <=  8'h00;      memory[57305] <=  8'h00;      memory[57306] <=  8'h00;      memory[57307] <=  8'h00;      memory[57308] <=  8'h00;      memory[57309] <=  8'h00;      memory[57310] <=  8'h00;      memory[57311] <=  8'h00;      memory[57312] <=  8'h00;      memory[57313] <=  8'h00;      memory[57314] <=  8'h00;      memory[57315] <=  8'h00;      memory[57316] <=  8'h00;      memory[57317] <=  8'h00;      memory[57318] <=  8'h00;      memory[57319] <=  8'h00;      memory[57320] <=  8'h00;      memory[57321] <=  8'h00;      memory[57322] <=  8'h00;      memory[57323] <=  8'h00;      memory[57324] <=  8'h00;      memory[57325] <=  8'h00;      memory[57326] <=  8'h00;      memory[57327] <=  8'h00;      memory[57328] <=  8'h00;      memory[57329] <=  8'h00;      memory[57330] <=  8'h00;      memory[57331] <=  8'h00;      memory[57332] <=  8'h00;      memory[57333] <=  8'h00;      memory[57334] <=  8'h00;      memory[57335] <=  8'h00;      memory[57336] <=  8'h00;      memory[57337] <=  8'h00;      memory[57338] <=  8'h00;      memory[57339] <=  8'h00;      memory[57340] <=  8'h00;      memory[57341] <=  8'h00;      memory[57342] <=  8'h00;      memory[57343] <=  8'h00;      memory[57344] <=  8'h00;      memory[57345] <=  8'h00;      memory[57346] <=  8'h00;      memory[57347] <=  8'h00;      memory[57348] <=  8'h00;      memory[57349] <=  8'h00;      memory[57350] <=  8'h00;      memory[57351] <=  8'h00;      memory[57352] <=  8'h00;      memory[57353] <=  8'h00;      memory[57354] <=  8'h00;      memory[57355] <=  8'h00;      memory[57356] <=  8'h00;      memory[57357] <=  8'h00;      memory[57358] <=  8'h00;      memory[57359] <=  8'h00;      memory[57360] <=  8'h00;      memory[57361] <=  8'h00;      memory[57362] <=  8'h00;      memory[57363] <=  8'h00;      memory[57364] <=  8'h00;      memory[57365] <=  8'h00;      memory[57366] <=  8'h00;      memory[57367] <=  8'h00;      memory[57368] <=  8'h00;      memory[57369] <=  8'h00;      memory[57370] <=  8'h00;      memory[57371] <=  8'h00;      memory[57372] <=  8'h00;      memory[57373] <=  8'h00;      memory[57374] <=  8'h00;      memory[57375] <=  8'h00;      memory[57376] <=  8'h00;      memory[57377] <=  8'h00;      memory[57378] <=  8'h00;      memory[57379] <=  8'h00;      memory[57380] <=  8'h00;      memory[57381] <=  8'h00;      memory[57382] <=  8'h00;      memory[57383] <=  8'h00;      memory[57384] <=  8'h00;      memory[57385] <=  8'h00;      memory[57386] <=  8'h00;      memory[57387] <=  8'h00;      memory[57388] <=  8'h00;      memory[57389] <=  8'h00;      memory[57390] <=  8'h00;      memory[57391] <=  8'h00;      memory[57392] <=  8'h00;      memory[57393] <=  8'h00;      memory[57394] <=  8'h00;      memory[57395] <=  8'h00;      memory[57396] <=  8'h00;      memory[57397] <=  8'h00;      memory[57398] <=  8'h00;      memory[57399] <=  8'h00;      memory[57400] <=  8'h00;      memory[57401] <=  8'h00;      memory[57402] <=  8'h00;      memory[57403] <=  8'h00;      memory[57404] <=  8'h00;      memory[57405] <=  8'h00;      memory[57406] <=  8'h00;      memory[57407] <=  8'h00;      memory[57408] <=  8'h00;      memory[57409] <=  8'h00;      memory[57410] <=  8'h00;      memory[57411] <=  8'h00;      memory[57412] <=  8'h00;      memory[57413] <=  8'h00;      memory[57414] <=  8'h00;      memory[57415] <=  8'h00;      memory[57416] <=  8'h00;      memory[57417] <=  8'h00;      memory[57418] <=  8'h00;      memory[57419] <=  8'h00;      memory[57420] <=  8'h00;      memory[57421] <=  8'h00;      memory[57422] <=  8'h00;      memory[57423] <=  8'h00;      memory[57424] <=  8'h00;      memory[57425] <=  8'h00;      memory[57426] <=  8'h00;      memory[57427] <=  8'h00;      memory[57428] <=  8'h00;      memory[57429] <=  8'h00;      memory[57430] <=  8'h00;      memory[57431] <=  8'h00;      memory[57432] <=  8'h00;      memory[57433] <=  8'h00;      memory[57434] <=  8'h00;      memory[57435] <=  8'h00;      memory[57436] <=  8'h00;      memory[57437] <=  8'h00;      memory[57438] <=  8'h00;      memory[57439] <=  8'h00;      memory[57440] <=  8'h00;      memory[57441] <=  8'h00;      memory[57442] <=  8'h00;      memory[57443] <=  8'h00;      memory[57444] <=  8'h00;      memory[57445] <=  8'h00;      memory[57446] <=  8'h00;      memory[57447] <=  8'h00;      memory[57448] <=  8'h00;      memory[57449] <=  8'h00;      memory[57450] <=  8'h00;      memory[57451] <=  8'h00;      memory[57452] <=  8'h00;      memory[57453] <=  8'h00;      memory[57454] <=  8'h00;      memory[57455] <=  8'h00;      memory[57456] <=  8'h00;      memory[57457] <=  8'h00;      memory[57458] <=  8'h00;      memory[57459] <=  8'h00;      memory[57460] <=  8'h00;      memory[57461] <=  8'h00;      memory[57462] <=  8'h00;      memory[57463] <=  8'h00;      memory[57464] <=  8'h00;      memory[57465] <=  8'h00;      memory[57466] <=  8'h00;      memory[57467] <=  8'h00;      memory[57468] <=  8'h00;      memory[57469] <=  8'h00;      memory[57470] <=  8'h00;      memory[57471] <=  8'h00;      memory[57472] <=  8'h00;      memory[57473] <=  8'h00;      memory[57474] <=  8'h00;      memory[57475] <=  8'h00;      memory[57476] <=  8'h00;      memory[57477] <=  8'h00;      memory[57478] <=  8'h00;      memory[57479] <=  8'h00;      memory[57480] <=  8'h00;      memory[57481] <=  8'h00;      memory[57482] <=  8'h00;      memory[57483] <=  8'h00;      memory[57484] <=  8'h00;      memory[57485] <=  8'h00;      memory[57486] <=  8'h00;      memory[57487] <=  8'h00;      memory[57488] <=  8'h00;      memory[57489] <=  8'h00;      memory[57490] <=  8'h00;      memory[57491] <=  8'h00;      memory[57492] <=  8'h00;      memory[57493] <=  8'h00;      memory[57494] <=  8'h00;      memory[57495] <=  8'h00;      memory[57496] <=  8'h00;      memory[57497] <=  8'h00;      memory[57498] <=  8'h00;      memory[57499] <=  8'h00;      memory[57500] <=  8'h00;      memory[57501] <=  8'h00;      memory[57502] <=  8'h00;      memory[57503] <=  8'h00;      memory[57504] <=  8'h00;      memory[57505] <=  8'h00;      memory[57506] <=  8'h00;      memory[57507] <=  8'h00;      memory[57508] <=  8'h00;      memory[57509] <=  8'h00;      memory[57510] <=  8'h00;      memory[57511] <=  8'h00;      memory[57512] <=  8'h00;      memory[57513] <=  8'h00;      memory[57514] <=  8'h00;      memory[57515] <=  8'h00;      memory[57516] <=  8'h00;      memory[57517] <=  8'h00;      memory[57518] <=  8'h00;      memory[57519] <=  8'h00;      memory[57520] <=  8'h00;      memory[57521] <=  8'h00;      memory[57522] <=  8'h00;      memory[57523] <=  8'h00;      memory[57524] <=  8'h00;      memory[57525] <=  8'h00;      memory[57526] <=  8'h00;      memory[57527] <=  8'h00;      memory[57528] <=  8'h00;      memory[57529] <=  8'h00;      memory[57530] <=  8'h00;      memory[57531] <=  8'h00;      memory[57532] <=  8'h00;      memory[57533] <=  8'h00;      memory[57534] <=  8'h00;      memory[57535] <=  8'h00;      memory[57536] <=  8'h00;      memory[57537] <=  8'h00;      memory[57538] <=  8'h00;      memory[57539] <=  8'h00;      memory[57540] <=  8'h00;      memory[57541] <=  8'h00;      memory[57542] <=  8'h00;      memory[57543] <=  8'h00;      memory[57544] <=  8'h00;      memory[57545] <=  8'h00;      memory[57546] <=  8'h00;      memory[57547] <=  8'h00;      memory[57548] <=  8'h00;      memory[57549] <=  8'h00;      memory[57550] <=  8'h00;      memory[57551] <=  8'h00;      memory[57552] <=  8'h00;      memory[57553] <=  8'h00;      memory[57554] <=  8'h00;      memory[57555] <=  8'h00;      memory[57556] <=  8'h00;      memory[57557] <=  8'h00;      memory[57558] <=  8'h00;      memory[57559] <=  8'h00;      memory[57560] <=  8'h00;      memory[57561] <=  8'h00;      memory[57562] <=  8'h00;      memory[57563] <=  8'h00;      memory[57564] <=  8'h00;      memory[57565] <=  8'h00;      memory[57566] <=  8'h00;      memory[57567] <=  8'h00;      memory[57568] <=  8'h00;      memory[57569] <=  8'h00;      memory[57570] <=  8'h00;      memory[57571] <=  8'h00;      memory[57572] <=  8'h00;      memory[57573] <=  8'h00;      memory[57574] <=  8'h00;      memory[57575] <=  8'h00;      memory[57576] <=  8'h00;      memory[57577] <=  8'h00;      memory[57578] <=  8'h00;      memory[57579] <=  8'h00;      memory[57580] <=  8'h00;      memory[57581] <=  8'h00;      memory[57582] <=  8'h00;      memory[57583] <=  8'h00;      memory[57584] <=  8'h00;      memory[57585] <=  8'h00;      memory[57586] <=  8'h00;      memory[57587] <=  8'h00;      memory[57588] <=  8'h00;      memory[57589] <=  8'h00;      memory[57590] <=  8'h00;      memory[57591] <=  8'h00;      memory[57592] <=  8'h00;      memory[57593] <=  8'h00;      memory[57594] <=  8'h00;      memory[57595] <=  8'h00;      memory[57596] <=  8'h00;      memory[57597] <=  8'h00;      memory[57598] <=  8'h00;      memory[57599] <=  8'h00;      memory[57600] <=  8'h00;      memory[57601] <=  8'h00;      memory[57602] <=  8'h00;      memory[57603] <=  8'h00;      memory[57604] <=  8'h00;      memory[57605] <=  8'h00;      memory[57606] <=  8'h00;      memory[57607] <=  8'h00;      memory[57608] <=  8'h00;      memory[57609] <=  8'h00;      memory[57610] <=  8'h00;      memory[57611] <=  8'h00;      memory[57612] <=  8'h00;      memory[57613] <=  8'h00;      memory[57614] <=  8'h00;      memory[57615] <=  8'h00;      memory[57616] <=  8'h00;      memory[57617] <=  8'h00;      memory[57618] <=  8'h00;      memory[57619] <=  8'h00;      memory[57620] <=  8'h00;      memory[57621] <=  8'h00;      memory[57622] <=  8'h00;      memory[57623] <=  8'h00;      memory[57624] <=  8'h00;      memory[57625] <=  8'h00;      memory[57626] <=  8'h00;      memory[57627] <=  8'h00;      memory[57628] <=  8'h00;      memory[57629] <=  8'h00;      memory[57630] <=  8'h00;      memory[57631] <=  8'h00;      memory[57632] <=  8'h00;      memory[57633] <=  8'h00;      memory[57634] <=  8'h00;      memory[57635] <=  8'h00;      memory[57636] <=  8'h00;      memory[57637] <=  8'h00;      memory[57638] <=  8'h00;      memory[57639] <=  8'h00;      memory[57640] <=  8'h00;      memory[57641] <=  8'h00;      memory[57642] <=  8'h00;      memory[57643] <=  8'h00;      memory[57644] <=  8'h00;      memory[57645] <=  8'h00;      memory[57646] <=  8'h00;      memory[57647] <=  8'h00;      memory[57648] <=  8'h00;      memory[57649] <=  8'h00;      memory[57650] <=  8'h00;      memory[57651] <=  8'h00;      memory[57652] <=  8'h00;      memory[57653] <=  8'h00;      memory[57654] <=  8'h00;      memory[57655] <=  8'h00;      memory[57656] <=  8'h00;      memory[57657] <=  8'h00;      memory[57658] <=  8'h00;      memory[57659] <=  8'h00;      memory[57660] <=  8'h00;      memory[57661] <=  8'h00;      memory[57662] <=  8'h00;      memory[57663] <=  8'h00;      memory[57664] <=  8'h00;      memory[57665] <=  8'h00;      memory[57666] <=  8'h00;      memory[57667] <=  8'h00;      memory[57668] <=  8'h00;      memory[57669] <=  8'h00;      memory[57670] <=  8'h00;      memory[57671] <=  8'h00;      memory[57672] <=  8'h00;      memory[57673] <=  8'h00;      memory[57674] <=  8'h00;      memory[57675] <=  8'h00;      memory[57676] <=  8'h00;      memory[57677] <=  8'h00;      memory[57678] <=  8'h00;      memory[57679] <=  8'h00;      memory[57680] <=  8'h00;      memory[57681] <=  8'h00;      memory[57682] <=  8'h00;      memory[57683] <=  8'h00;      memory[57684] <=  8'h00;      memory[57685] <=  8'h00;      memory[57686] <=  8'h00;      memory[57687] <=  8'h00;      memory[57688] <=  8'h00;      memory[57689] <=  8'h00;      memory[57690] <=  8'h00;      memory[57691] <=  8'h00;      memory[57692] <=  8'h00;      memory[57693] <=  8'h00;      memory[57694] <=  8'h00;      memory[57695] <=  8'h00;      memory[57696] <=  8'h00;      memory[57697] <=  8'h00;      memory[57698] <=  8'h00;      memory[57699] <=  8'h00;      memory[57700] <=  8'h00;      memory[57701] <=  8'h00;      memory[57702] <=  8'h00;      memory[57703] <=  8'h00;      memory[57704] <=  8'h00;      memory[57705] <=  8'h00;      memory[57706] <=  8'h00;      memory[57707] <=  8'h00;      memory[57708] <=  8'h00;      memory[57709] <=  8'h00;      memory[57710] <=  8'h00;      memory[57711] <=  8'h00;      memory[57712] <=  8'h00;      memory[57713] <=  8'h00;      memory[57714] <=  8'h00;      memory[57715] <=  8'h00;      memory[57716] <=  8'h00;      memory[57717] <=  8'h00;      memory[57718] <=  8'h00;      memory[57719] <=  8'h00;      memory[57720] <=  8'h00;      memory[57721] <=  8'h00;      memory[57722] <=  8'h00;      memory[57723] <=  8'h00;      memory[57724] <=  8'h00;      memory[57725] <=  8'h00;      memory[57726] <=  8'h00;      memory[57727] <=  8'h00;      memory[57728] <=  8'h00;      memory[57729] <=  8'h00;      memory[57730] <=  8'h00;      memory[57731] <=  8'h00;      memory[57732] <=  8'h00;      memory[57733] <=  8'h00;      memory[57734] <=  8'h00;      memory[57735] <=  8'h00;      memory[57736] <=  8'h00;      memory[57737] <=  8'h00;      memory[57738] <=  8'h00;      memory[57739] <=  8'h00;      memory[57740] <=  8'h00;      memory[57741] <=  8'h00;      memory[57742] <=  8'h00;      memory[57743] <=  8'h00;      memory[57744] <=  8'h00;      memory[57745] <=  8'h00;      memory[57746] <=  8'h00;      memory[57747] <=  8'h00;      memory[57748] <=  8'h00;      memory[57749] <=  8'h00;      memory[57750] <=  8'h00;      memory[57751] <=  8'h00;      memory[57752] <=  8'h00;      memory[57753] <=  8'h00;      memory[57754] <=  8'h00;      memory[57755] <=  8'h00;      memory[57756] <=  8'h00;      memory[57757] <=  8'h00;      memory[57758] <=  8'h00;      memory[57759] <=  8'h00;      memory[57760] <=  8'h00;      memory[57761] <=  8'h00;      memory[57762] <=  8'h00;      memory[57763] <=  8'h00;      memory[57764] <=  8'h00;      memory[57765] <=  8'h00;      memory[57766] <=  8'h00;      memory[57767] <=  8'h00;      memory[57768] <=  8'h00;      memory[57769] <=  8'h00;      memory[57770] <=  8'h00;      memory[57771] <=  8'h00;      memory[57772] <=  8'h00;      memory[57773] <=  8'h00;      memory[57774] <=  8'h00;      memory[57775] <=  8'h00;      memory[57776] <=  8'h00;      memory[57777] <=  8'h00;      memory[57778] <=  8'h00;      memory[57779] <=  8'h00;      memory[57780] <=  8'h00;      memory[57781] <=  8'h00;      memory[57782] <=  8'h00;      memory[57783] <=  8'h00;      memory[57784] <=  8'h00;      memory[57785] <=  8'h00;      memory[57786] <=  8'h00;      memory[57787] <=  8'h00;      memory[57788] <=  8'h00;      memory[57789] <=  8'h00;      memory[57790] <=  8'h00;      memory[57791] <=  8'h00;      memory[57792] <=  8'h00;      memory[57793] <=  8'h00;      memory[57794] <=  8'h00;      memory[57795] <=  8'h00;      memory[57796] <=  8'h00;      memory[57797] <=  8'h00;      memory[57798] <=  8'h00;      memory[57799] <=  8'h00;      memory[57800] <=  8'h00;      memory[57801] <=  8'h00;      memory[57802] <=  8'h00;      memory[57803] <=  8'h00;      memory[57804] <=  8'h00;      memory[57805] <=  8'h00;      memory[57806] <=  8'h00;      memory[57807] <=  8'h00;      memory[57808] <=  8'h00;      memory[57809] <=  8'h00;      memory[57810] <=  8'h00;      memory[57811] <=  8'h00;      memory[57812] <=  8'h00;      memory[57813] <=  8'h00;      memory[57814] <=  8'h00;      memory[57815] <=  8'h00;      memory[57816] <=  8'h00;      memory[57817] <=  8'h00;      memory[57818] <=  8'h00;      memory[57819] <=  8'h00;      memory[57820] <=  8'h00;      memory[57821] <=  8'h00;      memory[57822] <=  8'h00;      memory[57823] <=  8'h00;      memory[57824] <=  8'h00;      memory[57825] <=  8'h00;      memory[57826] <=  8'h00;      memory[57827] <=  8'h00;      memory[57828] <=  8'h00;      memory[57829] <=  8'h00;      memory[57830] <=  8'h00;      memory[57831] <=  8'h00;      memory[57832] <=  8'h00;      memory[57833] <=  8'h00;      memory[57834] <=  8'h00;      memory[57835] <=  8'h00;      memory[57836] <=  8'h00;      memory[57837] <=  8'h00;      memory[57838] <=  8'h00;      memory[57839] <=  8'h00;      memory[57840] <=  8'h00;      memory[57841] <=  8'h00;      memory[57842] <=  8'h00;      memory[57843] <=  8'h00;      memory[57844] <=  8'h00;      memory[57845] <=  8'h00;      memory[57846] <=  8'h00;      memory[57847] <=  8'h00;      memory[57848] <=  8'h00;      memory[57849] <=  8'h00;      memory[57850] <=  8'h00;      memory[57851] <=  8'h00;      memory[57852] <=  8'h00;      memory[57853] <=  8'h00;      memory[57854] <=  8'h00;      memory[57855] <=  8'h00;      memory[57856] <=  8'h00;      memory[57857] <=  8'h00;      memory[57858] <=  8'h00;      memory[57859] <=  8'h00;      memory[57860] <=  8'h00;      memory[57861] <=  8'h00;      memory[57862] <=  8'h00;      memory[57863] <=  8'h00;      memory[57864] <=  8'h00;      memory[57865] <=  8'h00;      memory[57866] <=  8'h00;      memory[57867] <=  8'h00;      memory[57868] <=  8'h00;      memory[57869] <=  8'h00;      memory[57870] <=  8'h00;      memory[57871] <=  8'h00;      memory[57872] <=  8'h00;      memory[57873] <=  8'h00;      memory[57874] <=  8'h00;      memory[57875] <=  8'h00;      memory[57876] <=  8'h00;      memory[57877] <=  8'h00;      memory[57878] <=  8'h00;      memory[57879] <=  8'h00;      memory[57880] <=  8'h00;      memory[57881] <=  8'h00;      memory[57882] <=  8'h00;      memory[57883] <=  8'h00;      memory[57884] <=  8'h00;      memory[57885] <=  8'h00;      memory[57886] <=  8'h00;      memory[57887] <=  8'h00;      memory[57888] <=  8'h00;      memory[57889] <=  8'h00;      memory[57890] <=  8'h00;      memory[57891] <=  8'h00;      memory[57892] <=  8'h00;      memory[57893] <=  8'h00;      memory[57894] <=  8'h00;      memory[57895] <=  8'h00;      memory[57896] <=  8'h00;      memory[57897] <=  8'h00;      memory[57898] <=  8'h00;      memory[57899] <=  8'h00;      memory[57900] <=  8'h00;      memory[57901] <=  8'h00;      memory[57902] <=  8'h00;      memory[57903] <=  8'h00;      memory[57904] <=  8'h00;      memory[57905] <=  8'h00;      memory[57906] <=  8'h00;      memory[57907] <=  8'h00;      memory[57908] <=  8'h00;      memory[57909] <=  8'h00;      memory[57910] <=  8'h00;      memory[57911] <=  8'h00;      memory[57912] <=  8'h00;      memory[57913] <=  8'h00;      memory[57914] <=  8'h00;      memory[57915] <=  8'h00;      memory[57916] <=  8'h00;      memory[57917] <=  8'h00;      memory[57918] <=  8'h00;      memory[57919] <=  8'h00;      memory[57920] <=  8'h00;      memory[57921] <=  8'h00;      memory[57922] <=  8'h00;      memory[57923] <=  8'h00;      memory[57924] <=  8'h00;      memory[57925] <=  8'h00;      memory[57926] <=  8'h00;      memory[57927] <=  8'h00;      memory[57928] <=  8'h00;      memory[57929] <=  8'h00;      memory[57930] <=  8'h00;      memory[57931] <=  8'h00;      memory[57932] <=  8'h00;      memory[57933] <=  8'h00;      memory[57934] <=  8'h00;      memory[57935] <=  8'h00;      memory[57936] <=  8'h00;      memory[57937] <=  8'h00;      memory[57938] <=  8'h00;      memory[57939] <=  8'h00;      memory[57940] <=  8'h00;      memory[57941] <=  8'h00;      memory[57942] <=  8'h00;      memory[57943] <=  8'h00;      memory[57944] <=  8'h00;      memory[57945] <=  8'h00;      memory[57946] <=  8'h00;      memory[57947] <=  8'h00;      memory[57948] <=  8'h00;      memory[57949] <=  8'h00;      memory[57950] <=  8'h00;      memory[57951] <=  8'h00;      memory[57952] <=  8'h00;      memory[57953] <=  8'h00;      memory[57954] <=  8'h00;      memory[57955] <=  8'h00;      memory[57956] <=  8'h00;      memory[57957] <=  8'h00;      memory[57958] <=  8'h00;      memory[57959] <=  8'h00;      memory[57960] <=  8'h00;      memory[57961] <=  8'h00;      memory[57962] <=  8'h00;      memory[57963] <=  8'h00;      memory[57964] <=  8'h00;      memory[57965] <=  8'h00;      memory[57966] <=  8'h00;      memory[57967] <=  8'h00;      memory[57968] <=  8'h00;      memory[57969] <=  8'h00;      memory[57970] <=  8'h00;      memory[57971] <=  8'h00;      memory[57972] <=  8'h00;      memory[57973] <=  8'h00;      memory[57974] <=  8'h00;      memory[57975] <=  8'h00;      memory[57976] <=  8'h00;      memory[57977] <=  8'h00;      memory[57978] <=  8'h00;      memory[57979] <=  8'h00;      memory[57980] <=  8'h00;      memory[57981] <=  8'h00;      memory[57982] <=  8'h00;      memory[57983] <=  8'h00;      memory[57984] <=  8'h00;      memory[57985] <=  8'h00;      memory[57986] <=  8'h00;      memory[57987] <=  8'h00;      memory[57988] <=  8'h00;      memory[57989] <=  8'h00;      memory[57990] <=  8'h00;      memory[57991] <=  8'h00;      memory[57992] <=  8'h00;      memory[57993] <=  8'h00;      memory[57994] <=  8'h00;      memory[57995] <=  8'h00;      memory[57996] <=  8'h00;      memory[57997] <=  8'h00;      memory[57998] <=  8'h00;      memory[57999] <=  8'h00;      memory[58000] <=  8'h00;      memory[58001] <=  8'h00;      memory[58002] <=  8'h00;      memory[58003] <=  8'h00;      memory[58004] <=  8'h00;      memory[58005] <=  8'h00;      memory[58006] <=  8'h00;      memory[58007] <=  8'h00;      memory[58008] <=  8'h00;      memory[58009] <=  8'h00;      memory[58010] <=  8'h00;      memory[58011] <=  8'h00;      memory[58012] <=  8'h00;      memory[58013] <=  8'h00;      memory[58014] <=  8'h00;      memory[58015] <=  8'h00;      memory[58016] <=  8'h00;      memory[58017] <=  8'h00;      memory[58018] <=  8'h00;      memory[58019] <=  8'h00;      memory[58020] <=  8'h00;      memory[58021] <=  8'h00;      memory[58022] <=  8'h00;      memory[58023] <=  8'h00;      memory[58024] <=  8'h00;      memory[58025] <=  8'h00;      memory[58026] <=  8'h00;      memory[58027] <=  8'h00;      memory[58028] <=  8'h00;      memory[58029] <=  8'h00;      memory[58030] <=  8'h00;      memory[58031] <=  8'h00;      memory[58032] <=  8'h00;      memory[58033] <=  8'h00;      memory[58034] <=  8'h00;      memory[58035] <=  8'h00;      memory[58036] <=  8'h00;      memory[58037] <=  8'h00;      memory[58038] <=  8'h00;      memory[58039] <=  8'h00;      memory[58040] <=  8'h00;      memory[58041] <=  8'h00;      memory[58042] <=  8'h00;      memory[58043] <=  8'h00;      memory[58044] <=  8'h00;      memory[58045] <=  8'h00;      memory[58046] <=  8'h00;      memory[58047] <=  8'h00;      memory[58048] <=  8'h00;      memory[58049] <=  8'h00;      memory[58050] <=  8'h00;      memory[58051] <=  8'h00;      memory[58052] <=  8'h00;      memory[58053] <=  8'h00;      memory[58054] <=  8'h00;      memory[58055] <=  8'h00;      memory[58056] <=  8'h00;      memory[58057] <=  8'h00;      memory[58058] <=  8'h00;      memory[58059] <=  8'h00;      memory[58060] <=  8'h00;      memory[58061] <=  8'h00;      memory[58062] <=  8'h00;      memory[58063] <=  8'h00;      memory[58064] <=  8'h00;      memory[58065] <=  8'h00;      memory[58066] <=  8'h00;      memory[58067] <=  8'h00;      memory[58068] <=  8'h00;      memory[58069] <=  8'h00;      memory[58070] <=  8'h00;      memory[58071] <=  8'h00;      memory[58072] <=  8'h00;      memory[58073] <=  8'h00;      memory[58074] <=  8'h00;      memory[58075] <=  8'h00;      memory[58076] <=  8'h00;      memory[58077] <=  8'h00;      memory[58078] <=  8'h00;      memory[58079] <=  8'h00;      memory[58080] <=  8'h00;      memory[58081] <=  8'h00;      memory[58082] <=  8'h00;      memory[58083] <=  8'h00;      memory[58084] <=  8'h00;      memory[58085] <=  8'h00;      memory[58086] <=  8'h00;      memory[58087] <=  8'h00;      memory[58088] <=  8'h00;      memory[58089] <=  8'h00;      memory[58090] <=  8'h00;      memory[58091] <=  8'h00;      memory[58092] <=  8'h00;      memory[58093] <=  8'h00;      memory[58094] <=  8'h00;      memory[58095] <=  8'h00;      memory[58096] <=  8'h00;      memory[58097] <=  8'h00;      memory[58098] <=  8'h00;      memory[58099] <=  8'h00;      memory[58100] <=  8'h00;      memory[58101] <=  8'h00;      memory[58102] <=  8'h00;      memory[58103] <=  8'h00;      memory[58104] <=  8'h00;      memory[58105] <=  8'h00;      memory[58106] <=  8'h00;      memory[58107] <=  8'h00;      memory[58108] <=  8'h00;      memory[58109] <=  8'h00;      memory[58110] <=  8'h00;      memory[58111] <=  8'h00;      memory[58112] <=  8'h00;      memory[58113] <=  8'h00;      memory[58114] <=  8'h00;      memory[58115] <=  8'h00;      memory[58116] <=  8'h00;      memory[58117] <=  8'h00;      memory[58118] <=  8'h00;      memory[58119] <=  8'h00;      memory[58120] <=  8'h00;      memory[58121] <=  8'h00;      memory[58122] <=  8'h00;      memory[58123] <=  8'h00;      memory[58124] <=  8'h00;      memory[58125] <=  8'h00;      memory[58126] <=  8'h00;      memory[58127] <=  8'h00;      memory[58128] <=  8'h00;      memory[58129] <=  8'h00;      memory[58130] <=  8'h00;      memory[58131] <=  8'h00;      memory[58132] <=  8'h00;      memory[58133] <=  8'h00;      memory[58134] <=  8'h00;      memory[58135] <=  8'h00;      memory[58136] <=  8'h00;      memory[58137] <=  8'h00;      memory[58138] <=  8'h00;      memory[58139] <=  8'h00;      memory[58140] <=  8'h00;      memory[58141] <=  8'h00;      memory[58142] <=  8'h00;      memory[58143] <=  8'h00;      memory[58144] <=  8'h00;      memory[58145] <=  8'h00;      memory[58146] <=  8'h00;      memory[58147] <=  8'h00;      memory[58148] <=  8'h00;      memory[58149] <=  8'h00;      memory[58150] <=  8'h00;      memory[58151] <=  8'h00;      memory[58152] <=  8'h00;      memory[58153] <=  8'h00;      memory[58154] <=  8'h00;      memory[58155] <=  8'h00;      memory[58156] <=  8'h00;      memory[58157] <=  8'h00;      memory[58158] <=  8'h00;      memory[58159] <=  8'h00;      memory[58160] <=  8'h00;      memory[58161] <=  8'h00;      memory[58162] <=  8'h00;      memory[58163] <=  8'h00;      memory[58164] <=  8'h00;      memory[58165] <=  8'h00;      memory[58166] <=  8'h00;      memory[58167] <=  8'h00;      memory[58168] <=  8'h00;      memory[58169] <=  8'h00;      memory[58170] <=  8'h00;      memory[58171] <=  8'h00;      memory[58172] <=  8'h00;      memory[58173] <=  8'h00;      memory[58174] <=  8'h00;      memory[58175] <=  8'h00;      memory[58176] <=  8'h00;      memory[58177] <=  8'h00;      memory[58178] <=  8'h00;      memory[58179] <=  8'h00;      memory[58180] <=  8'h00;      memory[58181] <=  8'h00;      memory[58182] <=  8'h00;      memory[58183] <=  8'h00;      memory[58184] <=  8'h00;      memory[58185] <=  8'h00;      memory[58186] <=  8'h00;      memory[58187] <=  8'h00;      memory[58188] <=  8'h00;      memory[58189] <=  8'h00;      memory[58190] <=  8'h00;      memory[58191] <=  8'h00;      memory[58192] <=  8'h00;      memory[58193] <=  8'h00;      memory[58194] <=  8'h00;      memory[58195] <=  8'h00;      memory[58196] <=  8'h00;      memory[58197] <=  8'h00;      memory[58198] <=  8'h00;      memory[58199] <=  8'h00;      memory[58200] <=  8'h00;      memory[58201] <=  8'h00;      memory[58202] <=  8'h00;      memory[58203] <=  8'h00;      memory[58204] <=  8'h00;      memory[58205] <=  8'h00;      memory[58206] <=  8'h00;      memory[58207] <=  8'h00;      memory[58208] <=  8'h00;      memory[58209] <=  8'h00;      memory[58210] <=  8'h00;      memory[58211] <=  8'h00;      memory[58212] <=  8'h00;      memory[58213] <=  8'h00;      memory[58214] <=  8'h00;      memory[58215] <=  8'h00;      memory[58216] <=  8'h00;      memory[58217] <=  8'h00;      memory[58218] <=  8'h00;      memory[58219] <=  8'h00;      memory[58220] <=  8'h00;      memory[58221] <=  8'h00;      memory[58222] <=  8'h00;      memory[58223] <=  8'h00;      memory[58224] <=  8'h00;      memory[58225] <=  8'h00;      memory[58226] <=  8'h00;      memory[58227] <=  8'h00;      memory[58228] <=  8'h00;      memory[58229] <=  8'h00;      memory[58230] <=  8'h00;      memory[58231] <=  8'h00;      memory[58232] <=  8'h00;      memory[58233] <=  8'h00;      memory[58234] <=  8'h00;      memory[58235] <=  8'h00;      memory[58236] <=  8'h00;      memory[58237] <=  8'h00;      memory[58238] <=  8'h00;      memory[58239] <=  8'h00;      memory[58240] <=  8'h00;      memory[58241] <=  8'h00;      memory[58242] <=  8'h00;      memory[58243] <=  8'h00;      memory[58244] <=  8'h00;      memory[58245] <=  8'h00;      memory[58246] <=  8'h00;      memory[58247] <=  8'h00;      memory[58248] <=  8'h00;      memory[58249] <=  8'h00;      memory[58250] <=  8'h00;      memory[58251] <=  8'h00;      memory[58252] <=  8'h00;      memory[58253] <=  8'h00;      memory[58254] <=  8'h00;      memory[58255] <=  8'h00;      memory[58256] <=  8'h00;      memory[58257] <=  8'h00;      memory[58258] <=  8'h00;      memory[58259] <=  8'h00;      memory[58260] <=  8'h00;      memory[58261] <=  8'h00;      memory[58262] <=  8'h00;      memory[58263] <=  8'h00;      memory[58264] <=  8'h00;      memory[58265] <=  8'h00;      memory[58266] <=  8'h00;      memory[58267] <=  8'h00;      memory[58268] <=  8'h00;      memory[58269] <=  8'h00;      memory[58270] <=  8'h00;      memory[58271] <=  8'h00;      memory[58272] <=  8'h00;      memory[58273] <=  8'h00;      memory[58274] <=  8'h00;      memory[58275] <=  8'h00;      memory[58276] <=  8'h00;      memory[58277] <=  8'h00;      memory[58278] <=  8'h00;      memory[58279] <=  8'h00;      memory[58280] <=  8'h00;      memory[58281] <=  8'h00;      memory[58282] <=  8'h00;      memory[58283] <=  8'h00;      memory[58284] <=  8'h00;      memory[58285] <=  8'h00;      memory[58286] <=  8'h00;      memory[58287] <=  8'h00;      memory[58288] <=  8'h00;      memory[58289] <=  8'h00;      memory[58290] <=  8'h00;      memory[58291] <=  8'h00;      memory[58292] <=  8'h00;      memory[58293] <=  8'h00;      memory[58294] <=  8'h00;      memory[58295] <=  8'h00;      memory[58296] <=  8'h00;      memory[58297] <=  8'h00;      memory[58298] <=  8'h00;      memory[58299] <=  8'h00;      memory[58300] <=  8'h00;      memory[58301] <=  8'h00;      memory[58302] <=  8'h00;      memory[58303] <=  8'h00;      memory[58304] <=  8'h00;      memory[58305] <=  8'h00;      memory[58306] <=  8'h00;      memory[58307] <=  8'h00;      memory[58308] <=  8'h00;      memory[58309] <=  8'h00;      memory[58310] <=  8'h00;      memory[58311] <=  8'h00;      memory[58312] <=  8'h00;      memory[58313] <=  8'h00;      memory[58314] <=  8'h00;      memory[58315] <=  8'h00;      memory[58316] <=  8'h00;      memory[58317] <=  8'h00;      memory[58318] <=  8'h00;      memory[58319] <=  8'h00;      memory[58320] <=  8'h00;      memory[58321] <=  8'h00;      memory[58322] <=  8'h00;      memory[58323] <=  8'h00;      memory[58324] <=  8'h00;      memory[58325] <=  8'h00;      memory[58326] <=  8'h00;      memory[58327] <=  8'h00;      memory[58328] <=  8'h00;      memory[58329] <=  8'h00;      memory[58330] <=  8'h00;      memory[58331] <=  8'h00;      memory[58332] <=  8'h00;      memory[58333] <=  8'h00;      memory[58334] <=  8'h00;      memory[58335] <=  8'h00;      memory[58336] <=  8'h00;      memory[58337] <=  8'h00;      memory[58338] <=  8'h00;      memory[58339] <=  8'h00;      memory[58340] <=  8'h00;      memory[58341] <=  8'h00;      memory[58342] <=  8'h00;      memory[58343] <=  8'h00;      memory[58344] <=  8'h00;      memory[58345] <=  8'h00;      memory[58346] <=  8'h00;      memory[58347] <=  8'h00;      memory[58348] <=  8'h00;      memory[58349] <=  8'h00;      memory[58350] <=  8'h00;      memory[58351] <=  8'h00;      memory[58352] <=  8'h00;      memory[58353] <=  8'h00;      memory[58354] <=  8'h00;      memory[58355] <=  8'h00;      memory[58356] <=  8'h00;      memory[58357] <=  8'h00;      memory[58358] <=  8'h00;      memory[58359] <=  8'h00;      memory[58360] <=  8'h00;      memory[58361] <=  8'h00;      memory[58362] <=  8'h00;      memory[58363] <=  8'h00;      memory[58364] <=  8'h00;      memory[58365] <=  8'h00;      memory[58366] <=  8'h00;      memory[58367] <=  8'h00;      memory[58368] <=  8'h00;      memory[58369] <=  8'h00;      memory[58370] <=  8'h00;      memory[58371] <=  8'h00;      memory[58372] <=  8'h00;      memory[58373] <=  8'h00;      memory[58374] <=  8'h00;      memory[58375] <=  8'h00;      memory[58376] <=  8'h00;      memory[58377] <=  8'h00;      memory[58378] <=  8'h00;      memory[58379] <=  8'h00;      memory[58380] <=  8'h00;      memory[58381] <=  8'h00;      memory[58382] <=  8'h00;      memory[58383] <=  8'h00;      memory[58384] <=  8'h00;      memory[58385] <=  8'h00;      memory[58386] <=  8'h00;      memory[58387] <=  8'h00;      memory[58388] <=  8'h00;      memory[58389] <=  8'h00;      memory[58390] <=  8'h00;      memory[58391] <=  8'h00;      memory[58392] <=  8'h00;      memory[58393] <=  8'h00;      memory[58394] <=  8'h00;      memory[58395] <=  8'h00;      memory[58396] <=  8'h00;      memory[58397] <=  8'h00;      memory[58398] <=  8'h00;      memory[58399] <=  8'h00;      memory[58400] <=  8'h00;      memory[58401] <=  8'h00;      memory[58402] <=  8'h00;      memory[58403] <=  8'h00;      memory[58404] <=  8'h00;      memory[58405] <=  8'h00;      memory[58406] <=  8'h00;      memory[58407] <=  8'h00;      memory[58408] <=  8'h00;      memory[58409] <=  8'h00;      memory[58410] <=  8'h00;      memory[58411] <=  8'h00;      memory[58412] <=  8'h00;      memory[58413] <=  8'h00;      memory[58414] <=  8'h00;      memory[58415] <=  8'h00;      memory[58416] <=  8'h00;      memory[58417] <=  8'h00;      memory[58418] <=  8'h00;      memory[58419] <=  8'h00;      memory[58420] <=  8'h00;      memory[58421] <=  8'h00;      memory[58422] <=  8'h00;      memory[58423] <=  8'h00;      memory[58424] <=  8'h00;      memory[58425] <=  8'h00;      memory[58426] <=  8'h00;      memory[58427] <=  8'h00;      memory[58428] <=  8'h00;      memory[58429] <=  8'h00;      memory[58430] <=  8'h00;      memory[58431] <=  8'h00;      memory[58432] <=  8'h00;      memory[58433] <=  8'h00;      memory[58434] <=  8'h00;      memory[58435] <=  8'h00;      memory[58436] <=  8'h00;      memory[58437] <=  8'h00;      memory[58438] <=  8'h00;      memory[58439] <=  8'h00;      memory[58440] <=  8'h00;      memory[58441] <=  8'h00;      memory[58442] <=  8'h00;      memory[58443] <=  8'h00;      memory[58444] <=  8'h00;      memory[58445] <=  8'h00;      memory[58446] <=  8'h00;      memory[58447] <=  8'h00;      memory[58448] <=  8'h00;      memory[58449] <=  8'h00;      memory[58450] <=  8'h00;      memory[58451] <=  8'h00;      memory[58452] <=  8'h00;      memory[58453] <=  8'h00;      memory[58454] <=  8'h00;      memory[58455] <=  8'h00;      memory[58456] <=  8'h00;      memory[58457] <=  8'h00;      memory[58458] <=  8'h00;      memory[58459] <=  8'h00;      memory[58460] <=  8'h00;      memory[58461] <=  8'h00;      memory[58462] <=  8'h00;      memory[58463] <=  8'h00;      memory[58464] <=  8'h00;      memory[58465] <=  8'h00;      memory[58466] <=  8'h00;      memory[58467] <=  8'h00;      memory[58468] <=  8'h00;      memory[58469] <=  8'h00;      memory[58470] <=  8'h00;      memory[58471] <=  8'h00;      memory[58472] <=  8'h00;      memory[58473] <=  8'h00;      memory[58474] <=  8'h00;      memory[58475] <=  8'h00;      memory[58476] <=  8'h00;      memory[58477] <=  8'h00;      memory[58478] <=  8'h00;      memory[58479] <=  8'h00;      memory[58480] <=  8'h00;      memory[58481] <=  8'h00;      memory[58482] <=  8'h00;      memory[58483] <=  8'h00;      memory[58484] <=  8'h00;      memory[58485] <=  8'h00;      memory[58486] <=  8'h00;      memory[58487] <=  8'h00;      memory[58488] <=  8'h00;      memory[58489] <=  8'h00;      memory[58490] <=  8'h00;      memory[58491] <=  8'h00;      memory[58492] <=  8'h00;      memory[58493] <=  8'h00;      memory[58494] <=  8'h00;      memory[58495] <=  8'h00;      memory[58496] <=  8'h00;      memory[58497] <=  8'h00;      memory[58498] <=  8'h00;      memory[58499] <=  8'h00;      memory[58500] <=  8'h00;      memory[58501] <=  8'h00;      memory[58502] <=  8'h00;      memory[58503] <=  8'h00;      memory[58504] <=  8'h00;      memory[58505] <=  8'h00;      memory[58506] <=  8'h00;      memory[58507] <=  8'h00;      memory[58508] <=  8'h00;      memory[58509] <=  8'h00;      memory[58510] <=  8'h00;      memory[58511] <=  8'h00;      memory[58512] <=  8'h00;      memory[58513] <=  8'h00;      memory[58514] <=  8'h00;      memory[58515] <=  8'h00;      memory[58516] <=  8'h00;      memory[58517] <=  8'h00;      memory[58518] <=  8'h00;      memory[58519] <=  8'h00;      memory[58520] <=  8'h00;      memory[58521] <=  8'h00;      memory[58522] <=  8'h00;      memory[58523] <=  8'h00;      memory[58524] <=  8'h00;      memory[58525] <=  8'h00;      memory[58526] <=  8'h00;      memory[58527] <=  8'h00;      memory[58528] <=  8'h00;      memory[58529] <=  8'h00;      memory[58530] <=  8'h00;      memory[58531] <=  8'h00;      memory[58532] <=  8'h00;      memory[58533] <=  8'h00;      memory[58534] <=  8'h00;      memory[58535] <=  8'h00;      memory[58536] <=  8'h00;      memory[58537] <=  8'h00;      memory[58538] <=  8'h00;      memory[58539] <=  8'h00;      memory[58540] <=  8'h00;      memory[58541] <=  8'h00;      memory[58542] <=  8'h00;      memory[58543] <=  8'h00;      memory[58544] <=  8'h00;      memory[58545] <=  8'h00;      memory[58546] <=  8'h00;      memory[58547] <=  8'h00;      memory[58548] <=  8'h00;      memory[58549] <=  8'h00;      memory[58550] <=  8'h00;      memory[58551] <=  8'h00;      memory[58552] <=  8'h00;      memory[58553] <=  8'h00;      memory[58554] <=  8'h00;      memory[58555] <=  8'h00;      memory[58556] <=  8'h00;      memory[58557] <=  8'h00;      memory[58558] <=  8'h00;      memory[58559] <=  8'h00;      memory[58560] <=  8'h00;      memory[58561] <=  8'h00;      memory[58562] <=  8'h00;      memory[58563] <=  8'h00;      memory[58564] <=  8'h00;      memory[58565] <=  8'h00;      memory[58566] <=  8'h00;      memory[58567] <=  8'h00;      memory[58568] <=  8'h00;      memory[58569] <=  8'h00;      memory[58570] <=  8'h00;      memory[58571] <=  8'h00;      memory[58572] <=  8'h00;      memory[58573] <=  8'h00;      memory[58574] <=  8'h00;      memory[58575] <=  8'h00;      memory[58576] <=  8'h00;      memory[58577] <=  8'h00;      memory[58578] <=  8'h00;      memory[58579] <=  8'h00;      memory[58580] <=  8'h00;      memory[58581] <=  8'h00;      memory[58582] <=  8'h00;      memory[58583] <=  8'h00;      memory[58584] <=  8'h00;      memory[58585] <=  8'h00;      memory[58586] <=  8'h00;      memory[58587] <=  8'h00;      memory[58588] <=  8'h00;      memory[58589] <=  8'h00;      memory[58590] <=  8'h00;      memory[58591] <=  8'h00;      memory[58592] <=  8'h00;      memory[58593] <=  8'h00;      memory[58594] <=  8'h00;      memory[58595] <=  8'h00;      memory[58596] <=  8'h00;      memory[58597] <=  8'h00;      memory[58598] <=  8'h00;      memory[58599] <=  8'h00;      memory[58600] <=  8'h00;      memory[58601] <=  8'h00;      memory[58602] <=  8'h00;      memory[58603] <=  8'h00;      memory[58604] <=  8'h00;      memory[58605] <=  8'h00;      memory[58606] <=  8'h00;      memory[58607] <=  8'h00;      memory[58608] <=  8'h00;      memory[58609] <=  8'h00;      memory[58610] <=  8'h00;      memory[58611] <=  8'h00;      memory[58612] <=  8'h00;      memory[58613] <=  8'h00;      memory[58614] <=  8'h00;      memory[58615] <=  8'h00;      memory[58616] <=  8'h00;      memory[58617] <=  8'h00;      memory[58618] <=  8'h00;      memory[58619] <=  8'h00;      memory[58620] <=  8'h00;      memory[58621] <=  8'h00;      memory[58622] <=  8'h00;      memory[58623] <=  8'h00;      memory[58624] <=  8'h00;      memory[58625] <=  8'h00;      memory[58626] <=  8'h00;      memory[58627] <=  8'h00;      memory[58628] <=  8'h00;      memory[58629] <=  8'h00;      memory[58630] <=  8'h00;      memory[58631] <=  8'h00;      memory[58632] <=  8'h00;      memory[58633] <=  8'h00;      memory[58634] <=  8'h00;      memory[58635] <=  8'h00;      memory[58636] <=  8'h00;      memory[58637] <=  8'h00;      memory[58638] <=  8'h00;      memory[58639] <=  8'h00;      memory[58640] <=  8'h00;      memory[58641] <=  8'h00;      memory[58642] <=  8'h00;      memory[58643] <=  8'h00;      memory[58644] <=  8'h00;      memory[58645] <=  8'h00;      memory[58646] <=  8'h00;      memory[58647] <=  8'h00;      memory[58648] <=  8'h00;      memory[58649] <=  8'h00;      memory[58650] <=  8'h00;      memory[58651] <=  8'h00;      memory[58652] <=  8'h00;      memory[58653] <=  8'h00;      memory[58654] <=  8'h00;      memory[58655] <=  8'h00;      memory[58656] <=  8'h00;      memory[58657] <=  8'h00;      memory[58658] <=  8'h00;      memory[58659] <=  8'h00;      memory[58660] <=  8'h00;      memory[58661] <=  8'h00;      memory[58662] <=  8'h00;      memory[58663] <=  8'h00;      memory[58664] <=  8'h00;      memory[58665] <=  8'h00;      memory[58666] <=  8'h00;      memory[58667] <=  8'h00;      memory[58668] <=  8'h00;      memory[58669] <=  8'h00;      memory[58670] <=  8'h00;      memory[58671] <=  8'h00;      memory[58672] <=  8'h00;      memory[58673] <=  8'h00;      memory[58674] <=  8'h00;      memory[58675] <=  8'h00;      memory[58676] <=  8'h00;      memory[58677] <=  8'h00;      memory[58678] <=  8'h00;      memory[58679] <=  8'h00;      memory[58680] <=  8'h00;      memory[58681] <=  8'h00;      memory[58682] <=  8'h00;      memory[58683] <=  8'h00;      memory[58684] <=  8'h00;      memory[58685] <=  8'h00;      memory[58686] <=  8'h00;      memory[58687] <=  8'h00;      memory[58688] <=  8'h00;      memory[58689] <=  8'h00;      memory[58690] <=  8'h00;      memory[58691] <=  8'h00;      memory[58692] <=  8'h00;      memory[58693] <=  8'h00;      memory[58694] <=  8'h00;      memory[58695] <=  8'h00;      memory[58696] <=  8'h00;      memory[58697] <=  8'h00;      memory[58698] <=  8'h00;      memory[58699] <=  8'h00;      memory[58700] <=  8'h00;      memory[58701] <=  8'h00;      memory[58702] <=  8'h00;      memory[58703] <=  8'h00;      memory[58704] <=  8'h00;      memory[58705] <=  8'h00;      memory[58706] <=  8'h00;      memory[58707] <=  8'h00;      memory[58708] <=  8'h00;      memory[58709] <=  8'h00;      memory[58710] <=  8'h00;      memory[58711] <=  8'h00;      memory[58712] <=  8'h00;      memory[58713] <=  8'h00;      memory[58714] <=  8'h00;      memory[58715] <=  8'h00;      memory[58716] <=  8'h00;      memory[58717] <=  8'h00;      memory[58718] <=  8'h00;      memory[58719] <=  8'h00;      memory[58720] <=  8'h00;      memory[58721] <=  8'h00;      memory[58722] <=  8'h00;      memory[58723] <=  8'h00;      memory[58724] <=  8'h00;      memory[58725] <=  8'h00;      memory[58726] <=  8'h00;      memory[58727] <=  8'h00;      memory[58728] <=  8'h00;      memory[58729] <=  8'h00;      memory[58730] <=  8'h00;      memory[58731] <=  8'h00;      memory[58732] <=  8'h00;      memory[58733] <=  8'h00;      memory[58734] <=  8'h00;      memory[58735] <=  8'h00;      memory[58736] <=  8'h00;      memory[58737] <=  8'h00;      memory[58738] <=  8'h00;      memory[58739] <=  8'h00;      memory[58740] <=  8'h00;      memory[58741] <=  8'h00;      memory[58742] <=  8'h00;      memory[58743] <=  8'h00;      memory[58744] <=  8'h00;      memory[58745] <=  8'h00;      memory[58746] <=  8'h00;      memory[58747] <=  8'h00;      memory[58748] <=  8'h00;      memory[58749] <=  8'h00;      memory[58750] <=  8'h00;      memory[58751] <=  8'h00;      memory[58752] <=  8'h00;      memory[58753] <=  8'h00;      memory[58754] <=  8'h00;      memory[58755] <=  8'h00;      memory[58756] <=  8'h00;      memory[58757] <=  8'h00;      memory[58758] <=  8'h00;      memory[58759] <=  8'h00;      memory[58760] <=  8'h00;      memory[58761] <=  8'h00;      memory[58762] <=  8'h00;      memory[58763] <=  8'h00;      memory[58764] <=  8'h00;      memory[58765] <=  8'h00;      memory[58766] <=  8'h00;      memory[58767] <=  8'h00;      memory[58768] <=  8'h00;      memory[58769] <=  8'h00;      memory[58770] <=  8'h00;      memory[58771] <=  8'h00;      memory[58772] <=  8'h00;      memory[58773] <=  8'h00;      memory[58774] <=  8'h00;      memory[58775] <=  8'h00;      memory[58776] <=  8'h00;      memory[58777] <=  8'h00;      memory[58778] <=  8'h00;      memory[58779] <=  8'h00;      memory[58780] <=  8'h00;      memory[58781] <=  8'h00;      memory[58782] <=  8'h00;      memory[58783] <=  8'h00;      memory[58784] <=  8'h00;      memory[58785] <=  8'h00;      memory[58786] <=  8'h00;      memory[58787] <=  8'h00;      memory[58788] <=  8'h00;      memory[58789] <=  8'h00;      memory[58790] <=  8'h00;      memory[58791] <=  8'h00;      memory[58792] <=  8'h00;      memory[58793] <=  8'h00;      memory[58794] <=  8'h00;      memory[58795] <=  8'h00;      memory[58796] <=  8'h00;      memory[58797] <=  8'h00;      memory[58798] <=  8'h00;      memory[58799] <=  8'h00;      memory[58800] <=  8'h00;      memory[58801] <=  8'h00;      memory[58802] <=  8'h00;      memory[58803] <=  8'h00;      memory[58804] <=  8'h00;      memory[58805] <=  8'h00;      memory[58806] <=  8'h00;      memory[58807] <=  8'h00;      memory[58808] <=  8'h00;      memory[58809] <=  8'h00;      memory[58810] <=  8'h00;      memory[58811] <=  8'h00;      memory[58812] <=  8'h00;      memory[58813] <=  8'h00;      memory[58814] <=  8'h00;      memory[58815] <=  8'h00;      memory[58816] <=  8'h00;      memory[58817] <=  8'h00;      memory[58818] <=  8'h00;      memory[58819] <=  8'h00;      memory[58820] <=  8'h00;      memory[58821] <=  8'h00;      memory[58822] <=  8'h00;      memory[58823] <=  8'h00;      memory[58824] <=  8'h00;      memory[58825] <=  8'h00;      memory[58826] <=  8'h00;      memory[58827] <=  8'h00;      memory[58828] <=  8'h00;      memory[58829] <=  8'h00;      memory[58830] <=  8'h00;      memory[58831] <=  8'h00;      memory[58832] <=  8'h00;      memory[58833] <=  8'h00;      memory[58834] <=  8'h00;      memory[58835] <=  8'h00;      memory[58836] <=  8'h00;      memory[58837] <=  8'h00;      memory[58838] <=  8'h00;      memory[58839] <=  8'h00;      memory[58840] <=  8'h00;      memory[58841] <=  8'h00;      memory[58842] <=  8'h00;      memory[58843] <=  8'h00;      memory[58844] <=  8'h00;      memory[58845] <=  8'h00;      memory[58846] <=  8'h00;      memory[58847] <=  8'h00;      memory[58848] <=  8'h00;      memory[58849] <=  8'h00;      memory[58850] <=  8'h00;      memory[58851] <=  8'h00;      memory[58852] <=  8'h00;      memory[58853] <=  8'h00;      memory[58854] <=  8'h00;      memory[58855] <=  8'h00;      memory[58856] <=  8'h00;      memory[58857] <=  8'h00;      memory[58858] <=  8'h00;      memory[58859] <=  8'h00;      memory[58860] <=  8'h00;      memory[58861] <=  8'h00;      memory[58862] <=  8'h00;      memory[58863] <=  8'h00;      memory[58864] <=  8'h00;      memory[58865] <=  8'h00;      memory[58866] <=  8'h00;      memory[58867] <=  8'h00;      memory[58868] <=  8'h00;      memory[58869] <=  8'h00;      memory[58870] <=  8'h00;      memory[58871] <=  8'h00;      memory[58872] <=  8'h00;      memory[58873] <=  8'h00;      memory[58874] <=  8'h00;      memory[58875] <=  8'h00;      memory[58876] <=  8'h00;      memory[58877] <=  8'h00;      memory[58878] <=  8'h00;      memory[58879] <=  8'h00;      memory[58880] <=  8'h00;      memory[58881] <=  8'h00;      memory[58882] <=  8'h00;      memory[58883] <=  8'h00;      memory[58884] <=  8'h00;      memory[58885] <=  8'h00;      memory[58886] <=  8'h00;      memory[58887] <=  8'h00;      memory[58888] <=  8'h00;      memory[58889] <=  8'h00;      memory[58890] <=  8'h00;      memory[58891] <=  8'h00;      memory[58892] <=  8'h00;      memory[58893] <=  8'h00;      memory[58894] <=  8'h00;      memory[58895] <=  8'h00;      memory[58896] <=  8'h00;      memory[58897] <=  8'h00;      memory[58898] <=  8'h00;      memory[58899] <=  8'h00;      memory[58900] <=  8'h00;      memory[58901] <=  8'h00;      memory[58902] <=  8'h00;      memory[58903] <=  8'h00;      memory[58904] <=  8'h00;      memory[58905] <=  8'h00;      memory[58906] <=  8'h00;      memory[58907] <=  8'h00;      memory[58908] <=  8'h00;      memory[58909] <=  8'h00;      memory[58910] <=  8'h00;      memory[58911] <=  8'h00;      memory[58912] <=  8'h00;      memory[58913] <=  8'h00;      memory[58914] <=  8'h00;      memory[58915] <=  8'h00;      memory[58916] <=  8'h00;      memory[58917] <=  8'h00;      memory[58918] <=  8'h00;      memory[58919] <=  8'h00;      memory[58920] <=  8'h00;      memory[58921] <=  8'h00;      memory[58922] <=  8'h00;      memory[58923] <=  8'h00;      memory[58924] <=  8'h00;      memory[58925] <=  8'h00;      memory[58926] <=  8'h00;      memory[58927] <=  8'h00;      memory[58928] <=  8'h00;      memory[58929] <=  8'h00;      memory[58930] <=  8'h00;      memory[58931] <=  8'h00;      memory[58932] <=  8'h00;      memory[58933] <=  8'h00;      memory[58934] <=  8'h00;      memory[58935] <=  8'h00;      memory[58936] <=  8'h00;      memory[58937] <=  8'h00;      memory[58938] <=  8'h00;      memory[58939] <=  8'h00;      memory[58940] <=  8'h00;      memory[58941] <=  8'h00;      memory[58942] <=  8'h00;      memory[58943] <=  8'h00;      memory[58944] <=  8'h00;      memory[58945] <=  8'h00;      memory[58946] <=  8'h00;      memory[58947] <=  8'h00;      memory[58948] <=  8'h00;      memory[58949] <=  8'h00;      memory[58950] <=  8'h00;      memory[58951] <=  8'h00;      memory[58952] <=  8'h00;      memory[58953] <=  8'h00;      memory[58954] <=  8'h00;      memory[58955] <=  8'h00;      memory[58956] <=  8'h00;      memory[58957] <=  8'h00;      memory[58958] <=  8'h00;      memory[58959] <=  8'h00;      memory[58960] <=  8'h00;      memory[58961] <=  8'h00;      memory[58962] <=  8'h00;      memory[58963] <=  8'h00;      memory[58964] <=  8'h00;      memory[58965] <=  8'h00;      memory[58966] <=  8'h00;      memory[58967] <=  8'h00;      memory[58968] <=  8'h00;      memory[58969] <=  8'h00;      memory[58970] <=  8'h00;      memory[58971] <=  8'h00;      memory[58972] <=  8'h00;      memory[58973] <=  8'h00;      memory[58974] <=  8'h00;      memory[58975] <=  8'h00;      memory[58976] <=  8'h00;      memory[58977] <=  8'h00;      memory[58978] <=  8'h00;      memory[58979] <=  8'h00;      memory[58980] <=  8'h00;      memory[58981] <=  8'h00;      memory[58982] <=  8'h00;      memory[58983] <=  8'h00;      memory[58984] <=  8'h00;      memory[58985] <=  8'h00;      memory[58986] <=  8'h00;      memory[58987] <=  8'h00;      memory[58988] <=  8'h00;      memory[58989] <=  8'h00;      memory[58990] <=  8'h00;      memory[58991] <=  8'h00;      memory[58992] <=  8'h00;      memory[58993] <=  8'h00;      memory[58994] <=  8'h00;      memory[58995] <=  8'h00;      memory[58996] <=  8'h00;      memory[58997] <=  8'h00;      memory[58998] <=  8'h00;      memory[58999] <=  8'h00;      memory[59000] <=  8'h00;      memory[59001] <=  8'h00;      memory[59002] <=  8'h00;      memory[59003] <=  8'h00;      memory[59004] <=  8'h00;      memory[59005] <=  8'h00;      memory[59006] <=  8'h00;      memory[59007] <=  8'h00;      memory[59008] <=  8'h00;      memory[59009] <=  8'h00;      memory[59010] <=  8'h00;      memory[59011] <=  8'h00;      memory[59012] <=  8'h00;      memory[59013] <=  8'h00;      memory[59014] <=  8'h00;      memory[59015] <=  8'h00;      memory[59016] <=  8'h00;      memory[59017] <=  8'h00;      memory[59018] <=  8'h00;      memory[59019] <=  8'h00;      memory[59020] <=  8'h00;      memory[59021] <=  8'h00;      memory[59022] <=  8'h00;      memory[59023] <=  8'h00;      memory[59024] <=  8'h00;      memory[59025] <=  8'h00;      memory[59026] <=  8'h00;      memory[59027] <=  8'h00;      memory[59028] <=  8'h00;      memory[59029] <=  8'h00;      memory[59030] <=  8'h00;      memory[59031] <=  8'h00;      memory[59032] <=  8'h00;      memory[59033] <=  8'h00;      memory[59034] <=  8'h00;      memory[59035] <=  8'h00;      memory[59036] <=  8'h00;      memory[59037] <=  8'h00;      memory[59038] <=  8'h00;      memory[59039] <=  8'h00;      memory[59040] <=  8'h00;      memory[59041] <=  8'h00;      memory[59042] <=  8'h00;      memory[59043] <=  8'h00;      memory[59044] <=  8'h00;      memory[59045] <=  8'h00;      memory[59046] <=  8'h00;      memory[59047] <=  8'h00;      memory[59048] <=  8'h00;      memory[59049] <=  8'h00;      memory[59050] <=  8'h00;      memory[59051] <=  8'h00;      memory[59052] <=  8'h00;      memory[59053] <=  8'h00;      memory[59054] <=  8'h00;      memory[59055] <=  8'h00;      memory[59056] <=  8'h00;      memory[59057] <=  8'h00;      memory[59058] <=  8'h00;      memory[59059] <=  8'h00;      memory[59060] <=  8'h00;      memory[59061] <=  8'h00;      memory[59062] <=  8'h00;      memory[59063] <=  8'h00;      memory[59064] <=  8'h00;      memory[59065] <=  8'h00;      memory[59066] <=  8'h00;      memory[59067] <=  8'h00;      memory[59068] <=  8'h00;      memory[59069] <=  8'h00;      memory[59070] <=  8'h00;      memory[59071] <=  8'h00;      memory[59072] <=  8'h00;      memory[59073] <=  8'h00;      memory[59074] <=  8'h00;      memory[59075] <=  8'h00;      memory[59076] <=  8'h00;      memory[59077] <=  8'h00;      memory[59078] <=  8'h00;      memory[59079] <=  8'h00;      memory[59080] <=  8'h00;      memory[59081] <=  8'h00;      memory[59082] <=  8'h00;      memory[59083] <=  8'h00;      memory[59084] <=  8'h00;      memory[59085] <=  8'h00;      memory[59086] <=  8'h00;      memory[59087] <=  8'h00;      memory[59088] <=  8'h00;      memory[59089] <=  8'h00;      memory[59090] <=  8'h00;      memory[59091] <=  8'h00;      memory[59092] <=  8'h00;      memory[59093] <=  8'h00;      memory[59094] <=  8'h00;      memory[59095] <=  8'h00;      memory[59096] <=  8'h00;      memory[59097] <=  8'h00;      memory[59098] <=  8'h00;      memory[59099] <=  8'h00;      memory[59100] <=  8'h00;      memory[59101] <=  8'h00;      memory[59102] <=  8'h00;      memory[59103] <=  8'h00;      memory[59104] <=  8'h00;      memory[59105] <=  8'h00;      memory[59106] <=  8'h00;      memory[59107] <=  8'h00;      memory[59108] <=  8'h00;      memory[59109] <=  8'h00;      memory[59110] <=  8'h00;      memory[59111] <=  8'h00;      memory[59112] <=  8'h00;      memory[59113] <=  8'h00;      memory[59114] <=  8'h00;      memory[59115] <=  8'h00;      memory[59116] <=  8'h00;      memory[59117] <=  8'h00;      memory[59118] <=  8'h00;      memory[59119] <=  8'h00;      memory[59120] <=  8'h00;      memory[59121] <=  8'h00;      memory[59122] <=  8'h00;      memory[59123] <=  8'h00;      memory[59124] <=  8'h00;      memory[59125] <=  8'h00;      memory[59126] <=  8'h00;      memory[59127] <=  8'h00;      memory[59128] <=  8'h00;      memory[59129] <=  8'h00;      memory[59130] <=  8'h00;      memory[59131] <=  8'h00;      memory[59132] <=  8'h00;      memory[59133] <=  8'h00;      memory[59134] <=  8'h00;      memory[59135] <=  8'h00;      memory[59136] <=  8'h00;      memory[59137] <=  8'h00;      memory[59138] <=  8'h00;      memory[59139] <=  8'h00;      memory[59140] <=  8'h00;      memory[59141] <=  8'h00;      memory[59142] <=  8'h00;      memory[59143] <=  8'h00;      memory[59144] <=  8'h00;      memory[59145] <=  8'h00;      memory[59146] <=  8'h00;      memory[59147] <=  8'h00;      memory[59148] <=  8'h00;      memory[59149] <=  8'h00;      memory[59150] <=  8'h00;      memory[59151] <=  8'h00;      memory[59152] <=  8'h00;      memory[59153] <=  8'h00;      memory[59154] <=  8'h00;      memory[59155] <=  8'h00;      memory[59156] <=  8'h00;      memory[59157] <=  8'h00;      memory[59158] <=  8'h00;      memory[59159] <=  8'h00;      memory[59160] <=  8'h00;      memory[59161] <=  8'h00;      memory[59162] <=  8'h00;      memory[59163] <=  8'h00;      memory[59164] <=  8'h00;      memory[59165] <=  8'h00;      memory[59166] <=  8'h00;      memory[59167] <=  8'h00;      memory[59168] <=  8'h00;      memory[59169] <=  8'h00;      memory[59170] <=  8'h00;      memory[59171] <=  8'h00;      memory[59172] <=  8'h00;      memory[59173] <=  8'h00;      memory[59174] <=  8'h00;      memory[59175] <=  8'h00;      memory[59176] <=  8'h00;      memory[59177] <=  8'h00;      memory[59178] <=  8'h00;      memory[59179] <=  8'h00;      memory[59180] <=  8'h00;      memory[59181] <=  8'h00;      memory[59182] <=  8'h00;      memory[59183] <=  8'h00;      memory[59184] <=  8'h00;      memory[59185] <=  8'h00;      memory[59186] <=  8'h00;      memory[59187] <=  8'h00;      memory[59188] <=  8'h00;      memory[59189] <=  8'h00;      memory[59190] <=  8'h00;      memory[59191] <=  8'h00;      memory[59192] <=  8'h00;      memory[59193] <=  8'h00;      memory[59194] <=  8'h00;      memory[59195] <=  8'h00;      memory[59196] <=  8'h00;      memory[59197] <=  8'h00;      memory[59198] <=  8'h00;      memory[59199] <=  8'h00;      memory[59200] <=  8'h00;      memory[59201] <=  8'h00;      memory[59202] <=  8'h00;      memory[59203] <=  8'h00;      memory[59204] <=  8'h00;      memory[59205] <=  8'h00;      memory[59206] <=  8'h00;      memory[59207] <=  8'h00;      memory[59208] <=  8'h00;      memory[59209] <=  8'h00;      memory[59210] <=  8'h00;      memory[59211] <=  8'h00;      memory[59212] <=  8'h00;      memory[59213] <=  8'h00;      memory[59214] <=  8'h00;      memory[59215] <=  8'h00;      memory[59216] <=  8'h00;      memory[59217] <=  8'h00;      memory[59218] <=  8'h00;      memory[59219] <=  8'h00;      memory[59220] <=  8'h00;      memory[59221] <=  8'h00;      memory[59222] <=  8'h00;      memory[59223] <=  8'h00;      memory[59224] <=  8'h00;      memory[59225] <=  8'h00;      memory[59226] <=  8'h00;      memory[59227] <=  8'h00;      memory[59228] <=  8'h00;      memory[59229] <=  8'h00;      memory[59230] <=  8'h00;      memory[59231] <=  8'h00;      memory[59232] <=  8'h00;      memory[59233] <=  8'h00;      memory[59234] <=  8'h00;      memory[59235] <=  8'h00;      memory[59236] <=  8'h00;      memory[59237] <=  8'h00;      memory[59238] <=  8'h00;      memory[59239] <=  8'h00;      memory[59240] <=  8'h00;      memory[59241] <=  8'h00;      memory[59242] <=  8'h00;      memory[59243] <=  8'h00;      memory[59244] <=  8'h00;      memory[59245] <=  8'h00;      memory[59246] <=  8'h00;      memory[59247] <=  8'h00;      memory[59248] <=  8'h00;      memory[59249] <=  8'h00;      memory[59250] <=  8'h00;      memory[59251] <=  8'h00;      memory[59252] <=  8'h00;      memory[59253] <=  8'h00;      memory[59254] <=  8'h00;      memory[59255] <=  8'h00;      memory[59256] <=  8'h00;      memory[59257] <=  8'h00;      memory[59258] <=  8'h00;      memory[59259] <=  8'h00;      memory[59260] <=  8'h00;      memory[59261] <=  8'h00;      memory[59262] <=  8'h00;      memory[59263] <=  8'h00;      memory[59264] <=  8'h00;      memory[59265] <=  8'h00;      memory[59266] <=  8'h00;      memory[59267] <=  8'h00;      memory[59268] <=  8'h00;      memory[59269] <=  8'h00;      memory[59270] <=  8'h00;      memory[59271] <=  8'h00;      memory[59272] <=  8'h00;      memory[59273] <=  8'h00;      memory[59274] <=  8'h00;      memory[59275] <=  8'h00;      memory[59276] <=  8'h00;      memory[59277] <=  8'h00;      memory[59278] <=  8'h00;      memory[59279] <=  8'h00;      memory[59280] <=  8'h00;      memory[59281] <=  8'h00;      memory[59282] <=  8'h00;      memory[59283] <=  8'h00;      memory[59284] <=  8'h00;      memory[59285] <=  8'h00;      memory[59286] <=  8'h00;      memory[59287] <=  8'h00;      memory[59288] <=  8'h00;      memory[59289] <=  8'h00;      memory[59290] <=  8'h00;      memory[59291] <=  8'h00;      memory[59292] <=  8'h00;      memory[59293] <=  8'h00;      memory[59294] <=  8'h00;      memory[59295] <=  8'h00;      memory[59296] <=  8'h00;      memory[59297] <=  8'h00;      memory[59298] <=  8'h00;      memory[59299] <=  8'h00;      memory[59300] <=  8'h00;      memory[59301] <=  8'h00;      memory[59302] <=  8'h00;      memory[59303] <=  8'h00;      memory[59304] <=  8'h00;      memory[59305] <=  8'h00;      memory[59306] <=  8'h00;      memory[59307] <=  8'h00;      memory[59308] <=  8'h00;      memory[59309] <=  8'h00;      memory[59310] <=  8'h00;      memory[59311] <=  8'h00;      memory[59312] <=  8'h00;      memory[59313] <=  8'h00;      memory[59314] <=  8'h00;      memory[59315] <=  8'h00;      memory[59316] <=  8'h00;      memory[59317] <=  8'h00;      memory[59318] <=  8'h00;      memory[59319] <=  8'h00;      memory[59320] <=  8'h00;      memory[59321] <=  8'h00;      memory[59322] <=  8'h00;      memory[59323] <=  8'h00;      memory[59324] <=  8'h00;      memory[59325] <=  8'h00;      memory[59326] <=  8'h00;      memory[59327] <=  8'h00;      memory[59328] <=  8'h00;      memory[59329] <=  8'h00;      memory[59330] <=  8'h00;      memory[59331] <=  8'h00;      memory[59332] <=  8'h00;      memory[59333] <=  8'h00;      memory[59334] <=  8'h00;      memory[59335] <=  8'h00;      memory[59336] <=  8'h00;      memory[59337] <=  8'h00;      memory[59338] <=  8'h00;      memory[59339] <=  8'h00;      memory[59340] <=  8'h00;      memory[59341] <=  8'h00;      memory[59342] <=  8'h00;      memory[59343] <=  8'h00;      memory[59344] <=  8'h00;      memory[59345] <=  8'h00;      memory[59346] <=  8'h00;      memory[59347] <=  8'h00;      memory[59348] <=  8'h00;      memory[59349] <=  8'h00;      memory[59350] <=  8'h00;      memory[59351] <=  8'h00;      memory[59352] <=  8'h00;      memory[59353] <=  8'h00;      memory[59354] <=  8'h00;      memory[59355] <=  8'h00;      memory[59356] <=  8'h00;      memory[59357] <=  8'h00;      memory[59358] <=  8'h00;      memory[59359] <=  8'h00;      memory[59360] <=  8'h00;      memory[59361] <=  8'h00;      memory[59362] <=  8'h00;      memory[59363] <=  8'h00;      memory[59364] <=  8'h00;      memory[59365] <=  8'h00;      memory[59366] <=  8'h00;      memory[59367] <=  8'h00;      memory[59368] <=  8'h00;      memory[59369] <=  8'h00;      memory[59370] <=  8'h00;      memory[59371] <=  8'h00;      memory[59372] <=  8'h00;      memory[59373] <=  8'h00;      memory[59374] <=  8'h00;      memory[59375] <=  8'h00;      memory[59376] <=  8'h00;      memory[59377] <=  8'h00;      memory[59378] <=  8'h00;      memory[59379] <=  8'h00;      memory[59380] <=  8'h00;      memory[59381] <=  8'h00;      memory[59382] <=  8'h00;      memory[59383] <=  8'h00;      memory[59384] <=  8'h00;      memory[59385] <=  8'h00;      memory[59386] <=  8'h00;      memory[59387] <=  8'h00;      memory[59388] <=  8'h00;      memory[59389] <=  8'h00;      memory[59390] <=  8'h00;      memory[59391] <=  8'h00;      memory[59392] <=  8'h00;      memory[59393] <=  8'h00;      memory[59394] <=  8'h00;      memory[59395] <=  8'h00;      memory[59396] <=  8'h00;      memory[59397] <=  8'h00;      memory[59398] <=  8'h00;      memory[59399] <=  8'h00;      memory[59400] <=  8'h00;      memory[59401] <=  8'h00;      memory[59402] <=  8'h00;      memory[59403] <=  8'h00;      memory[59404] <=  8'h00;      memory[59405] <=  8'h00;      memory[59406] <=  8'h00;      memory[59407] <=  8'h00;      memory[59408] <=  8'h00;      memory[59409] <=  8'h00;      memory[59410] <=  8'h00;      memory[59411] <=  8'h00;      memory[59412] <=  8'h00;      memory[59413] <=  8'h00;      memory[59414] <=  8'h00;      memory[59415] <=  8'h00;      memory[59416] <=  8'h00;      memory[59417] <=  8'h00;      memory[59418] <=  8'h00;      memory[59419] <=  8'h00;      memory[59420] <=  8'h00;      memory[59421] <=  8'h00;      memory[59422] <=  8'h00;      memory[59423] <=  8'h00;      memory[59424] <=  8'h00;      memory[59425] <=  8'h00;      memory[59426] <=  8'h00;      memory[59427] <=  8'h00;      memory[59428] <=  8'h00;      memory[59429] <=  8'h00;      memory[59430] <=  8'h00;      memory[59431] <=  8'h00;      memory[59432] <=  8'h00;      memory[59433] <=  8'h00;      memory[59434] <=  8'h00;      memory[59435] <=  8'h00;      memory[59436] <=  8'h00;      memory[59437] <=  8'h00;      memory[59438] <=  8'h00;      memory[59439] <=  8'h00;      memory[59440] <=  8'h00;      memory[59441] <=  8'h00;      memory[59442] <=  8'h00;      memory[59443] <=  8'h00;      memory[59444] <=  8'h00;      memory[59445] <=  8'h00;      memory[59446] <=  8'h00;      memory[59447] <=  8'h00;      memory[59448] <=  8'h00;      memory[59449] <=  8'h00;      memory[59450] <=  8'h00;      memory[59451] <=  8'h00;      memory[59452] <=  8'h00;      memory[59453] <=  8'h00;      memory[59454] <=  8'h00;      memory[59455] <=  8'h00;      memory[59456] <=  8'h00;      memory[59457] <=  8'h00;      memory[59458] <=  8'h00;      memory[59459] <=  8'h00;      memory[59460] <=  8'h00;      memory[59461] <=  8'h00;      memory[59462] <=  8'h00;      memory[59463] <=  8'h00;      memory[59464] <=  8'h00;      memory[59465] <=  8'h00;      memory[59466] <=  8'h00;      memory[59467] <=  8'h00;      memory[59468] <=  8'h00;      memory[59469] <=  8'h00;      memory[59470] <=  8'h00;      memory[59471] <=  8'h00;      memory[59472] <=  8'h00;      memory[59473] <=  8'h00;      memory[59474] <=  8'h00;      memory[59475] <=  8'h00;      memory[59476] <=  8'h00;      memory[59477] <=  8'h00;      memory[59478] <=  8'h00;      memory[59479] <=  8'h00;      memory[59480] <=  8'h00;      memory[59481] <=  8'h00;      memory[59482] <=  8'h00;      memory[59483] <=  8'h00;      memory[59484] <=  8'h00;      memory[59485] <=  8'h00;      memory[59486] <=  8'h00;      memory[59487] <=  8'h00;      memory[59488] <=  8'h00;      memory[59489] <=  8'h00;      memory[59490] <=  8'h00;      memory[59491] <=  8'h00;      memory[59492] <=  8'h00;      memory[59493] <=  8'h00;      memory[59494] <=  8'h00;      memory[59495] <=  8'h00;      memory[59496] <=  8'h00;      memory[59497] <=  8'h00;      memory[59498] <=  8'h00;      memory[59499] <=  8'h00;      memory[59500] <=  8'h00;      memory[59501] <=  8'h00;      memory[59502] <=  8'h00;      memory[59503] <=  8'h00;      memory[59504] <=  8'h00;      memory[59505] <=  8'h00;      memory[59506] <=  8'h00;      memory[59507] <=  8'h00;      memory[59508] <=  8'h00;      memory[59509] <=  8'h00;      memory[59510] <=  8'h00;      memory[59511] <=  8'h00;      memory[59512] <=  8'h00;      memory[59513] <=  8'h00;      memory[59514] <=  8'h00;      memory[59515] <=  8'h00;      memory[59516] <=  8'h00;      memory[59517] <=  8'h00;      memory[59518] <=  8'h00;      memory[59519] <=  8'h00;      memory[59520] <=  8'h00;      memory[59521] <=  8'h00;      memory[59522] <=  8'h00;      memory[59523] <=  8'h00;      memory[59524] <=  8'h00;      memory[59525] <=  8'h00;      memory[59526] <=  8'h00;      memory[59527] <=  8'h00;      memory[59528] <=  8'h00;      memory[59529] <=  8'h00;      memory[59530] <=  8'h00;      memory[59531] <=  8'h00;      memory[59532] <=  8'h00;      memory[59533] <=  8'h00;      memory[59534] <=  8'h00;      memory[59535] <=  8'h00;      memory[59536] <=  8'h00;      memory[59537] <=  8'h00;      memory[59538] <=  8'h00;      memory[59539] <=  8'h00;      memory[59540] <=  8'h00;      memory[59541] <=  8'h00;      memory[59542] <=  8'h00;      memory[59543] <=  8'h00;      memory[59544] <=  8'h00;      memory[59545] <=  8'h00;      memory[59546] <=  8'h00;      memory[59547] <=  8'h00;      memory[59548] <=  8'h00;      memory[59549] <=  8'h00;      memory[59550] <=  8'h00;      memory[59551] <=  8'h00;      memory[59552] <=  8'h00;      memory[59553] <=  8'h00;      memory[59554] <=  8'h00;      memory[59555] <=  8'h00;      memory[59556] <=  8'h00;      memory[59557] <=  8'h00;      memory[59558] <=  8'h00;      memory[59559] <=  8'h00;      memory[59560] <=  8'h00;      memory[59561] <=  8'h00;      memory[59562] <=  8'h00;      memory[59563] <=  8'h00;      memory[59564] <=  8'h00;      memory[59565] <=  8'h00;      memory[59566] <=  8'h00;      memory[59567] <=  8'h00;      memory[59568] <=  8'h00;      memory[59569] <=  8'h00;      memory[59570] <=  8'h00;      memory[59571] <=  8'h00;      memory[59572] <=  8'h00;      memory[59573] <=  8'h00;      memory[59574] <=  8'h00;      memory[59575] <=  8'h00;      memory[59576] <=  8'h00;      memory[59577] <=  8'h00;      memory[59578] <=  8'h00;      memory[59579] <=  8'h00;      memory[59580] <=  8'h00;      memory[59581] <=  8'h00;      memory[59582] <=  8'h00;      memory[59583] <=  8'h00;      memory[59584] <=  8'h00;      memory[59585] <=  8'h00;      memory[59586] <=  8'h00;      memory[59587] <=  8'h00;      memory[59588] <=  8'h00;      memory[59589] <=  8'h00;      memory[59590] <=  8'h00;      memory[59591] <=  8'h00;      memory[59592] <=  8'h00;      memory[59593] <=  8'h00;      memory[59594] <=  8'h00;      memory[59595] <=  8'h00;      memory[59596] <=  8'h00;      memory[59597] <=  8'h00;      memory[59598] <=  8'h00;      memory[59599] <=  8'h00;      memory[59600] <=  8'h00;      memory[59601] <=  8'h00;      memory[59602] <=  8'h00;      memory[59603] <=  8'h00;      memory[59604] <=  8'h00;      memory[59605] <=  8'h00;      memory[59606] <=  8'h00;      memory[59607] <=  8'h00;      memory[59608] <=  8'h00;      memory[59609] <=  8'h00;      memory[59610] <=  8'h00;      memory[59611] <=  8'h00;      memory[59612] <=  8'h00;      memory[59613] <=  8'h00;      memory[59614] <=  8'h00;      memory[59615] <=  8'h00;      memory[59616] <=  8'h00;      memory[59617] <=  8'h00;      memory[59618] <=  8'h00;      memory[59619] <=  8'h00;      memory[59620] <=  8'h00;      memory[59621] <=  8'h00;      memory[59622] <=  8'h00;      memory[59623] <=  8'h00;      memory[59624] <=  8'h00;      memory[59625] <=  8'h00;      memory[59626] <=  8'h00;      memory[59627] <=  8'h00;      memory[59628] <=  8'h00;      memory[59629] <=  8'h00;      memory[59630] <=  8'h00;      memory[59631] <=  8'h00;      memory[59632] <=  8'h00;      memory[59633] <=  8'h00;      memory[59634] <=  8'h00;      memory[59635] <=  8'h00;      memory[59636] <=  8'h00;      memory[59637] <=  8'h00;      memory[59638] <=  8'h00;      memory[59639] <=  8'h00;      memory[59640] <=  8'h00;      memory[59641] <=  8'h00;      memory[59642] <=  8'h00;      memory[59643] <=  8'h00;      memory[59644] <=  8'h00;      memory[59645] <=  8'h00;      memory[59646] <=  8'h00;      memory[59647] <=  8'h00;      memory[59648] <=  8'h00;      memory[59649] <=  8'h00;      memory[59650] <=  8'h00;      memory[59651] <=  8'h00;      memory[59652] <=  8'h00;      memory[59653] <=  8'h00;      memory[59654] <=  8'h00;      memory[59655] <=  8'h00;      memory[59656] <=  8'h00;      memory[59657] <=  8'h00;      memory[59658] <=  8'h00;      memory[59659] <=  8'h00;      memory[59660] <=  8'h00;      memory[59661] <=  8'h00;      memory[59662] <=  8'h00;      memory[59663] <=  8'h00;      memory[59664] <=  8'h00;      memory[59665] <=  8'h00;      memory[59666] <=  8'h00;      memory[59667] <=  8'h00;      memory[59668] <=  8'h00;      memory[59669] <=  8'h00;      memory[59670] <=  8'h00;      memory[59671] <=  8'h00;      memory[59672] <=  8'h00;      memory[59673] <=  8'h00;      memory[59674] <=  8'h00;      memory[59675] <=  8'h00;      memory[59676] <=  8'h00;      memory[59677] <=  8'h00;      memory[59678] <=  8'h00;      memory[59679] <=  8'h00;      memory[59680] <=  8'h00;      memory[59681] <=  8'h00;      memory[59682] <=  8'h00;      memory[59683] <=  8'h00;      memory[59684] <=  8'h00;      memory[59685] <=  8'h00;      memory[59686] <=  8'h00;      memory[59687] <=  8'h00;      memory[59688] <=  8'h00;      memory[59689] <=  8'h00;      memory[59690] <=  8'h00;      memory[59691] <=  8'h00;      memory[59692] <=  8'h00;      memory[59693] <=  8'h00;      memory[59694] <=  8'h00;      memory[59695] <=  8'h00;      memory[59696] <=  8'h00;      memory[59697] <=  8'h00;      memory[59698] <=  8'h00;      memory[59699] <=  8'h00;      memory[59700] <=  8'h00;      memory[59701] <=  8'h00;      memory[59702] <=  8'h00;      memory[59703] <=  8'h00;      memory[59704] <=  8'h00;      memory[59705] <=  8'h00;      memory[59706] <=  8'h00;      memory[59707] <=  8'h00;      memory[59708] <=  8'h00;      memory[59709] <=  8'h00;      memory[59710] <=  8'h00;      memory[59711] <=  8'h00;      memory[59712] <=  8'h00;      memory[59713] <=  8'h00;      memory[59714] <=  8'h00;      memory[59715] <=  8'h00;      memory[59716] <=  8'h00;      memory[59717] <=  8'h00;      memory[59718] <=  8'h00;      memory[59719] <=  8'h00;      memory[59720] <=  8'h00;      memory[59721] <=  8'h00;      memory[59722] <=  8'h00;      memory[59723] <=  8'h00;      memory[59724] <=  8'h00;      memory[59725] <=  8'h00;      memory[59726] <=  8'h00;      memory[59727] <=  8'h00;      memory[59728] <=  8'h00;      memory[59729] <=  8'h00;      memory[59730] <=  8'h00;      memory[59731] <=  8'h00;      memory[59732] <=  8'h00;      memory[59733] <=  8'h00;      memory[59734] <=  8'h00;      memory[59735] <=  8'h00;      memory[59736] <=  8'h00;      memory[59737] <=  8'h00;      memory[59738] <=  8'h00;      memory[59739] <=  8'h00;      memory[59740] <=  8'h00;      memory[59741] <=  8'h00;      memory[59742] <=  8'h00;      memory[59743] <=  8'h00;      memory[59744] <=  8'h00;      memory[59745] <=  8'h00;      memory[59746] <=  8'h00;      memory[59747] <=  8'h00;      memory[59748] <=  8'h00;      memory[59749] <=  8'h00;      memory[59750] <=  8'h00;      memory[59751] <=  8'h00;      memory[59752] <=  8'h00;      memory[59753] <=  8'h00;      memory[59754] <=  8'h00;      memory[59755] <=  8'h00;      memory[59756] <=  8'h00;      memory[59757] <=  8'h00;      memory[59758] <=  8'h00;      memory[59759] <=  8'h00;      memory[59760] <=  8'h00;      memory[59761] <=  8'h00;      memory[59762] <=  8'h00;      memory[59763] <=  8'h00;      memory[59764] <=  8'h00;      memory[59765] <=  8'h00;      memory[59766] <=  8'h00;      memory[59767] <=  8'h00;      memory[59768] <=  8'h00;      memory[59769] <=  8'h00;      memory[59770] <=  8'h00;      memory[59771] <=  8'h00;      memory[59772] <=  8'h00;      memory[59773] <=  8'h00;      memory[59774] <=  8'h00;      memory[59775] <=  8'h00;      memory[59776] <=  8'h00;      memory[59777] <=  8'h00;      memory[59778] <=  8'h00;      memory[59779] <=  8'h00;      memory[59780] <=  8'h00;      memory[59781] <=  8'h00;      memory[59782] <=  8'h00;      memory[59783] <=  8'h00;      memory[59784] <=  8'h00;      memory[59785] <=  8'h00;      memory[59786] <=  8'h00;      memory[59787] <=  8'h00;      memory[59788] <=  8'h00;      memory[59789] <=  8'h00;      memory[59790] <=  8'h00;      memory[59791] <=  8'h00;      memory[59792] <=  8'h00;      memory[59793] <=  8'h00;      memory[59794] <=  8'h00;      memory[59795] <=  8'h00;      memory[59796] <=  8'h00;      memory[59797] <=  8'h00;      memory[59798] <=  8'h00;      memory[59799] <=  8'h00;      memory[59800] <=  8'h00;      memory[59801] <=  8'h00;      memory[59802] <=  8'h00;      memory[59803] <=  8'h00;      memory[59804] <=  8'h00;      memory[59805] <=  8'h00;      memory[59806] <=  8'h00;      memory[59807] <=  8'h00;      memory[59808] <=  8'h00;      memory[59809] <=  8'h00;      memory[59810] <=  8'h00;      memory[59811] <=  8'h00;      memory[59812] <=  8'h00;      memory[59813] <=  8'h00;      memory[59814] <=  8'h00;      memory[59815] <=  8'h00;      memory[59816] <=  8'h00;      memory[59817] <=  8'h00;      memory[59818] <=  8'h00;      memory[59819] <=  8'h00;      memory[59820] <=  8'h00;      memory[59821] <=  8'h00;      memory[59822] <=  8'h00;      memory[59823] <=  8'h00;      memory[59824] <=  8'h00;      memory[59825] <=  8'h00;      memory[59826] <=  8'h00;      memory[59827] <=  8'h00;      memory[59828] <=  8'h00;      memory[59829] <=  8'h00;      memory[59830] <=  8'h00;      memory[59831] <=  8'h00;      memory[59832] <=  8'h00;      memory[59833] <=  8'h00;      memory[59834] <=  8'h00;      memory[59835] <=  8'h00;      memory[59836] <=  8'h00;      memory[59837] <=  8'h00;      memory[59838] <=  8'h00;      memory[59839] <=  8'h00;      memory[59840] <=  8'h00;      memory[59841] <=  8'h00;      memory[59842] <=  8'h00;      memory[59843] <=  8'h00;      memory[59844] <=  8'h00;      memory[59845] <=  8'h00;      memory[59846] <=  8'h00;      memory[59847] <=  8'h00;      memory[59848] <=  8'h00;      memory[59849] <=  8'h00;      memory[59850] <=  8'h00;      memory[59851] <=  8'h00;      memory[59852] <=  8'h00;      memory[59853] <=  8'h00;      memory[59854] <=  8'h00;      memory[59855] <=  8'h00;      memory[59856] <=  8'h00;      memory[59857] <=  8'h00;      memory[59858] <=  8'h00;      memory[59859] <=  8'h00;      memory[59860] <=  8'h00;      memory[59861] <=  8'h00;      memory[59862] <=  8'h00;      memory[59863] <=  8'h00;      memory[59864] <=  8'h00;      memory[59865] <=  8'h00;      memory[59866] <=  8'h00;      memory[59867] <=  8'h00;      memory[59868] <=  8'h00;      memory[59869] <=  8'h00;      memory[59870] <=  8'h00;      memory[59871] <=  8'h00;      memory[59872] <=  8'h00;      memory[59873] <=  8'h00;      memory[59874] <=  8'h00;      memory[59875] <=  8'h00;      memory[59876] <=  8'h00;      memory[59877] <=  8'h00;      memory[59878] <=  8'h00;      memory[59879] <=  8'h00;      memory[59880] <=  8'h00;      memory[59881] <=  8'h00;      memory[59882] <=  8'h00;      memory[59883] <=  8'h00;      memory[59884] <=  8'h00;      memory[59885] <=  8'h00;      memory[59886] <=  8'h00;      memory[59887] <=  8'h00;      memory[59888] <=  8'h00;      memory[59889] <=  8'h00;      memory[59890] <=  8'h00;      memory[59891] <=  8'h00;      memory[59892] <=  8'h00;      memory[59893] <=  8'h00;      memory[59894] <=  8'h00;      memory[59895] <=  8'h00;      memory[59896] <=  8'h00;      memory[59897] <=  8'h00;      memory[59898] <=  8'h00;      memory[59899] <=  8'h00;      memory[59900] <=  8'h00;      memory[59901] <=  8'h00;      memory[59902] <=  8'h00;      memory[59903] <=  8'h00;      memory[59904] <=  8'h00;      memory[59905] <=  8'h00;      memory[59906] <=  8'h00;      memory[59907] <=  8'h00;      memory[59908] <=  8'h00;      memory[59909] <=  8'h00;      memory[59910] <=  8'h00;      memory[59911] <=  8'h00;      memory[59912] <=  8'h00;      memory[59913] <=  8'h00;      memory[59914] <=  8'h00;      memory[59915] <=  8'h00;      memory[59916] <=  8'h00;      memory[59917] <=  8'h00;      memory[59918] <=  8'h00;      memory[59919] <=  8'h00;      memory[59920] <=  8'h00;      memory[59921] <=  8'h00;      memory[59922] <=  8'h00;      memory[59923] <=  8'h00;      memory[59924] <=  8'h00;      memory[59925] <=  8'h00;      memory[59926] <=  8'h00;      memory[59927] <=  8'h00;      memory[59928] <=  8'h00;      memory[59929] <=  8'h00;      memory[59930] <=  8'h00;      memory[59931] <=  8'h00;      memory[59932] <=  8'h00;      memory[59933] <=  8'h00;      memory[59934] <=  8'h00;      memory[59935] <=  8'h00;      memory[59936] <=  8'h00;      memory[59937] <=  8'h00;      memory[59938] <=  8'h00;      memory[59939] <=  8'h00;      memory[59940] <=  8'h00;      memory[59941] <=  8'h00;      memory[59942] <=  8'h00;      memory[59943] <=  8'h00;      memory[59944] <=  8'h00;      memory[59945] <=  8'h00;      memory[59946] <=  8'h00;      memory[59947] <=  8'h00;      memory[59948] <=  8'h00;      memory[59949] <=  8'h00;      memory[59950] <=  8'h00;      memory[59951] <=  8'h00;      memory[59952] <=  8'h00;      memory[59953] <=  8'h00;      memory[59954] <=  8'h00;      memory[59955] <=  8'h00;      memory[59956] <=  8'h00;      memory[59957] <=  8'h00;      memory[59958] <=  8'h00;      memory[59959] <=  8'h00;      memory[59960] <=  8'h00;      memory[59961] <=  8'h00;      memory[59962] <=  8'h00;      memory[59963] <=  8'h00;      memory[59964] <=  8'h00;      memory[59965] <=  8'h00;      memory[59966] <=  8'h00;      memory[59967] <=  8'h00;      memory[59968] <=  8'h00;      memory[59969] <=  8'h00;      memory[59970] <=  8'h00;      memory[59971] <=  8'h00;      memory[59972] <=  8'h00;      memory[59973] <=  8'h00;      memory[59974] <=  8'h00;      memory[59975] <=  8'h00;      memory[59976] <=  8'h00;      memory[59977] <=  8'h00;      memory[59978] <=  8'h00;      memory[59979] <=  8'h00;      memory[59980] <=  8'h00;      memory[59981] <=  8'h00;      memory[59982] <=  8'h00;      memory[59983] <=  8'h00;      memory[59984] <=  8'h00;      memory[59985] <=  8'h00;      memory[59986] <=  8'h00;      memory[59987] <=  8'h00;      memory[59988] <=  8'h00;      memory[59989] <=  8'h00;      memory[59990] <=  8'h00;      memory[59991] <=  8'h00;      memory[59992] <=  8'h00;      memory[59993] <=  8'h00;      memory[59994] <=  8'h00;      memory[59995] <=  8'h00;      memory[59996] <=  8'h00;      memory[59997] <=  8'h00;      memory[59998] <=  8'h00;      memory[59999] <=  8'h00;      memory[60000] <=  8'h00;      memory[60001] <=  8'h00;      memory[60002] <=  8'h00;      memory[60003] <=  8'h00;      memory[60004] <=  8'h00;      memory[60005] <=  8'h00;      memory[60006] <=  8'h00;      memory[60007] <=  8'h00;      memory[60008] <=  8'h00;      memory[60009] <=  8'h00;      memory[60010] <=  8'h00;      memory[60011] <=  8'h00;      memory[60012] <=  8'h00;      memory[60013] <=  8'h00;      memory[60014] <=  8'h00;      memory[60015] <=  8'h00;      memory[60016] <=  8'h00;      memory[60017] <=  8'h00;      memory[60018] <=  8'h00;      memory[60019] <=  8'h00;      memory[60020] <=  8'h00;      memory[60021] <=  8'h00;      memory[60022] <=  8'h00;      memory[60023] <=  8'h00;      memory[60024] <=  8'h00;      memory[60025] <=  8'h00;      memory[60026] <=  8'h00;      memory[60027] <=  8'h00;      memory[60028] <=  8'h00;      memory[60029] <=  8'h00;      memory[60030] <=  8'h00;      memory[60031] <=  8'h00;      memory[60032] <=  8'h00;      memory[60033] <=  8'h00;      memory[60034] <=  8'h00;      memory[60035] <=  8'h00;      memory[60036] <=  8'h00;      memory[60037] <=  8'h00;      memory[60038] <=  8'h00;      memory[60039] <=  8'h00;      memory[60040] <=  8'h00;      memory[60041] <=  8'h00;      memory[60042] <=  8'h00;      memory[60043] <=  8'h00;      memory[60044] <=  8'h00;      memory[60045] <=  8'h00;      memory[60046] <=  8'h00;      memory[60047] <=  8'h00;      memory[60048] <=  8'h00;      memory[60049] <=  8'h00;      memory[60050] <=  8'h00;      memory[60051] <=  8'h00;      memory[60052] <=  8'h00;      memory[60053] <=  8'h00;      memory[60054] <=  8'h00;      memory[60055] <=  8'h00;      memory[60056] <=  8'h00;      memory[60057] <=  8'h00;      memory[60058] <=  8'h00;      memory[60059] <=  8'h00;      memory[60060] <=  8'h00;      memory[60061] <=  8'h00;      memory[60062] <=  8'h00;      memory[60063] <=  8'h00;      memory[60064] <=  8'h00;      memory[60065] <=  8'h00;      memory[60066] <=  8'h00;      memory[60067] <=  8'h00;      memory[60068] <=  8'h00;      memory[60069] <=  8'h00;      memory[60070] <=  8'h00;      memory[60071] <=  8'h00;      memory[60072] <=  8'h00;      memory[60073] <=  8'h00;      memory[60074] <=  8'h00;      memory[60075] <=  8'h00;      memory[60076] <=  8'h00;      memory[60077] <=  8'h00;      memory[60078] <=  8'h00;      memory[60079] <=  8'h00;      memory[60080] <=  8'h00;      memory[60081] <=  8'h00;      memory[60082] <=  8'h00;      memory[60083] <=  8'h00;      memory[60084] <=  8'h00;      memory[60085] <=  8'h00;      memory[60086] <=  8'h00;      memory[60087] <=  8'h00;      memory[60088] <=  8'h00;      memory[60089] <=  8'h00;      memory[60090] <=  8'h00;      memory[60091] <=  8'h00;      memory[60092] <=  8'h00;      memory[60093] <=  8'h00;      memory[60094] <=  8'h00;      memory[60095] <=  8'h00;      memory[60096] <=  8'h00;      memory[60097] <=  8'h00;      memory[60098] <=  8'h00;      memory[60099] <=  8'h00;      memory[60100] <=  8'h00;      memory[60101] <=  8'h00;      memory[60102] <=  8'h00;      memory[60103] <=  8'h00;      memory[60104] <=  8'h00;      memory[60105] <=  8'h00;      memory[60106] <=  8'h00;      memory[60107] <=  8'h00;      memory[60108] <=  8'h00;      memory[60109] <=  8'h00;      memory[60110] <=  8'h00;      memory[60111] <=  8'h00;      memory[60112] <=  8'h00;      memory[60113] <=  8'h00;      memory[60114] <=  8'h00;      memory[60115] <=  8'h00;      memory[60116] <=  8'h00;      memory[60117] <=  8'h00;      memory[60118] <=  8'h00;      memory[60119] <=  8'h00;      memory[60120] <=  8'h00;      memory[60121] <=  8'h00;      memory[60122] <=  8'h00;      memory[60123] <=  8'h00;      memory[60124] <=  8'h00;      memory[60125] <=  8'h00;      memory[60126] <=  8'h00;      memory[60127] <=  8'h00;      memory[60128] <=  8'h00;      memory[60129] <=  8'h00;      memory[60130] <=  8'h00;      memory[60131] <=  8'h00;      memory[60132] <=  8'h00;      memory[60133] <=  8'h00;      memory[60134] <=  8'h00;      memory[60135] <=  8'h00;      memory[60136] <=  8'h00;      memory[60137] <=  8'h00;      memory[60138] <=  8'h00;      memory[60139] <=  8'h00;      memory[60140] <=  8'h00;      memory[60141] <=  8'h00;      memory[60142] <=  8'h00;      memory[60143] <=  8'h00;      memory[60144] <=  8'h00;      memory[60145] <=  8'h00;      memory[60146] <=  8'h00;      memory[60147] <=  8'h00;      memory[60148] <=  8'h00;      memory[60149] <=  8'h00;      memory[60150] <=  8'h00;      memory[60151] <=  8'h00;      memory[60152] <=  8'h00;      memory[60153] <=  8'h00;      memory[60154] <=  8'h00;      memory[60155] <=  8'h00;      memory[60156] <=  8'h00;      memory[60157] <=  8'h00;      memory[60158] <=  8'h00;      memory[60159] <=  8'h00;      memory[60160] <=  8'h00;      memory[60161] <=  8'h00;      memory[60162] <=  8'h00;      memory[60163] <=  8'h00;      memory[60164] <=  8'h00;      memory[60165] <=  8'h00;      memory[60166] <=  8'h00;      memory[60167] <=  8'h00;      memory[60168] <=  8'h00;      memory[60169] <=  8'h00;      memory[60170] <=  8'h00;      memory[60171] <=  8'h00;      memory[60172] <=  8'h00;      memory[60173] <=  8'h00;      memory[60174] <=  8'h00;      memory[60175] <=  8'h00;      memory[60176] <=  8'h00;      memory[60177] <=  8'h00;      memory[60178] <=  8'h00;      memory[60179] <=  8'h00;      memory[60180] <=  8'h00;      memory[60181] <=  8'h00;      memory[60182] <=  8'h00;      memory[60183] <=  8'h00;      memory[60184] <=  8'h00;      memory[60185] <=  8'h00;      memory[60186] <=  8'h00;      memory[60187] <=  8'h00;      memory[60188] <=  8'h00;      memory[60189] <=  8'h00;      memory[60190] <=  8'h00;      memory[60191] <=  8'h00;      memory[60192] <=  8'h00;      memory[60193] <=  8'h00;      memory[60194] <=  8'h00;      memory[60195] <=  8'h00;      memory[60196] <=  8'h00;      memory[60197] <=  8'h00;      memory[60198] <=  8'h00;      memory[60199] <=  8'h00;      memory[60200] <=  8'h00;      memory[60201] <=  8'h00;      memory[60202] <=  8'h00;      memory[60203] <=  8'h00;      memory[60204] <=  8'h00;      memory[60205] <=  8'h00;      memory[60206] <=  8'h00;      memory[60207] <=  8'h00;      memory[60208] <=  8'h00;      memory[60209] <=  8'h00;      memory[60210] <=  8'h00;      memory[60211] <=  8'h00;      memory[60212] <=  8'h00;      memory[60213] <=  8'h00;      memory[60214] <=  8'h00;      memory[60215] <=  8'h00;      memory[60216] <=  8'h00;      memory[60217] <=  8'h00;      memory[60218] <=  8'h00;      memory[60219] <=  8'h00;      memory[60220] <=  8'h00;      memory[60221] <=  8'h00;      memory[60222] <=  8'h00;      memory[60223] <=  8'h00;      memory[60224] <=  8'h00;      memory[60225] <=  8'h00;      memory[60226] <=  8'h00;      memory[60227] <=  8'h00;      memory[60228] <=  8'h00;      memory[60229] <=  8'h00;      memory[60230] <=  8'h00;      memory[60231] <=  8'h00;      memory[60232] <=  8'h00;      memory[60233] <=  8'h00;      memory[60234] <=  8'h00;      memory[60235] <=  8'h00;      memory[60236] <=  8'h00;      memory[60237] <=  8'h00;      memory[60238] <=  8'h00;      memory[60239] <=  8'h00;      memory[60240] <=  8'h00;      memory[60241] <=  8'h00;      memory[60242] <=  8'h00;      memory[60243] <=  8'h00;      memory[60244] <=  8'h00;      memory[60245] <=  8'h00;      memory[60246] <=  8'h00;      memory[60247] <=  8'h00;      memory[60248] <=  8'h00;      memory[60249] <=  8'h00;      memory[60250] <=  8'h00;      memory[60251] <=  8'h00;      memory[60252] <=  8'h00;      memory[60253] <=  8'h00;      memory[60254] <=  8'h00;      memory[60255] <=  8'h00;      memory[60256] <=  8'h00;      memory[60257] <=  8'h00;      memory[60258] <=  8'h00;      memory[60259] <=  8'h00;      memory[60260] <=  8'h00;      memory[60261] <=  8'h00;      memory[60262] <=  8'h00;      memory[60263] <=  8'h00;      memory[60264] <=  8'h00;      memory[60265] <=  8'h00;      memory[60266] <=  8'h00;      memory[60267] <=  8'h00;      memory[60268] <=  8'h00;      memory[60269] <=  8'h00;      memory[60270] <=  8'h00;      memory[60271] <=  8'h00;      memory[60272] <=  8'h00;      memory[60273] <=  8'h00;      memory[60274] <=  8'h00;      memory[60275] <=  8'h00;      memory[60276] <=  8'h00;      memory[60277] <=  8'h00;      memory[60278] <=  8'h00;      memory[60279] <=  8'h00;      memory[60280] <=  8'h00;      memory[60281] <=  8'h00;      memory[60282] <=  8'h00;      memory[60283] <=  8'h00;      memory[60284] <=  8'h00;      memory[60285] <=  8'h00;      memory[60286] <=  8'h00;      memory[60287] <=  8'h00;      memory[60288] <=  8'h00;      memory[60289] <=  8'h00;      memory[60290] <=  8'h00;      memory[60291] <=  8'h00;      memory[60292] <=  8'h00;      memory[60293] <=  8'h00;      memory[60294] <=  8'h00;      memory[60295] <=  8'h00;      memory[60296] <=  8'h00;      memory[60297] <=  8'h00;      memory[60298] <=  8'h00;      memory[60299] <=  8'h00;      memory[60300] <=  8'h00;      memory[60301] <=  8'h00;      memory[60302] <=  8'h00;      memory[60303] <=  8'h00;      memory[60304] <=  8'h00;      memory[60305] <=  8'h00;      memory[60306] <=  8'h00;      memory[60307] <=  8'h00;      memory[60308] <=  8'h00;      memory[60309] <=  8'h00;      memory[60310] <=  8'h00;      memory[60311] <=  8'h00;      memory[60312] <=  8'h00;      memory[60313] <=  8'h00;      memory[60314] <=  8'h00;      memory[60315] <=  8'h00;      memory[60316] <=  8'h00;      memory[60317] <=  8'h00;      memory[60318] <=  8'h00;      memory[60319] <=  8'h00;      memory[60320] <=  8'h00;      memory[60321] <=  8'h00;      memory[60322] <=  8'h00;      memory[60323] <=  8'h00;      memory[60324] <=  8'h00;      memory[60325] <=  8'h00;      memory[60326] <=  8'h00;      memory[60327] <=  8'h00;      memory[60328] <=  8'h00;      memory[60329] <=  8'h00;      memory[60330] <=  8'h00;      memory[60331] <=  8'h00;      memory[60332] <=  8'h00;      memory[60333] <=  8'h00;      memory[60334] <=  8'h00;      memory[60335] <=  8'h00;      memory[60336] <=  8'h00;      memory[60337] <=  8'h00;      memory[60338] <=  8'h00;      memory[60339] <=  8'h00;      memory[60340] <=  8'h00;      memory[60341] <=  8'h00;      memory[60342] <=  8'h00;      memory[60343] <=  8'h00;      memory[60344] <=  8'h00;      memory[60345] <=  8'h00;      memory[60346] <=  8'h00;      memory[60347] <=  8'h00;      memory[60348] <=  8'h00;      memory[60349] <=  8'h00;      memory[60350] <=  8'h00;      memory[60351] <=  8'h00;      memory[60352] <=  8'h00;      memory[60353] <=  8'h00;      memory[60354] <=  8'h00;      memory[60355] <=  8'h00;      memory[60356] <=  8'h00;      memory[60357] <=  8'h00;      memory[60358] <=  8'h00;      memory[60359] <=  8'h00;      memory[60360] <=  8'h00;      memory[60361] <=  8'h00;      memory[60362] <=  8'h00;      memory[60363] <=  8'h00;      memory[60364] <=  8'h00;      memory[60365] <=  8'h00;      memory[60366] <=  8'h00;      memory[60367] <=  8'h00;      memory[60368] <=  8'h00;      memory[60369] <=  8'h00;      memory[60370] <=  8'h00;      memory[60371] <=  8'h00;      memory[60372] <=  8'h00;      memory[60373] <=  8'h00;      memory[60374] <=  8'h00;      memory[60375] <=  8'h00;      memory[60376] <=  8'h00;      memory[60377] <=  8'h00;      memory[60378] <=  8'h00;      memory[60379] <=  8'h00;      memory[60380] <=  8'h00;      memory[60381] <=  8'h00;      memory[60382] <=  8'h00;      memory[60383] <=  8'h00;      memory[60384] <=  8'h00;      memory[60385] <=  8'h00;      memory[60386] <=  8'h00;      memory[60387] <=  8'h00;      memory[60388] <=  8'h00;      memory[60389] <=  8'h00;      memory[60390] <=  8'h00;      memory[60391] <=  8'h00;      memory[60392] <=  8'h00;      memory[60393] <=  8'h00;      memory[60394] <=  8'h00;      memory[60395] <=  8'h00;      memory[60396] <=  8'h00;      memory[60397] <=  8'h00;      memory[60398] <=  8'h00;      memory[60399] <=  8'h00;      memory[60400] <=  8'h00;      memory[60401] <=  8'h00;      memory[60402] <=  8'h00;      memory[60403] <=  8'h00;      memory[60404] <=  8'h00;      memory[60405] <=  8'h00;      memory[60406] <=  8'h00;      memory[60407] <=  8'h00;      memory[60408] <=  8'h00;      memory[60409] <=  8'h00;      memory[60410] <=  8'h00;      memory[60411] <=  8'h00;      memory[60412] <=  8'h00;      memory[60413] <=  8'h00;      memory[60414] <=  8'h00;      memory[60415] <=  8'h00;      memory[60416] <=  8'h00;      memory[60417] <=  8'h00;      memory[60418] <=  8'h00;      memory[60419] <=  8'h00;      memory[60420] <=  8'h00;      memory[60421] <=  8'h00;      memory[60422] <=  8'h00;      memory[60423] <=  8'h00;      memory[60424] <=  8'h00;      memory[60425] <=  8'h00;      memory[60426] <=  8'h00;      memory[60427] <=  8'h00;      memory[60428] <=  8'h00;      memory[60429] <=  8'h00;      memory[60430] <=  8'h00;      memory[60431] <=  8'h00;      memory[60432] <=  8'h00;      memory[60433] <=  8'h00;      memory[60434] <=  8'h00;      memory[60435] <=  8'h00;      memory[60436] <=  8'h00;      memory[60437] <=  8'h00;      memory[60438] <=  8'h00;      memory[60439] <=  8'h00;      memory[60440] <=  8'h00;      memory[60441] <=  8'h00;      memory[60442] <=  8'h00;      memory[60443] <=  8'h00;      memory[60444] <=  8'h00;      memory[60445] <=  8'h00;      memory[60446] <=  8'h00;      memory[60447] <=  8'h00;      memory[60448] <=  8'h00;      memory[60449] <=  8'h00;      memory[60450] <=  8'h00;      memory[60451] <=  8'h00;      memory[60452] <=  8'h00;      memory[60453] <=  8'h00;      memory[60454] <=  8'h00;      memory[60455] <=  8'h00;      memory[60456] <=  8'h00;      memory[60457] <=  8'h00;      memory[60458] <=  8'h00;      memory[60459] <=  8'h00;      memory[60460] <=  8'h00;      memory[60461] <=  8'h00;      memory[60462] <=  8'h00;      memory[60463] <=  8'h00;      memory[60464] <=  8'h00;      memory[60465] <=  8'h00;      memory[60466] <=  8'h00;      memory[60467] <=  8'h00;      memory[60468] <=  8'h00;      memory[60469] <=  8'h00;      memory[60470] <=  8'h00;      memory[60471] <=  8'h00;      memory[60472] <=  8'h00;      memory[60473] <=  8'h00;      memory[60474] <=  8'h00;      memory[60475] <=  8'h00;      memory[60476] <=  8'h00;      memory[60477] <=  8'h00;      memory[60478] <=  8'h00;      memory[60479] <=  8'h00;      memory[60480] <=  8'h00;      memory[60481] <=  8'h00;      memory[60482] <=  8'h00;      memory[60483] <=  8'h00;      memory[60484] <=  8'h00;      memory[60485] <=  8'h00;      memory[60486] <=  8'h00;      memory[60487] <=  8'h00;      memory[60488] <=  8'h00;      memory[60489] <=  8'h00;      memory[60490] <=  8'h00;      memory[60491] <=  8'h00;      memory[60492] <=  8'h00;      memory[60493] <=  8'h00;      memory[60494] <=  8'h00;      memory[60495] <=  8'h00;      memory[60496] <=  8'h00;      memory[60497] <=  8'h00;      memory[60498] <=  8'h00;      memory[60499] <=  8'h00;      memory[60500] <=  8'h00;      memory[60501] <=  8'h00;      memory[60502] <=  8'h00;      memory[60503] <=  8'h00;      memory[60504] <=  8'h00;      memory[60505] <=  8'h00;      memory[60506] <=  8'h00;      memory[60507] <=  8'h00;      memory[60508] <=  8'h00;      memory[60509] <=  8'h00;      memory[60510] <=  8'h00;      memory[60511] <=  8'h00;      memory[60512] <=  8'h00;      memory[60513] <=  8'h00;      memory[60514] <=  8'h00;      memory[60515] <=  8'h00;      memory[60516] <=  8'h00;      memory[60517] <=  8'h00;      memory[60518] <=  8'h00;      memory[60519] <=  8'h00;      memory[60520] <=  8'h00;      memory[60521] <=  8'h00;      memory[60522] <=  8'h00;      memory[60523] <=  8'h00;      memory[60524] <=  8'h00;      memory[60525] <=  8'h00;      memory[60526] <=  8'h00;      memory[60527] <=  8'h00;      memory[60528] <=  8'h00;      memory[60529] <=  8'h00;      memory[60530] <=  8'h00;      memory[60531] <=  8'h00;      memory[60532] <=  8'h00;      memory[60533] <=  8'h00;      memory[60534] <=  8'h00;      memory[60535] <=  8'h00;      memory[60536] <=  8'h00;      memory[60537] <=  8'h00;      memory[60538] <=  8'h00;      memory[60539] <=  8'h00;      memory[60540] <=  8'h00;      memory[60541] <=  8'h00;      memory[60542] <=  8'h00;      memory[60543] <=  8'h00;      memory[60544] <=  8'h00;      memory[60545] <=  8'h00;      memory[60546] <=  8'h00;      memory[60547] <=  8'h00;      memory[60548] <=  8'h00;      memory[60549] <=  8'h00;      memory[60550] <=  8'h00;      memory[60551] <=  8'h00;      memory[60552] <=  8'h00;      memory[60553] <=  8'h00;      memory[60554] <=  8'h00;      memory[60555] <=  8'h00;      memory[60556] <=  8'h00;      memory[60557] <=  8'h00;      memory[60558] <=  8'h00;      memory[60559] <=  8'h00;      memory[60560] <=  8'h00;      memory[60561] <=  8'h00;      memory[60562] <=  8'h00;      memory[60563] <=  8'h00;      memory[60564] <=  8'h00;      memory[60565] <=  8'h00;      memory[60566] <=  8'h00;      memory[60567] <=  8'h00;      memory[60568] <=  8'h00;      memory[60569] <=  8'h00;      memory[60570] <=  8'h00;      memory[60571] <=  8'h00;      memory[60572] <=  8'h00;      memory[60573] <=  8'h00;      memory[60574] <=  8'h00;      memory[60575] <=  8'h00;      memory[60576] <=  8'h00;      memory[60577] <=  8'h00;      memory[60578] <=  8'h00;      memory[60579] <=  8'h00;      memory[60580] <=  8'h00;      memory[60581] <=  8'h00;      memory[60582] <=  8'h00;      memory[60583] <=  8'h00;      memory[60584] <=  8'h00;      memory[60585] <=  8'h00;      memory[60586] <=  8'h00;      memory[60587] <=  8'h00;      memory[60588] <=  8'h00;      memory[60589] <=  8'h00;      memory[60590] <=  8'h00;      memory[60591] <=  8'h00;      memory[60592] <=  8'h00;      memory[60593] <=  8'h00;      memory[60594] <=  8'h00;      memory[60595] <=  8'h00;      memory[60596] <=  8'h00;      memory[60597] <=  8'h00;      memory[60598] <=  8'h00;      memory[60599] <=  8'h00;      memory[60600] <=  8'h00;      memory[60601] <=  8'h00;      memory[60602] <=  8'h00;      memory[60603] <=  8'h00;      memory[60604] <=  8'h00;      memory[60605] <=  8'h00;      memory[60606] <=  8'h00;      memory[60607] <=  8'h00;      memory[60608] <=  8'h00;      memory[60609] <=  8'h00;      memory[60610] <=  8'h00;      memory[60611] <=  8'h00;      memory[60612] <=  8'h00;      memory[60613] <=  8'h00;      memory[60614] <=  8'h00;      memory[60615] <=  8'h00;      memory[60616] <=  8'h00;      memory[60617] <=  8'h00;      memory[60618] <=  8'h00;      memory[60619] <=  8'h00;      memory[60620] <=  8'h00;      memory[60621] <=  8'h00;      memory[60622] <=  8'h00;      memory[60623] <=  8'h00;      memory[60624] <=  8'h00;      memory[60625] <=  8'h00;      memory[60626] <=  8'h00;      memory[60627] <=  8'h00;      memory[60628] <=  8'h00;      memory[60629] <=  8'h00;      memory[60630] <=  8'h00;      memory[60631] <=  8'h00;      memory[60632] <=  8'h00;      memory[60633] <=  8'h00;      memory[60634] <=  8'h00;      memory[60635] <=  8'h00;      memory[60636] <=  8'h00;      memory[60637] <=  8'h00;      memory[60638] <=  8'h00;      memory[60639] <=  8'h00;      memory[60640] <=  8'h00;      memory[60641] <=  8'h00;      memory[60642] <=  8'h00;      memory[60643] <=  8'h00;      memory[60644] <=  8'h00;      memory[60645] <=  8'h00;      memory[60646] <=  8'h00;      memory[60647] <=  8'h00;      memory[60648] <=  8'h00;      memory[60649] <=  8'h00;      memory[60650] <=  8'h00;      memory[60651] <=  8'h00;      memory[60652] <=  8'h00;      memory[60653] <=  8'h00;      memory[60654] <=  8'h00;      memory[60655] <=  8'h00;      memory[60656] <=  8'h00;      memory[60657] <=  8'h00;      memory[60658] <=  8'h00;      memory[60659] <=  8'h00;      memory[60660] <=  8'h00;      memory[60661] <=  8'h00;      memory[60662] <=  8'h00;      memory[60663] <=  8'h00;      memory[60664] <=  8'h00;      memory[60665] <=  8'h00;      memory[60666] <=  8'h00;      memory[60667] <=  8'h00;      memory[60668] <=  8'h00;      memory[60669] <=  8'h00;      memory[60670] <=  8'h00;      memory[60671] <=  8'h00;      memory[60672] <=  8'h00;      memory[60673] <=  8'h00;      memory[60674] <=  8'h00;      memory[60675] <=  8'h00;      memory[60676] <=  8'h00;      memory[60677] <=  8'h00;      memory[60678] <=  8'h00;      memory[60679] <=  8'h00;      memory[60680] <=  8'h00;      memory[60681] <=  8'h00;      memory[60682] <=  8'h00;      memory[60683] <=  8'h00;      memory[60684] <=  8'h00;      memory[60685] <=  8'h00;      memory[60686] <=  8'h00;      memory[60687] <=  8'h00;      memory[60688] <=  8'h00;      memory[60689] <=  8'h00;      memory[60690] <=  8'h00;      memory[60691] <=  8'h00;      memory[60692] <=  8'h00;      memory[60693] <=  8'h00;      memory[60694] <=  8'h00;      memory[60695] <=  8'h00;      memory[60696] <=  8'h00;      memory[60697] <=  8'h00;      memory[60698] <=  8'h00;      memory[60699] <=  8'h00;      memory[60700] <=  8'h00;      memory[60701] <=  8'h00;      memory[60702] <=  8'h00;      memory[60703] <=  8'h00;      memory[60704] <=  8'h00;      memory[60705] <=  8'h00;      memory[60706] <=  8'h00;      memory[60707] <=  8'h00;      memory[60708] <=  8'h00;      memory[60709] <=  8'h00;      memory[60710] <=  8'h00;      memory[60711] <=  8'h00;      memory[60712] <=  8'h00;      memory[60713] <=  8'h00;      memory[60714] <=  8'h00;      memory[60715] <=  8'h00;      memory[60716] <=  8'h00;      memory[60717] <=  8'h00;      memory[60718] <=  8'h00;      memory[60719] <=  8'h00;      memory[60720] <=  8'h00;      memory[60721] <=  8'h00;      memory[60722] <=  8'h00;      memory[60723] <=  8'h00;      memory[60724] <=  8'h00;      memory[60725] <=  8'h00;      memory[60726] <=  8'h00;      memory[60727] <=  8'h00;      memory[60728] <=  8'h00;      memory[60729] <=  8'h00;      memory[60730] <=  8'h00;      memory[60731] <=  8'h00;      memory[60732] <=  8'h00;      memory[60733] <=  8'h00;      memory[60734] <=  8'h00;      memory[60735] <=  8'h00;      memory[60736] <=  8'h00;      memory[60737] <=  8'h00;      memory[60738] <=  8'h00;      memory[60739] <=  8'h00;      memory[60740] <=  8'h00;      memory[60741] <=  8'h00;      memory[60742] <=  8'h00;      memory[60743] <=  8'h00;      memory[60744] <=  8'h00;      memory[60745] <=  8'h00;      memory[60746] <=  8'h00;      memory[60747] <=  8'h00;      memory[60748] <=  8'h00;      memory[60749] <=  8'h00;      memory[60750] <=  8'h00;      memory[60751] <=  8'h00;      memory[60752] <=  8'h00;      memory[60753] <=  8'h00;      memory[60754] <=  8'h00;      memory[60755] <=  8'h00;      memory[60756] <=  8'h00;      memory[60757] <=  8'h00;      memory[60758] <=  8'h00;      memory[60759] <=  8'h00;      memory[60760] <=  8'h00;      memory[60761] <=  8'h00;      memory[60762] <=  8'h00;      memory[60763] <=  8'h00;      memory[60764] <=  8'h00;      memory[60765] <=  8'h00;      memory[60766] <=  8'h00;      memory[60767] <=  8'h00;      memory[60768] <=  8'h00;      memory[60769] <=  8'h00;      memory[60770] <=  8'h00;      memory[60771] <=  8'h00;      memory[60772] <=  8'h00;      memory[60773] <=  8'h00;      memory[60774] <=  8'h00;      memory[60775] <=  8'h00;      memory[60776] <=  8'h00;      memory[60777] <=  8'h00;      memory[60778] <=  8'h00;      memory[60779] <=  8'h00;      memory[60780] <=  8'h00;      memory[60781] <=  8'h00;      memory[60782] <=  8'h00;      memory[60783] <=  8'h00;      memory[60784] <=  8'h00;      memory[60785] <=  8'h00;      memory[60786] <=  8'h00;      memory[60787] <=  8'h00;      memory[60788] <=  8'h00;      memory[60789] <=  8'h00;      memory[60790] <=  8'h00;      memory[60791] <=  8'h00;      memory[60792] <=  8'h00;      memory[60793] <=  8'h00;      memory[60794] <=  8'h00;      memory[60795] <=  8'h00;      memory[60796] <=  8'h00;      memory[60797] <=  8'h00;      memory[60798] <=  8'h00;      memory[60799] <=  8'h00;      memory[60800] <=  8'h00;      memory[60801] <=  8'h00;      memory[60802] <=  8'h00;      memory[60803] <=  8'h00;      memory[60804] <=  8'h00;      memory[60805] <=  8'h00;      memory[60806] <=  8'h00;      memory[60807] <=  8'h00;      memory[60808] <=  8'h00;      memory[60809] <=  8'h00;      memory[60810] <=  8'h00;      memory[60811] <=  8'h00;      memory[60812] <=  8'h00;      memory[60813] <=  8'h00;      memory[60814] <=  8'h00;      memory[60815] <=  8'h00;      memory[60816] <=  8'h00;      memory[60817] <=  8'h00;      memory[60818] <=  8'h00;      memory[60819] <=  8'h00;      memory[60820] <=  8'h00;      memory[60821] <=  8'h00;      memory[60822] <=  8'h00;      memory[60823] <=  8'h00;      memory[60824] <=  8'h00;      memory[60825] <=  8'h00;      memory[60826] <=  8'h00;      memory[60827] <=  8'h00;      memory[60828] <=  8'h00;      memory[60829] <=  8'h00;      memory[60830] <=  8'h00;      memory[60831] <=  8'h00;      memory[60832] <=  8'h00;      memory[60833] <=  8'h00;      memory[60834] <=  8'h00;      memory[60835] <=  8'h00;      memory[60836] <=  8'h00;      memory[60837] <=  8'h00;      memory[60838] <=  8'h00;      memory[60839] <=  8'h00;      memory[60840] <=  8'h00;      memory[60841] <=  8'h00;      memory[60842] <=  8'h00;      memory[60843] <=  8'h00;      memory[60844] <=  8'h00;      memory[60845] <=  8'h00;      memory[60846] <=  8'h00;      memory[60847] <=  8'h00;      memory[60848] <=  8'h00;      memory[60849] <=  8'h00;      memory[60850] <=  8'h00;      memory[60851] <=  8'h00;      memory[60852] <=  8'h00;      memory[60853] <=  8'h00;      memory[60854] <=  8'h00;      memory[60855] <=  8'h00;      memory[60856] <=  8'h00;      memory[60857] <=  8'h00;      memory[60858] <=  8'h00;      memory[60859] <=  8'h00;      memory[60860] <=  8'h00;      memory[60861] <=  8'h00;      memory[60862] <=  8'h00;      memory[60863] <=  8'h00;      memory[60864] <=  8'h00;      memory[60865] <=  8'h00;      memory[60866] <=  8'h00;      memory[60867] <=  8'h00;      memory[60868] <=  8'h00;      memory[60869] <=  8'h00;      memory[60870] <=  8'h00;      memory[60871] <=  8'h00;      memory[60872] <=  8'h00;      memory[60873] <=  8'h00;      memory[60874] <=  8'h00;      memory[60875] <=  8'h00;      memory[60876] <=  8'h00;      memory[60877] <=  8'h00;      memory[60878] <=  8'h00;      memory[60879] <=  8'h00;      memory[60880] <=  8'h00;      memory[60881] <=  8'h00;      memory[60882] <=  8'h00;      memory[60883] <=  8'h00;      memory[60884] <=  8'h00;      memory[60885] <=  8'h00;      memory[60886] <=  8'h00;      memory[60887] <=  8'h00;      memory[60888] <=  8'h00;      memory[60889] <=  8'h00;      memory[60890] <=  8'h00;      memory[60891] <=  8'h00;      memory[60892] <=  8'h00;      memory[60893] <=  8'h00;      memory[60894] <=  8'h00;      memory[60895] <=  8'h00;      memory[60896] <=  8'h00;      memory[60897] <=  8'h00;      memory[60898] <=  8'h00;      memory[60899] <=  8'h00;      memory[60900] <=  8'h00;      memory[60901] <=  8'h00;      memory[60902] <=  8'h00;      memory[60903] <=  8'h00;      memory[60904] <=  8'h00;      memory[60905] <=  8'h00;      memory[60906] <=  8'h00;      memory[60907] <=  8'h00;      memory[60908] <=  8'h00;      memory[60909] <=  8'h00;      memory[60910] <=  8'h00;      memory[60911] <=  8'h00;      memory[60912] <=  8'h00;      memory[60913] <=  8'h00;      memory[60914] <=  8'h00;      memory[60915] <=  8'h00;      memory[60916] <=  8'h00;      memory[60917] <=  8'h00;      memory[60918] <=  8'h00;      memory[60919] <=  8'h00;      memory[60920] <=  8'h00;      memory[60921] <=  8'h00;      memory[60922] <=  8'h00;      memory[60923] <=  8'h00;      memory[60924] <=  8'h00;      memory[60925] <=  8'h00;      memory[60926] <=  8'h00;      memory[60927] <=  8'h00;      memory[60928] <=  8'h00;      memory[60929] <=  8'h00;      memory[60930] <=  8'h00;      memory[60931] <=  8'h00;      memory[60932] <=  8'h00;      memory[60933] <=  8'h00;      memory[60934] <=  8'h00;      memory[60935] <=  8'h00;      memory[60936] <=  8'h00;      memory[60937] <=  8'h00;      memory[60938] <=  8'h00;      memory[60939] <=  8'h00;      memory[60940] <=  8'h00;      memory[60941] <=  8'h00;      memory[60942] <=  8'h00;      memory[60943] <=  8'h00;      memory[60944] <=  8'h00;      memory[60945] <=  8'h00;      memory[60946] <=  8'h00;      memory[60947] <=  8'h00;      memory[60948] <=  8'h00;      memory[60949] <=  8'h00;      memory[60950] <=  8'h00;      memory[60951] <=  8'h00;      memory[60952] <=  8'h00;      memory[60953] <=  8'h00;      memory[60954] <=  8'h00;      memory[60955] <=  8'h00;      memory[60956] <=  8'h00;      memory[60957] <=  8'h00;      memory[60958] <=  8'h00;      memory[60959] <=  8'h00;      memory[60960] <=  8'h00;      memory[60961] <=  8'h00;      memory[60962] <=  8'h00;      memory[60963] <=  8'h00;      memory[60964] <=  8'h00;      memory[60965] <=  8'h00;      memory[60966] <=  8'h00;      memory[60967] <=  8'h00;      memory[60968] <=  8'h00;      memory[60969] <=  8'h00;      memory[60970] <=  8'h00;      memory[60971] <=  8'h00;      memory[60972] <=  8'h00;      memory[60973] <=  8'h00;      memory[60974] <=  8'h00;      memory[60975] <=  8'h00;      memory[60976] <=  8'h00;      memory[60977] <=  8'h00;      memory[60978] <=  8'h00;      memory[60979] <=  8'h00;      memory[60980] <=  8'h00;      memory[60981] <=  8'h00;      memory[60982] <=  8'h00;      memory[60983] <=  8'h00;      memory[60984] <=  8'h00;      memory[60985] <=  8'h00;      memory[60986] <=  8'h00;      memory[60987] <=  8'h00;      memory[60988] <=  8'h00;      memory[60989] <=  8'h00;      memory[60990] <=  8'h00;      memory[60991] <=  8'h00;      memory[60992] <=  8'h00;      memory[60993] <=  8'h00;      memory[60994] <=  8'h00;      memory[60995] <=  8'h00;      memory[60996] <=  8'h00;      memory[60997] <=  8'h00;      memory[60998] <=  8'h00;      memory[60999] <=  8'h00;      memory[61000] <=  8'h00;      memory[61001] <=  8'h00;      memory[61002] <=  8'h00;      memory[61003] <=  8'h00;      memory[61004] <=  8'h00;      memory[61005] <=  8'h00;      memory[61006] <=  8'h00;      memory[61007] <=  8'h00;      memory[61008] <=  8'h00;      memory[61009] <=  8'h00;      memory[61010] <=  8'h00;      memory[61011] <=  8'h00;      memory[61012] <=  8'h00;      memory[61013] <=  8'h00;      memory[61014] <=  8'h00;      memory[61015] <=  8'h00;      memory[61016] <=  8'h00;      memory[61017] <=  8'h00;      memory[61018] <=  8'h00;      memory[61019] <=  8'h00;      memory[61020] <=  8'h00;      memory[61021] <=  8'h00;      memory[61022] <=  8'h00;      memory[61023] <=  8'h00;      memory[61024] <=  8'h00;      memory[61025] <=  8'h00;      memory[61026] <=  8'h00;      memory[61027] <=  8'h00;      memory[61028] <=  8'h00;      memory[61029] <=  8'h00;      memory[61030] <=  8'h00;      memory[61031] <=  8'h00;      memory[61032] <=  8'h00;      memory[61033] <=  8'h00;      memory[61034] <=  8'h00;      memory[61035] <=  8'h00;      memory[61036] <=  8'h00;      memory[61037] <=  8'h00;      memory[61038] <=  8'h00;      memory[61039] <=  8'h00;      memory[61040] <=  8'h00;      memory[61041] <=  8'h00;      memory[61042] <=  8'h00;      memory[61043] <=  8'h00;      memory[61044] <=  8'h00;      memory[61045] <=  8'h00;      memory[61046] <=  8'h00;      memory[61047] <=  8'h00;      memory[61048] <=  8'h00;      memory[61049] <=  8'h00;      memory[61050] <=  8'h00;      memory[61051] <=  8'h00;      memory[61052] <=  8'h00;      memory[61053] <=  8'h00;      memory[61054] <=  8'h00;      memory[61055] <=  8'h00;      memory[61056] <=  8'h00;      memory[61057] <=  8'h00;      memory[61058] <=  8'h00;      memory[61059] <=  8'h00;      memory[61060] <=  8'h00;      memory[61061] <=  8'h00;      memory[61062] <=  8'h00;      memory[61063] <=  8'h00;      memory[61064] <=  8'h00;      memory[61065] <=  8'h00;      memory[61066] <=  8'h00;      memory[61067] <=  8'h00;      memory[61068] <=  8'h00;      memory[61069] <=  8'h00;      memory[61070] <=  8'h00;      memory[61071] <=  8'h00;      memory[61072] <=  8'h00;      memory[61073] <=  8'h00;      memory[61074] <=  8'h00;      memory[61075] <=  8'h00;      memory[61076] <=  8'h00;      memory[61077] <=  8'h00;      memory[61078] <=  8'h00;      memory[61079] <=  8'h00;      memory[61080] <=  8'h00;      memory[61081] <=  8'h00;      memory[61082] <=  8'h00;      memory[61083] <=  8'h00;      memory[61084] <=  8'h00;      memory[61085] <=  8'h00;      memory[61086] <=  8'h00;      memory[61087] <=  8'h00;      memory[61088] <=  8'h00;      memory[61089] <=  8'h00;      memory[61090] <=  8'h00;      memory[61091] <=  8'h00;      memory[61092] <=  8'h00;      memory[61093] <=  8'h00;      memory[61094] <=  8'h00;      memory[61095] <=  8'h00;      memory[61096] <=  8'h00;      memory[61097] <=  8'h00;      memory[61098] <=  8'h00;      memory[61099] <=  8'h00;      memory[61100] <=  8'h00;      memory[61101] <=  8'h00;      memory[61102] <=  8'h00;      memory[61103] <=  8'h00;      memory[61104] <=  8'h00;      memory[61105] <=  8'h00;      memory[61106] <=  8'h00;      memory[61107] <=  8'h00;      memory[61108] <=  8'h00;      memory[61109] <=  8'h00;      memory[61110] <=  8'h00;      memory[61111] <=  8'h00;      memory[61112] <=  8'h00;      memory[61113] <=  8'h00;      memory[61114] <=  8'h00;      memory[61115] <=  8'h00;      memory[61116] <=  8'h00;      memory[61117] <=  8'h00;      memory[61118] <=  8'h00;      memory[61119] <=  8'h00;      memory[61120] <=  8'h00;      memory[61121] <=  8'h00;      memory[61122] <=  8'h00;      memory[61123] <=  8'h00;      memory[61124] <=  8'h00;      memory[61125] <=  8'h00;      memory[61126] <=  8'h00;      memory[61127] <=  8'h00;      memory[61128] <=  8'h00;      memory[61129] <=  8'h00;      memory[61130] <=  8'h00;      memory[61131] <=  8'h00;      memory[61132] <=  8'h00;      memory[61133] <=  8'h00;      memory[61134] <=  8'h00;      memory[61135] <=  8'h00;      memory[61136] <=  8'h00;      memory[61137] <=  8'h00;      memory[61138] <=  8'h00;      memory[61139] <=  8'h00;      memory[61140] <=  8'h00;      memory[61141] <=  8'h00;      memory[61142] <=  8'h00;      memory[61143] <=  8'h00;      memory[61144] <=  8'h00;      memory[61145] <=  8'h00;      memory[61146] <=  8'h00;      memory[61147] <=  8'h00;      memory[61148] <=  8'h00;      memory[61149] <=  8'h00;      memory[61150] <=  8'h00;      memory[61151] <=  8'h00;      memory[61152] <=  8'h00;      memory[61153] <=  8'h00;      memory[61154] <=  8'h00;      memory[61155] <=  8'h00;      memory[61156] <=  8'h00;      memory[61157] <=  8'h00;      memory[61158] <=  8'h00;      memory[61159] <=  8'h00;      memory[61160] <=  8'h00;      memory[61161] <=  8'h00;      memory[61162] <=  8'h00;      memory[61163] <=  8'h00;      memory[61164] <=  8'h00;      memory[61165] <=  8'h00;      memory[61166] <=  8'h00;      memory[61167] <=  8'h00;      memory[61168] <=  8'h00;      memory[61169] <=  8'h00;      memory[61170] <=  8'h00;      memory[61171] <=  8'h00;      memory[61172] <=  8'h00;      memory[61173] <=  8'h00;      memory[61174] <=  8'h00;      memory[61175] <=  8'h00;      memory[61176] <=  8'h00;      memory[61177] <=  8'h00;      memory[61178] <=  8'h00;      memory[61179] <=  8'h00;      memory[61180] <=  8'h00;      memory[61181] <=  8'h00;      memory[61182] <=  8'h00;      memory[61183] <=  8'h00;      memory[61184] <=  8'h00;      memory[61185] <=  8'h00;      memory[61186] <=  8'h00;      memory[61187] <=  8'h00;      memory[61188] <=  8'h00;      memory[61189] <=  8'h00;      memory[61190] <=  8'h00;      memory[61191] <=  8'h00;      memory[61192] <=  8'h00;      memory[61193] <=  8'h00;      memory[61194] <=  8'h00;      memory[61195] <=  8'h00;      memory[61196] <=  8'h00;      memory[61197] <=  8'h00;      memory[61198] <=  8'h00;      memory[61199] <=  8'h00;      memory[61200] <=  8'h00;      memory[61201] <=  8'h00;      memory[61202] <=  8'h00;      memory[61203] <=  8'h00;      memory[61204] <=  8'h00;      memory[61205] <=  8'h00;      memory[61206] <=  8'h00;      memory[61207] <=  8'h00;      memory[61208] <=  8'h00;      memory[61209] <=  8'h00;      memory[61210] <=  8'h00;      memory[61211] <=  8'h00;      memory[61212] <=  8'h00;      memory[61213] <=  8'h00;      memory[61214] <=  8'h00;      memory[61215] <=  8'h00;      memory[61216] <=  8'h00;      memory[61217] <=  8'h00;      memory[61218] <=  8'h00;      memory[61219] <=  8'h00;      memory[61220] <=  8'h00;      memory[61221] <=  8'h00;      memory[61222] <=  8'h00;      memory[61223] <=  8'h00;      memory[61224] <=  8'h00;      memory[61225] <=  8'h00;      memory[61226] <=  8'h00;      memory[61227] <=  8'h00;      memory[61228] <=  8'h00;      memory[61229] <=  8'h00;      memory[61230] <=  8'h00;      memory[61231] <=  8'h00;      memory[61232] <=  8'h00;      memory[61233] <=  8'h00;      memory[61234] <=  8'h00;      memory[61235] <=  8'h00;      memory[61236] <=  8'h00;      memory[61237] <=  8'h00;      memory[61238] <=  8'h00;      memory[61239] <=  8'h00;      memory[61240] <=  8'h00;      memory[61241] <=  8'h00;      memory[61242] <=  8'h00;      memory[61243] <=  8'h00;      memory[61244] <=  8'h00;      memory[61245] <=  8'h00;      memory[61246] <=  8'h00;      memory[61247] <=  8'h00;      memory[61248] <=  8'h00;      memory[61249] <=  8'h00;      memory[61250] <=  8'h00;      memory[61251] <=  8'h00;      memory[61252] <=  8'h00;      memory[61253] <=  8'h00;      memory[61254] <=  8'h00;      memory[61255] <=  8'h00;      memory[61256] <=  8'h00;      memory[61257] <=  8'h00;      memory[61258] <=  8'h00;      memory[61259] <=  8'h00;      memory[61260] <=  8'h00;      memory[61261] <=  8'h00;      memory[61262] <=  8'h00;      memory[61263] <=  8'h00;      memory[61264] <=  8'h00;      memory[61265] <=  8'h00;      memory[61266] <=  8'h00;      memory[61267] <=  8'h00;      memory[61268] <=  8'h00;      memory[61269] <=  8'h00;      memory[61270] <=  8'h00;      memory[61271] <=  8'h00;      memory[61272] <=  8'h00;      memory[61273] <=  8'h00;      memory[61274] <=  8'h00;      memory[61275] <=  8'h00;      memory[61276] <=  8'h00;      memory[61277] <=  8'h00;      memory[61278] <=  8'h00;      memory[61279] <=  8'h00;      memory[61280] <=  8'h00;      memory[61281] <=  8'h00;      memory[61282] <=  8'h00;      memory[61283] <=  8'h00;      memory[61284] <=  8'h00;      memory[61285] <=  8'h00;      memory[61286] <=  8'h00;      memory[61287] <=  8'h00;      memory[61288] <=  8'h00;      memory[61289] <=  8'h00;      memory[61290] <=  8'h00;      memory[61291] <=  8'h00;      memory[61292] <=  8'h00;      memory[61293] <=  8'h00;      memory[61294] <=  8'h00;      memory[61295] <=  8'h00;      memory[61296] <=  8'h00;      memory[61297] <=  8'h00;      memory[61298] <=  8'h00;      memory[61299] <=  8'h00;      memory[61300] <=  8'h00;      memory[61301] <=  8'h00;      memory[61302] <=  8'h00;      memory[61303] <=  8'h00;      memory[61304] <=  8'h00;      memory[61305] <=  8'h00;      memory[61306] <=  8'h00;      memory[61307] <=  8'h00;      memory[61308] <=  8'h00;      memory[61309] <=  8'h00;      memory[61310] <=  8'h00;      memory[61311] <=  8'h00;      memory[61312] <=  8'h00;      memory[61313] <=  8'h00;      memory[61314] <=  8'h00;      memory[61315] <=  8'h00;      memory[61316] <=  8'h00;      memory[61317] <=  8'h00;      memory[61318] <=  8'h00;      memory[61319] <=  8'h00;      memory[61320] <=  8'h00;      memory[61321] <=  8'h00;      memory[61322] <=  8'h00;      memory[61323] <=  8'h00;      memory[61324] <=  8'h00;      memory[61325] <=  8'h00;      memory[61326] <=  8'h00;      memory[61327] <=  8'h00;      memory[61328] <=  8'h00;      memory[61329] <=  8'h00;      memory[61330] <=  8'h00;      memory[61331] <=  8'h00;      memory[61332] <=  8'h00;      memory[61333] <=  8'h00;      memory[61334] <=  8'h00;      memory[61335] <=  8'h00;      memory[61336] <=  8'h00;      memory[61337] <=  8'h00;      memory[61338] <=  8'h00;      memory[61339] <=  8'h00;      memory[61340] <=  8'h00;      memory[61341] <=  8'h00;      memory[61342] <=  8'h00;      memory[61343] <=  8'h00;      memory[61344] <=  8'h00;      memory[61345] <=  8'h00;      memory[61346] <=  8'h00;      memory[61347] <=  8'h00;      memory[61348] <=  8'h00;      memory[61349] <=  8'h00;      memory[61350] <=  8'h00;      memory[61351] <=  8'h00;      memory[61352] <=  8'h00;      memory[61353] <=  8'h00;      memory[61354] <=  8'h00;      memory[61355] <=  8'h00;      memory[61356] <=  8'h00;      memory[61357] <=  8'h00;      memory[61358] <=  8'h00;      memory[61359] <=  8'h00;      memory[61360] <=  8'h00;      memory[61361] <=  8'h00;      memory[61362] <=  8'h00;      memory[61363] <=  8'h00;      memory[61364] <=  8'h00;      memory[61365] <=  8'h00;      memory[61366] <=  8'h00;      memory[61367] <=  8'h00;      memory[61368] <=  8'h00;      memory[61369] <=  8'h00;      memory[61370] <=  8'h00;      memory[61371] <=  8'h00;      memory[61372] <=  8'h00;      memory[61373] <=  8'h00;      memory[61374] <=  8'h00;      memory[61375] <=  8'h00;      memory[61376] <=  8'h00;      memory[61377] <=  8'h00;      memory[61378] <=  8'h00;      memory[61379] <=  8'h00;      memory[61380] <=  8'h00;      memory[61381] <=  8'h00;      memory[61382] <=  8'h00;      memory[61383] <=  8'h00;      memory[61384] <=  8'h00;      memory[61385] <=  8'h00;      memory[61386] <=  8'h00;      memory[61387] <=  8'h00;      memory[61388] <=  8'h00;      memory[61389] <=  8'h00;      memory[61390] <=  8'h00;      memory[61391] <=  8'h00;      memory[61392] <=  8'h00;      memory[61393] <=  8'h00;      memory[61394] <=  8'h00;      memory[61395] <=  8'h00;      memory[61396] <=  8'h00;      memory[61397] <=  8'h00;      memory[61398] <=  8'h00;      memory[61399] <=  8'h00;      memory[61400] <=  8'h00;      memory[61401] <=  8'h00;      memory[61402] <=  8'h00;      memory[61403] <=  8'h00;      memory[61404] <=  8'h00;      memory[61405] <=  8'h00;      memory[61406] <=  8'h00;      memory[61407] <=  8'h00;      memory[61408] <=  8'h00;      memory[61409] <=  8'h00;      memory[61410] <=  8'h00;      memory[61411] <=  8'h00;      memory[61412] <=  8'h00;      memory[61413] <=  8'h00;      memory[61414] <=  8'h00;      memory[61415] <=  8'h00;      memory[61416] <=  8'h00;      memory[61417] <=  8'h00;      memory[61418] <=  8'h00;      memory[61419] <=  8'h00;      memory[61420] <=  8'h00;      memory[61421] <=  8'h00;      memory[61422] <=  8'h00;      memory[61423] <=  8'h00;      memory[61424] <=  8'h00;      memory[61425] <=  8'h00;      memory[61426] <=  8'h00;      memory[61427] <=  8'h00;      memory[61428] <=  8'h00;      memory[61429] <=  8'h00;      memory[61430] <=  8'h00;      memory[61431] <=  8'h00;      memory[61432] <=  8'h00;      memory[61433] <=  8'h00;      memory[61434] <=  8'h00;      memory[61435] <=  8'h00;      memory[61436] <=  8'h00;      memory[61437] <=  8'h00;      memory[61438] <=  8'h00;      memory[61439] <=  8'h00;      memory[61440] <=  8'h00;      memory[61441] <=  8'h00;      memory[61442] <=  8'h00;      memory[61443] <=  8'h00;      memory[61444] <=  8'h00;      memory[61445] <=  8'h00;      memory[61446] <=  8'h00;      memory[61447] <=  8'h00;      memory[61448] <=  8'h00;      memory[61449] <=  8'h00;      memory[61450] <=  8'h00;      memory[61451] <=  8'h00;      memory[61452] <=  8'h00;      memory[61453] <=  8'h00;      memory[61454] <=  8'h00;      memory[61455] <=  8'h00;      memory[61456] <=  8'h00;      memory[61457] <=  8'h00;      memory[61458] <=  8'h00;      memory[61459] <=  8'h00;      memory[61460] <=  8'h00;      memory[61461] <=  8'h00;      memory[61462] <=  8'h00;      memory[61463] <=  8'h00;      memory[61464] <=  8'h00;      memory[61465] <=  8'h00;      memory[61466] <=  8'h00;      memory[61467] <=  8'h00;      memory[61468] <=  8'h00;      memory[61469] <=  8'h00;      memory[61470] <=  8'h00;      memory[61471] <=  8'h00;      memory[61472] <=  8'h00;      memory[61473] <=  8'h00;      memory[61474] <=  8'h00;      memory[61475] <=  8'h00;      memory[61476] <=  8'h00;      memory[61477] <=  8'h00;      memory[61478] <=  8'h00;      memory[61479] <=  8'h00;      memory[61480] <=  8'h00;      memory[61481] <=  8'h00;      memory[61482] <=  8'h00;      memory[61483] <=  8'h00;      memory[61484] <=  8'h00;      memory[61485] <=  8'h00;      memory[61486] <=  8'h00;      memory[61487] <=  8'h00;      memory[61488] <=  8'h00;      memory[61489] <=  8'h00;      memory[61490] <=  8'h00;      memory[61491] <=  8'h00;      memory[61492] <=  8'h00;      memory[61493] <=  8'h00;      memory[61494] <=  8'h00;      memory[61495] <=  8'h00;      memory[61496] <=  8'h00;      memory[61497] <=  8'h00;      memory[61498] <=  8'h00;      memory[61499] <=  8'h00;      memory[61500] <=  8'h00;      memory[61501] <=  8'h00;      memory[61502] <=  8'h00;      memory[61503] <=  8'h00;      memory[61504] <=  8'h00;      memory[61505] <=  8'h00;      memory[61506] <=  8'h00;      memory[61507] <=  8'h00;      memory[61508] <=  8'h00;      memory[61509] <=  8'h00;      memory[61510] <=  8'h00;      memory[61511] <=  8'h00;      memory[61512] <=  8'h00;      memory[61513] <=  8'h00;      memory[61514] <=  8'h00;      memory[61515] <=  8'h00;      memory[61516] <=  8'h00;      memory[61517] <=  8'h00;      memory[61518] <=  8'h00;      memory[61519] <=  8'h00;      memory[61520] <=  8'h00;      memory[61521] <=  8'h00;      memory[61522] <=  8'h00;      memory[61523] <=  8'h00;      memory[61524] <=  8'h00;      memory[61525] <=  8'h00;      memory[61526] <=  8'h00;      memory[61527] <=  8'h00;      memory[61528] <=  8'h00;      memory[61529] <=  8'h00;      memory[61530] <=  8'h00;      memory[61531] <=  8'h00;      memory[61532] <=  8'h00;      memory[61533] <=  8'h00;      memory[61534] <=  8'h00;      memory[61535] <=  8'h00;      memory[61536] <=  8'h00;      memory[61537] <=  8'h00;      memory[61538] <=  8'h00;      memory[61539] <=  8'h00;      memory[61540] <=  8'h00;      memory[61541] <=  8'h00;      memory[61542] <=  8'h00;      memory[61543] <=  8'h00;      memory[61544] <=  8'h00;      memory[61545] <=  8'h00;      memory[61546] <=  8'h00;      memory[61547] <=  8'h00;      memory[61548] <=  8'h00;      memory[61549] <=  8'h00;      memory[61550] <=  8'h00;      memory[61551] <=  8'h00;      memory[61552] <=  8'h00;      memory[61553] <=  8'h00;      memory[61554] <=  8'h00;      memory[61555] <=  8'h00;      memory[61556] <=  8'h00;      memory[61557] <=  8'h00;      memory[61558] <=  8'h00;      memory[61559] <=  8'h00;      memory[61560] <=  8'h00;      memory[61561] <=  8'h00;      memory[61562] <=  8'h00;      memory[61563] <=  8'h00;      memory[61564] <=  8'h00;      memory[61565] <=  8'h00;      memory[61566] <=  8'h00;      memory[61567] <=  8'h00;      memory[61568] <=  8'h00;      memory[61569] <=  8'h00;      memory[61570] <=  8'h00;      memory[61571] <=  8'h00;      memory[61572] <=  8'h00;      memory[61573] <=  8'h00;      memory[61574] <=  8'h00;      memory[61575] <=  8'h00;      memory[61576] <=  8'h00;      memory[61577] <=  8'h00;      memory[61578] <=  8'h00;      memory[61579] <=  8'h00;      memory[61580] <=  8'h00;      memory[61581] <=  8'h00;      memory[61582] <=  8'h00;      memory[61583] <=  8'h00;      memory[61584] <=  8'h00;      memory[61585] <=  8'h00;      memory[61586] <=  8'h00;      memory[61587] <=  8'h00;      memory[61588] <=  8'h00;      memory[61589] <=  8'h00;      memory[61590] <=  8'h00;      memory[61591] <=  8'h00;      memory[61592] <=  8'h00;      memory[61593] <=  8'h00;      memory[61594] <=  8'h00;      memory[61595] <=  8'h00;      memory[61596] <=  8'h00;      memory[61597] <=  8'h00;      memory[61598] <=  8'h00;      memory[61599] <=  8'h00;      memory[61600] <=  8'h00;      memory[61601] <=  8'h00;      memory[61602] <=  8'h00;      memory[61603] <=  8'h00;      memory[61604] <=  8'h00;      memory[61605] <=  8'h00;      memory[61606] <=  8'h00;      memory[61607] <=  8'h00;      memory[61608] <=  8'h00;      memory[61609] <=  8'h00;      memory[61610] <=  8'h00;      memory[61611] <=  8'h00;      memory[61612] <=  8'h00;      memory[61613] <=  8'h00;      memory[61614] <=  8'h00;      memory[61615] <=  8'h00;      memory[61616] <=  8'h00;      memory[61617] <=  8'h00;      memory[61618] <=  8'h00;      memory[61619] <=  8'h00;      memory[61620] <=  8'h00;      memory[61621] <=  8'h00;      memory[61622] <=  8'h00;      memory[61623] <=  8'h00;      memory[61624] <=  8'h00;      memory[61625] <=  8'h00;      memory[61626] <=  8'h00;      memory[61627] <=  8'h00;      memory[61628] <=  8'h00;      memory[61629] <=  8'h00;      memory[61630] <=  8'h00;      memory[61631] <=  8'h00;      memory[61632] <=  8'h00;      memory[61633] <=  8'h00;      memory[61634] <=  8'h00;      memory[61635] <=  8'h00;      memory[61636] <=  8'h00;      memory[61637] <=  8'h00;      memory[61638] <=  8'h00;      memory[61639] <=  8'h00;      memory[61640] <=  8'h00;      memory[61641] <=  8'h00;      memory[61642] <=  8'h00;      memory[61643] <=  8'h00;      memory[61644] <=  8'h00;      memory[61645] <=  8'h00;      memory[61646] <=  8'h00;      memory[61647] <=  8'h00;      memory[61648] <=  8'h00;      memory[61649] <=  8'h00;      memory[61650] <=  8'h00;      memory[61651] <=  8'h00;      memory[61652] <=  8'h00;      memory[61653] <=  8'h00;      memory[61654] <=  8'h00;      memory[61655] <=  8'h00;      memory[61656] <=  8'h00;      memory[61657] <=  8'h00;      memory[61658] <=  8'h00;      memory[61659] <=  8'h00;      memory[61660] <=  8'h00;      memory[61661] <=  8'h00;      memory[61662] <=  8'h00;      memory[61663] <=  8'h00;      memory[61664] <=  8'h00;      memory[61665] <=  8'h00;      memory[61666] <=  8'h00;      memory[61667] <=  8'h00;      memory[61668] <=  8'h00;      memory[61669] <=  8'h00;      memory[61670] <=  8'h00;      memory[61671] <=  8'h00;      memory[61672] <=  8'h00;      memory[61673] <=  8'h00;      memory[61674] <=  8'h00;      memory[61675] <=  8'h00;      memory[61676] <=  8'h00;      memory[61677] <=  8'h00;      memory[61678] <=  8'h00;      memory[61679] <=  8'h00;      memory[61680] <=  8'h00;      memory[61681] <=  8'h00;      memory[61682] <=  8'h00;      memory[61683] <=  8'h00;      memory[61684] <=  8'h00;      memory[61685] <=  8'h00;      memory[61686] <=  8'h00;      memory[61687] <=  8'h00;      memory[61688] <=  8'h00;      memory[61689] <=  8'h00;      memory[61690] <=  8'h00;      memory[61691] <=  8'h00;      memory[61692] <=  8'h00;      memory[61693] <=  8'h00;      memory[61694] <=  8'h00;      memory[61695] <=  8'h00;      memory[61696] <=  8'h00;      memory[61697] <=  8'h00;      memory[61698] <=  8'h00;      memory[61699] <=  8'h00;      memory[61700] <=  8'h00;      memory[61701] <=  8'h00;      memory[61702] <=  8'h00;      memory[61703] <=  8'h00;      memory[61704] <=  8'h00;      memory[61705] <=  8'h00;      memory[61706] <=  8'h00;      memory[61707] <=  8'h00;      memory[61708] <=  8'h00;      memory[61709] <=  8'h00;      memory[61710] <=  8'h00;      memory[61711] <=  8'h00;      memory[61712] <=  8'h00;      memory[61713] <=  8'h00;      memory[61714] <=  8'h00;      memory[61715] <=  8'h00;      memory[61716] <=  8'h00;      memory[61717] <=  8'h00;      memory[61718] <=  8'h00;      memory[61719] <=  8'h00;      memory[61720] <=  8'h00;      memory[61721] <=  8'h00;      memory[61722] <=  8'h00;      memory[61723] <=  8'h00;      memory[61724] <=  8'h00;      memory[61725] <=  8'h00;      memory[61726] <=  8'h00;      memory[61727] <=  8'h00;      memory[61728] <=  8'h00;      memory[61729] <=  8'h00;      memory[61730] <=  8'h00;      memory[61731] <=  8'h00;      memory[61732] <=  8'h00;      memory[61733] <=  8'h00;      memory[61734] <=  8'h00;      memory[61735] <=  8'h00;      memory[61736] <=  8'h00;      memory[61737] <=  8'h00;      memory[61738] <=  8'h00;      memory[61739] <=  8'h00;      memory[61740] <=  8'h00;      memory[61741] <=  8'h00;      memory[61742] <=  8'h00;      memory[61743] <=  8'h00;      memory[61744] <=  8'h00;      memory[61745] <=  8'h00;      memory[61746] <=  8'h00;      memory[61747] <=  8'h00;      memory[61748] <=  8'h00;      memory[61749] <=  8'h00;      memory[61750] <=  8'h00;      memory[61751] <=  8'h00;      memory[61752] <=  8'h00;      memory[61753] <=  8'h00;      memory[61754] <=  8'h00;      memory[61755] <=  8'h00;      memory[61756] <=  8'h00;      memory[61757] <=  8'h00;      memory[61758] <=  8'h00;      memory[61759] <=  8'h00;      memory[61760] <=  8'h00;      memory[61761] <=  8'h00;      memory[61762] <=  8'h00;      memory[61763] <=  8'h00;      memory[61764] <=  8'h00;      memory[61765] <=  8'h00;      memory[61766] <=  8'h00;      memory[61767] <=  8'h00;      memory[61768] <=  8'h00;      memory[61769] <=  8'h00;      memory[61770] <=  8'h00;      memory[61771] <=  8'h00;      memory[61772] <=  8'h00;      memory[61773] <=  8'h00;      memory[61774] <=  8'h00;      memory[61775] <=  8'h00;      memory[61776] <=  8'h00;      memory[61777] <=  8'h00;      memory[61778] <=  8'h00;      memory[61779] <=  8'h00;      memory[61780] <=  8'h00;      memory[61781] <=  8'h00;      memory[61782] <=  8'h00;      memory[61783] <=  8'h00;      memory[61784] <=  8'h00;      memory[61785] <=  8'h00;      memory[61786] <=  8'h00;      memory[61787] <=  8'h00;      memory[61788] <=  8'h00;      memory[61789] <=  8'h00;      memory[61790] <=  8'h00;      memory[61791] <=  8'h00;      memory[61792] <=  8'h00;      memory[61793] <=  8'h00;      memory[61794] <=  8'h00;      memory[61795] <=  8'h00;      memory[61796] <=  8'h00;      memory[61797] <=  8'h00;      memory[61798] <=  8'h00;      memory[61799] <=  8'h00;      memory[61800] <=  8'h00;      memory[61801] <=  8'h00;      memory[61802] <=  8'h00;      memory[61803] <=  8'h00;      memory[61804] <=  8'h00;      memory[61805] <=  8'h00;      memory[61806] <=  8'h00;      memory[61807] <=  8'h00;      memory[61808] <=  8'h00;      memory[61809] <=  8'h00;      memory[61810] <=  8'h00;      memory[61811] <=  8'h00;      memory[61812] <=  8'h00;      memory[61813] <=  8'h00;      memory[61814] <=  8'h00;      memory[61815] <=  8'h00;      memory[61816] <=  8'h00;      memory[61817] <=  8'h00;      memory[61818] <=  8'h00;      memory[61819] <=  8'h00;      memory[61820] <=  8'h00;      memory[61821] <=  8'h00;      memory[61822] <=  8'h00;      memory[61823] <=  8'h00;      memory[61824] <=  8'h00;      memory[61825] <=  8'h00;      memory[61826] <=  8'h00;      memory[61827] <=  8'h00;      memory[61828] <=  8'h00;      memory[61829] <=  8'h00;      memory[61830] <=  8'h00;      memory[61831] <=  8'h00;      memory[61832] <=  8'h00;      memory[61833] <=  8'h00;      memory[61834] <=  8'h00;      memory[61835] <=  8'h00;      memory[61836] <=  8'h00;      memory[61837] <=  8'h00;      memory[61838] <=  8'h00;      memory[61839] <=  8'h00;      memory[61840] <=  8'h00;      memory[61841] <=  8'h00;      memory[61842] <=  8'h00;      memory[61843] <=  8'h00;      memory[61844] <=  8'h00;      memory[61845] <=  8'h00;      memory[61846] <=  8'h00;      memory[61847] <=  8'h00;      memory[61848] <=  8'h00;      memory[61849] <=  8'h00;      memory[61850] <=  8'h00;      memory[61851] <=  8'h00;      memory[61852] <=  8'h00;      memory[61853] <=  8'h00;      memory[61854] <=  8'h00;      memory[61855] <=  8'h00;      memory[61856] <=  8'h00;      memory[61857] <=  8'h00;      memory[61858] <=  8'h00;      memory[61859] <=  8'h00;      memory[61860] <=  8'h00;      memory[61861] <=  8'h00;      memory[61862] <=  8'h00;      memory[61863] <=  8'h00;      memory[61864] <=  8'h00;      memory[61865] <=  8'h00;      memory[61866] <=  8'h00;      memory[61867] <=  8'h00;      memory[61868] <=  8'h00;      memory[61869] <=  8'h00;      memory[61870] <=  8'h00;      memory[61871] <=  8'h00;      memory[61872] <=  8'h00;      memory[61873] <=  8'h00;      memory[61874] <=  8'h00;      memory[61875] <=  8'h00;      memory[61876] <=  8'h00;      memory[61877] <=  8'h00;      memory[61878] <=  8'h00;      memory[61879] <=  8'h00;      memory[61880] <=  8'h00;      memory[61881] <=  8'h00;      memory[61882] <=  8'h00;      memory[61883] <=  8'h00;      memory[61884] <=  8'h00;      memory[61885] <=  8'h00;      memory[61886] <=  8'h00;      memory[61887] <=  8'h00;      memory[61888] <=  8'h00;      memory[61889] <=  8'h00;      memory[61890] <=  8'h00;      memory[61891] <=  8'h00;      memory[61892] <=  8'h00;      memory[61893] <=  8'h00;      memory[61894] <=  8'h00;      memory[61895] <=  8'h00;      memory[61896] <=  8'h00;      memory[61897] <=  8'h00;      memory[61898] <=  8'h00;      memory[61899] <=  8'h00;      memory[61900] <=  8'h00;      memory[61901] <=  8'h00;      memory[61902] <=  8'h00;      memory[61903] <=  8'h00;      memory[61904] <=  8'h00;      memory[61905] <=  8'h00;      memory[61906] <=  8'h00;      memory[61907] <=  8'h00;      memory[61908] <=  8'h00;      memory[61909] <=  8'h00;      memory[61910] <=  8'h00;      memory[61911] <=  8'h00;      memory[61912] <=  8'h00;      memory[61913] <=  8'h00;      memory[61914] <=  8'h00;      memory[61915] <=  8'h00;      memory[61916] <=  8'h00;      memory[61917] <=  8'h00;      memory[61918] <=  8'h00;      memory[61919] <=  8'h00;      memory[61920] <=  8'h00;      memory[61921] <=  8'h00;      memory[61922] <=  8'h00;      memory[61923] <=  8'h00;      memory[61924] <=  8'h00;      memory[61925] <=  8'h00;      memory[61926] <=  8'h00;      memory[61927] <=  8'h00;      memory[61928] <=  8'h00;      memory[61929] <=  8'h00;      memory[61930] <=  8'h00;      memory[61931] <=  8'h00;      memory[61932] <=  8'h00;      memory[61933] <=  8'h00;      memory[61934] <=  8'h00;      memory[61935] <=  8'h00;      memory[61936] <=  8'h00;      memory[61937] <=  8'h00;      memory[61938] <=  8'h00;      memory[61939] <=  8'h00;      memory[61940] <=  8'h00;      memory[61941] <=  8'h00;      memory[61942] <=  8'h00;      memory[61943] <=  8'h00;      memory[61944] <=  8'h00;      memory[61945] <=  8'h00;      memory[61946] <=  8'h00;      memory[61947] <=  8'h00;      memory[61948] <=  8'h00;      memory[61949] <=  8'h00;      memory[61950] <=  8'h00;      memory[61951] <=  8'h00;      memory[61952] <=  8'h00;      memory[61953] <=  8'h00;      memory[61954] <=  8'h00;      memory[61955] <=  8'h00;      memory[61956] <=  8'h00;      memory[61957] <=  8'h00;      memory[61958] <=  8'h00;      memory[61959] <=  8'h00;      memory[61960] <=  8'h00;      memory[61961] <=  8'h00;      memory[61962] <=  8'h00;      memory[61963] <=  8'h00;      memory[61964] <=  8'h00;      memory[61965] <=  8'h00;      memory[61966] <=  8'h00;      memory[61967] <=  8'h00;      memory[61968] <=  8'h00;      memory[61969] <=  8'h00;      memory[61970] <=  8'h00;      memory[61971] <=  8'h00;      memory[61972] <=  8'h00;      memory[61973] <=  8'h00;      memory[61974] <=  8'h00;      memory[61975] <=  8'h00;      memory[61976] <=  8'h00;      memory[61977] <=  8'h00;      memory[61978] <=  8'h00;      memory[61979] <=  8'h00;      memory[61980] <=  8'h00;      memory[61981] <=  8'h00;      memory[61982] <=  8'h00;      memory[61983] <=  8'h00;      memory[61984] <=  8'h00;      memory[61985] <=  8'h00;      memory[61986] <=  8'h00;      memory[61987] <=  8'h00;      memory[61988] <=  8'h00;      memory[61989] <=  8'h00;      memory[61990] <=  8'h00;      memory[61991] <=  8'h00;      memory[61992] <=  8'h00;      memory[61993] <=  8'h00;      memory[61994] <=  8'h00;      memory[61995] <=  8'h00;      memory[61996] <=  8'h00;      memory[61997] <=  8'h00;      memory[61998] <=  8'h00;      memory[61999] <=  8'h00;      memory[62000] <=  8'h00;      memory[62001] <=  8'h00;      memory[62002] <=  8'h00;      memory[62003] <=  8'h00;      memory[62004] <=  8'h00;      memory[62005] <=  8'h00;      memory[62006] <=  8'h00;      memory[62007] <=  8'h00;      memory[62008] <=  8'h00;      memory[62009] <=  8'h00;      memory[62010] <=  8'h00;      memory[62011] <=  8'h00;      memory[62012] <=  8'h00;      memory[62013] <=  8'h00;      memory[62014] <=  8'h00;      memory[62015] <=  8'h00;      memory[62016] <=  8'h00;      memory[62017] <=  8'h00;      memory[62018] <=  8'h00;      memory[62019] <=  8'h00;      memory[62020] <=  8'h00;      memory[62021] <=  8'h00;      memory[62022] <=  8'h00;      memory[62023] <=  8'h00;      memory[62024] <=  8'h00;      memory[62025] <=  8'h00;      memory[62026] <=  8'h00;      memory[62027] <=  8'h00;      memory[62028] <=  8'h00;      memory[62029] <=  8'h00;      memory[62030] <=  8'h00;      memory[62031] <=  8'h00;      memory[62032] <=  8'h00;      memory[62033] <=  8'h00;      memory[62034] <=  8'h00;      memory[62035] <=  8'h00;      memory[62036] <=  8'h00;      memory[62037] <=  8'h00;      memory[62038] <=  8'h00;      memory[62039] <=  8'h00;      memory[62040] <=  8'h00;      memory[62041] <=  8'h00;      memory[62042] <=  8'h00;      memory[62043] <=  8'h00;      memory[62044] <=  8'h00;      memory[62045] <=  8'h00;      memory[62046] <=  8'h00;      memory[62047] <=  8'h00;      memory[62048] <=  8'h00;      memory[62049] <=  8'h00;      memory[62050] <=  8'h00;      memory[62051] <=  8'h00;      memory[62052] <=  8'h00;      memory[62053] <=  8'h00;      memory[62054] <=  8'h00;      memory[62055] <=  8'h00;      memory[62056] <=  8'h00;      memory[62057] <=  8'h00;      memory[62058] <=  8'h00;      memory[62059] <=  8'h00;      memory[62060] <=  8'h00;      memory[62061] <=  8'h00;      memory[62062] <=  8'h00;      memory[62063] <=  8'h00;      memory[62064] <=  8'h00;      memory[62065] <=  8'h00;      memory[62066] <=  8'h00;      memory[62067] <=  8'h00;      memory[62068] <=  8'h00;      memory[62069] <=  8'h00;      memory[62070] <=  8'h00;      memory[62071] <=  8'h00;      memory[62072] <=  8'h00;      memory[62073] <=  8'h00;      memory[62074] <=  8'h00;      memory[62075] <=  8'h00;      memory[62076] <=  8'h00;      memory[62077] <=  8'h00;      memory[62078] <=  8'h00;      memory[62079] <=  8'h00;      memory[62080] <=  8'h00;      memory[62081] <=  8'h00;      memory[62082] <=  8'h00;      memory[62083] <=  8'h00;      memory[62084] <=  8'h00;      memory[62085] <=  8'h00;      memory[62086] <=  8'h00;      memory[62087] <=  8'h00;      memory[62088] <=  8'h00;      memory[62089] <=  8'h00;      memory[62090] <=  8'h00;      memory[62091] <=  8'h00;      memory[62092] <=  8'h00;      memory[62093] <=  8'h00;      memory[62094] <=  8'h00;      memory[62095] <=  8'h00;      memory[62096] <=  8'h00;      memory[62097] <=  8'h00;      memory[62098] <=  8'h00;      memory[62099] <=  8'h00;      memory[62100] <=  8'h00;      memory[62101] <=  8'h00;      memory[62102] <=  8'h00;      memory[62103] <=  8'h00;      memory[62104] <=  8'h00;      memory[62105] <=  8'h00;      memory[62106] <=  8'h00;      memory[62107] <=  8'h00;      memory[62108] <=  8'h00;      memory[62109] <=  8'h00;      memory[62110] <=  8'h00;      memory[62111] <=  8'h00;      memory[62112] <=  8'h00;      memory[62113] <=  8'h00;      memory[62114] <=  8'h00;      memory[62115] <=  8'h00;      memory[62116] <=  8'h00;      memory[62117] <=  8'h00;      memory[62118] <=  8'h00;      memory[62119] <=  8'h00;      memory[62120] <=  8'h00;      memory[62121] <=  8'h00;      memory[62122] <=  8'h00;      memory[62123] <=  8'h00;      memory[62124] <=  8'h00;      memory[62125] <=  8'h00;      memory[62126] <=  8'h00;      memory[62127] <=  8'h00;      memory[62128] <=  8'h00;      memory[62129] <=  8'h00;      memory[62130] <=  8'h00;      memory[62131] <=  8'h00;      memory[62132] <=  8'h00;      memory[62133] <=  8'h00;      memory[62134] <=  8'h00;      memory[62135] <=  8'h00;      memory[62136] <=  8'h00;      memory[62137] <=  8'h00;      memory[62138] <=  8'h00;      memory[62139] <=  8'h00;      memory[62140] <=  8'h00;      memory[62141] <=  8'h00;      memory[62142] <=  8'h00;      memory[62143] <=  8'h00;      memory[62144] <=  8'h00;      memory[62145] <=  8'h00;      memory[62146] <=  8'h00;      memory[62147] <=  8'h00;      memory[62148] <=  8'h00;      memory[62149] <=  8'h00;      memory[62150] <=  8'h00;      memory[62151] <=  8'h00;      memory[62152] <=  8'h00;      memory[62153] <=  8'h00;      memory[62154] <=  8'h00;      memory[62155] <=  8'h00;      memory[62156] <=  8'h00;      memory[62157] <=  8'h00;      memory[62158] <=  8'h00;      memory[62159] <=  8'h00;      memory[62160] <=  8'h00;      memory[62161] <=  8'h00;      memory[62162] <=  8'h00;      memory[62163] <=  8'h00;      memory[62164] <=  8'h00;      memory[62165] <=  8'h00;      memory[62166] <=  8'h00;      memory[62167] <=  8'h00;      memory[62168] <=  8'h00;      memory[62169] <=  8'h00;      memory[62170] <=  8'h00;      memory[62171] <=  8'h00;      memory[62172] <=  8'h00;      memory[62173] <=  8'h00;      memory[62174] <=  8'h00;      memory[62175] <=  8'h00;      memory[62176] <=  8'h00;      memory[62177] <=  8'h00;      memory[62178] <=  8'h00;      memory[62179] <=  8'h00;      memory[62180] <=  8'h00;      memory[62181] <=  8'h00;      memory[62182] <=  8'h00;      memory[62183] <=  8'h00;      memory[62184] <=  8'h00;      memory[62185] <=  8'h00;      memory[62186] <=  8'h00;      memory[62187] <=  8'h00;      memory[62188] <=  8'h00;      memory[62189] <=  8'h00;      memory[62190] <=  8'h00;      memory[62191] <=  8'h00;      memory[62192] <=  8'h00;      memory[62193] <=  8'h00;      memory[62194] <=  8'h00;      memory[62195] <=  8'h00;      memory[62196] <=  8'h00;      memory[62197] <=  8'h00;      memory[62198] <=  8'h00;      memory[62199] <=  8'h00;      memory[62200] <=  8'h00;      memory[62201] <=  8'h00;      memory[62202] <=  8'h00;      memory[62203] <=  8'h00;      memory[62204] <=  8'h00;      memory[62205] <=  8'h00;      memory[62206] <=  8'h00;      memory[62207] <=  8'h00;      memory[62208] <=  8'h00;      memory[62209] <=  8'h00;      memory[62210] <=  8'h00;      memory[62211] <=  8'h00;      memory[62212] <=  8'h00;      memory[62213] <=  8'h00;      memory[62214] <=  8'h00;      memory[62215] <=  8'h00;      memory[62216] <=  8'h00;      memory[62217] <=  8'h00;      memory[62218] <=  8'h00;      memory[62219] <=  8'h00;      memory[62220] <=  8'h00;      memory[62221] <=  8'h00;      memory[62222] <=  8'h00;      memory[62223] <=  8'h00;      memory[62224] <=  8'h00;      memory[62225] <=  8'h00;      memory[62226] <=  8'h00;      memory[62227] <=  8'h00;      memory[62228] <=  8'h00;      memory[62229] <=  8'h00;      memory[62230] <=  8'h00;      memory[62231] <=  8'h00;      memory[62232] <=  8'h00;      memory[62233] <=  8'h00;      memory[62234] <=  8'h00;      memory[62235] <=  8'h00;      memory[62236] <=  8'h00;      memory[62237] <=  8'h00;      memory[62238] <=  8'h00;      memory[62239] <=  8'h00;      memory[62240] <=  8'h00;      memory[62241] <=  8'h00;      memory[62242] <=  8'h00;      memory[62243] <=  8'h00;      memory[62244] <=  8'h00;      memory[62245] <=  8'h00;      memory[62246] <=  8'h00;      memory[62247] <=  8'h00;      memory[62248] <=  8'h00;      memory[62249] <=  8'h00;      memory[62250] <=  8'h00;      memory[62251] <=  8'h00;      memory[62252] <=  8'h00;      memory[62253] <=  8'h00;      memory[62254] <=  8'h00;      memory[62255] <=  8'h00;      memory[62256] <=  8'h00;      memory[62257] <=  8'h00;      memory[62258] <=  8'h00;      memory[62259] <=  8'h00;      memory[62260] <=  8'h00;      memory[62261] <=  8'h00;      memory[62262] <=  8'h00;      memory[62263] <=  8'h00;      memory[62264] <=  8'h00;      memory[62265] <=  8'h00;      memory[62266] <=  8'h00;      memory[62267] <=  8'h00;      memory[62268] <=  8'h00;      memory[62269] <=  8'h00;      memory[62270] <=  8'h00;      memory[62271] <=  8'h00;      memory[62272] <=  8'h00;      memory[62273] <=  8'h00;      memory[62274] <=  8'h00;      memory[62275] <=  8'h00;      memory[62276] <=  8'h00;      memory[62277] <=  8'h00;      memory[62278] <=  8'h00;      memory[62279] <=  8'h00;      memory[62280] <=  8'h00;      memory[62281] <=  8'h00;      memory[62282] <=  8'h00;      memory[62283] <=  8'h00;      memory[62284] <=  8'h00;      memory[62285] <=  8'h00;      memory[62286] <=  8'h00;      memory[62287] <=  8'h00;      memory[62288] <=  8'h00;      memory[62289] <=  8'h00;      memory[62290] <=  8'h00;      memory[62291] <=  8'h00;      memory[62292] <=  8'h00;      memory[62293] <=  8'h00;      memory[62294] <=  8'h00;      memory[62295] <=  8'h00;      memory[62296] <=  8'h00;      memory[62297] <=  8'h00;      memory[62298] <=  8'h00;      memory[62299] <=  8'h00;      memory[62300] <=  8'h00;      memory[62301] <=  8'h00;      memory[62302] <=  8'h00;      memory[62303] <=  8'h00;      memory[62304] <=  8'h00;      memory[62305] <=  8'h00;      memory[62306] <=  8'h00;      memory[62307] <=  8'h00;      memory[62308] <=  8'h00;      memory[62309] <=  8'h00;      memory[62310] <=  8'h00;      memory[62311] <=  8'h00;      memory[62312] <=  8'h00;      memory[62313] <=  8'h00;      memory[62314] <=  8'h00;      memory[62315] <=  8'h00;      memory[62316] <=  8'h00;      memory[62317] <=  8'h00;      memory[62318] <=  8'h00;      memory[62319] <=  8'h00;      memory[62320] <=  8'h00;      memory[62321] <=  8'h00;      memory[62322] <=  8'h00;      memory[62323] <=  8'h00;      memory[62324] <=  8'h00;      memory[62325] <=  8'h00;      memory[62326] <=  8'h00;      memory[62327] <=  8'h00;      memory[62328] <=  8'h00;      memory[62329] <=  8'h00;      memory[62330] <=  8'h00;      memory[62331] <=  8'h00;      memory[62332] <=  8'h00;      memory[62333] <=  8'h00;      memory[62334] <=  8'h00;      memory[62335] <=  8'h00;      memory[62336] <=  8'h00;      memory[62337] <=  8'h00;      memory[62338] <=  8'h00;      memory[62339] <=  8'h00;      memory[62340] <=  8'h00;      memory[62341] <=  8'h00;      memory[62342] <=  8'h00;      memory[62343] <=  8'h00;      memory[62344] <=  8'h00;      memory[62345] <=  8'h00;      memory[62346] <=  8'h00;      memory[62347] <=  8'h00;      memory[62348] <=  8'h00;      memory[62349] <=  8'h00;      memory[62350] <=  8'h00;      memory[62351] <=  8'h00;      memory[62352] <=  8'h00;      memory[62353] <=  8'h00;      memory[62354] <=  8'h00;      memory[62355] <=  8'h00;      memory[62356] <=  8'h00;      memory[62357] <=  8'h00;      memory[62358] <=  8'h00;      memory[62359] <=  8'h00;      memory[62360] <=  8'h00;      memory[62361] <=  8'h00;      memory[62362] <=  8'h00;      memory[62363] <=  8'h00;      memory[62364] <=  8'h00;      memory[62365] <=  8'h00;      memory[62366] <=  8'h00;      memory[62367] <=  8'h00;      memory[62368] <=  8'h00;      memory[62369] <=  8'h00;      memory[62370] <=  8'h00;      memory[62371] <=  8'h00;      memory[62372] <=  8'h00;      memory[62373] <=  8'h00;      memory[62374] <=  8'h00;      memory[62375] <=  8'h00;      memory[62376] <=  8'h00;      memory[62377] <=  8'h00;      memory[62378] <=  8'h00;      memory[62379] <=  8'h00;      memory[62380] <=  8'h00;      memory[62381] <=  8'h00;      memory[62382] <=  8'h00;      memory[62383] <=  8'h00;      memory[62384] <=  8'h00;      memory[62385] <=  8'h00;      memory[62386] <=  8'h00;      memory[62387] <=  8'h00;      memory[62388] <=  8'h00;      memory[62389] <=  8'h00;      memory[62390] <=  8'h00;      memory[62391] <=  8'h00;      memory[62392] <=  8'h00;      memory[62393] <=  8'h00;      memory[62394] <=  8'h00;      memory[62395] <=  8'h00;      memory[62396] <=  8'h00;      memory[62397] <=  8'h00;      memory[62398] <=  8'h00;      memory[62399] <=  8'h00;      memory[62400] <=  8'h00;      memory[62401] <=  8'h00;      memory[62402] <=  8'h00;      memory[62403] <=  8'h00;      memory[62404] <=  8'h00;      memory[62405] <=  8'h00;      memory[62406] <=  8'h00;      memory[62407] <=  8'h00;      memory[62408] <=  8'h00;      memory[62409] <=  8'h00;      memory[62410] <=  8'h00;      memory[62411] <=  8'h00;      memory[62412] <=  8'h00;      memory[62413] <=  8'h00;      memory[62414] <=  8'h00;      memory[62415] <=  8'h00;      memory[62416] <=  8'h00;      memory[62417] <=  8'h00;      memory[62418] <=  8'h00;      memory[62419] <=  8'h00;      memory[62420] <=  8'h00;      memory[62421] <=  8'h00;      memory[62422] <=  8'h00;      memory[62423] <=  8'h00;      memory[62424] <=  8'h00;      memory[62425] <=  8'h00;      memory[62426] <=  8'h00;      memory[62427] <=  8'h00;      memory[62428] <=  8'h00;      memory[62429] <=  8'h00;      memory[62430] <=  8'h00;      memory[62431] <=  8'h00;      memory[62432] <=  8'h00;      memory[62433] <=  8'h00;      memory[62434] <=  8'h00;      memory[62435] <=  8'h00;      memory[62436] <=  8'h00;      memory[62437] <=  8'h00;      memory[62438] <=  8'h00;      memory[62439] <=  8'h00;      memory[62440] <=  8'h00;      memory[62441] <=  8'h00;      memory[62442] <=  8'h00;      memory[62443] <=  8'h00;      memory[62444] <=  8'h00;      memory[62445] <=  8'h00;      memory[62446] <=  8'h00;      memory[62447] <=  8'h00;      memory[62448] <=  8'h00;      memory[62449] <=  8'h00;      memory[62450] <=  8'h00;      memory[62451] <=  8'h00;      memory[62452] <=  8'h00;      memory[62453] <=  8'h00;      memory[62454] <=  8'h00;      memory[62455] <=  8'h00;      memory[62456] <=  8'h00;      memory[62457] <=  8'h00;      memory[62458] <=  8'h00;      memory[62459] <=  8'h00;      memory[62460] <=  8'h00;      memory[62461] <=  8'h00;      memory[62462] <=  8'h00;      memory[62463] <=  8'h00;      memory[62464] <=  8'h00;      memory[62465] <=  8'h00;      memory[62466] <=  8'h00;      memory[62467] <=  8'h00;      memory[62468] <=  8'h00;      memory[62469] <=  8'h00;      memory[62470] <=  8'h00;      memory[62471] <=  8'h00;      memory[62472] <=  8'h00;      memory[62473] <=  8'h00;      memory[62474] <=  8'h00;      memory[62475] <=  8'h00;      memory[62476] <=  8'h00;      memory[62477] <=  8'h00;      memory[62478] <=  8'h00;      memory[62479] <=  8'h00;      memory[62480] <=  8'h00;      memory[62481] <=  8'h00;      memory[62482] <=  8'h00;      memory[62483] <=  8'h00;      memory[62484] <=  8'h00;      memory[62485] <=  8'h00;      memory[62486] <=  8'h00;      memory[62487] <=  8'h00;      memory[62488] <=  8'h00;      memory[62489] <=  8'h00;      memory[62490] <=  8'h00;      memory[62491] <=  8'h00;      memory[62492] <=  8'h00;      memory[62493] <=  8'h00;      memory[62494] <=  8'h00;      memory[62495] <=  8'h00;      memory[62496] <=  8'h00;      memory[62497] <=  8'h00;      memory[62498] <=  8'h00;      memory[62499] <=  8'h00;      memory[62500] <=  8'h00;      memory[62501] <=  8'h00;      memory[62502] <=  8'h00;      memory[62503] <=  8'h00;      memory[62504] <=  8'h00;      memory[62505] <=  8'h00;      memory[62506] <=  8'h00;      memory[62507] <=  8'h00;      memory[62508] <=  8'h00;      memory[62509] <=  8'h00;      memory[62510] <=  8'h00;      memory[62511] <=  8'h00;      memory[62512] <=  8'h00;      memory[62513] <=  8'h00;      memory[62514] <=  8'h00;      memory[62515] <=  8'h00;      memory[62516] <=  8'h00;      memory[62517] <=  8'h00;      memory[62518] <=  8'h00;      memory[62519] <=  8'h00;      memory[62520] <=  8'h00;      memory[62521] <=  8'h00;      memory[62522] <=  8'h00;      memory[62523] <=  8'h00;      memory[62524] <=  8'h00;      memory[62525] <=  8'h00;      memory[62526] <=  8'h00;      memory[62527] <=  8'h00;      memory[62528] <=  8'h00;      memory[62529] <=  8'h00;      memory[62530] <=  8'h00;      memory[62531] <=  8'h00;      memory[62532] <=  8'h00;      memory[62533] <=  8'h00;      memory[62534] <=  8'h00;      memory[62535] <=  8'h00;      memory[62536] <=  8'h00;      memory[62537] <=  8'h00;      memory[62538] <=  8'h00;      memory[62539] <=  8'h00;      memory[62540] <=  8'h00;      memory[62541] <=  8'h00;      memory[62542] <=  8'h00;      memory[62543] <=  8'h00;      memory[62544] <=  8'h00;      memory[62545] <=  8'h00;      memory[62546] <=  8'h00;      memory[62547] <=  8'h00;      memory[62548] <=  8'h00;      memory[62549] <=  8'h00;      memory[62550] <=  8'h00;      memory[62551] <=  8'h00;      memory[62552] <=  8'h00;      memory[62553] <=  8'h00;      memory[62554] <=  8'h00;      memory[62555] <=  8'h00;      memory[62556] <=  8'h00;      memory[62557] <=  8'h00;      memory[62558] <=  8'h00;      memory[62559] <=  8'h00;      memory[62560] <=  8'h00;      memory[62561] <=  8'h00;      memory[62562] <=  8'h00;      memory[62563] <=  8'h00;      memory[62564] <=  8'h00;      memory[62565] <=  8'h00;      memory[62566] <=  8'h00;      memory[62567] <=  8'h00;      memory[62568] <=  8'h00;      memory[62569] <=  8'h00;      memory[62570] <=  8'h00;      memory[62571] <=  8'h00;      memory[62572] <=  8'h00;      memory[62573] <=  8'h00;      memory[62574] <=  8'h00;      memory[62575] <=  8'h00;      memory[62576] <=  8'h00;      memory[62577] <=  8'h00;      memory[62578] <=  8'h00;      memory[62579] <=  8'h00;      memory[62580] <=  8'h00;      memory[62581] <=  8'h00;      memory[62582] <=  8'h00;      memory[62583] <=  8'h00;      memory[62584] <=  8'h00;      memory[62585] <=  8'h00;      memory[62586] <=  8'h00;      memory[62587] <=  8'h00;      memory[62588] <=  8'h00;      memory[62589] <=  8'h00;      memory[62590] <=  8'h00;      memory[62591] <=  8'h00;      memory[62592] <=  8'h00;      memory[62593] <=  8'h00;      memory[62594] <=  8'h00;      memory[62595] <=  8'h00;      memory[62596] <=  8'h00;      memory[62597] <=  8'h00;      memory[62598] <=  8'h00;      memory[62599] <=  8'h00;      memory[62600] <=  8'h00;      memory[62601] <=  8'h00;      memory[62602] <=  8'h00;      memory[62603] <=  8'h00;      memory[62604] <=  8'h00;      memory[62605] <=  8'h00;      memory[62606] <=  8'h00;      memory[62607] <=  8'h00;      memory[62608] <=  8'h00;      memory[62609] <=  8'h00;      memory[62610] <=  8'h00;      memory[62611] <=  8'h00;      memory[62612] <=  8'h00;      memory[62613] <=  8'h00;      memory[62614] <=  8'h00;      memory[62615] <=  8'h00;      memory[62616] <=  8'h00;      memory[62617] <=  8'h00;      memory[62618] <=  8'h00;      memory[62619] <=  8'h00;      memory[62620] <=  8'h00;      memory[62621] <=  8'h00;      memory[62622] <=  8'h00;      memory[62623] <=  8'h00;      memory[62624] <=  8'h00;      memory[62625] <=  8'h00;      memory[62626] <=  8'h00;      memory[62627] <=  8'h00;      memory[62628] <=  8'h00;      memory[62629] <=  8'h00;      memory[62630] <=  8'h00;      memory[62631] <=  8'h00;      memory[62632] <=  8'h00;      memory[62633] <=  8'h00;      memory[62634] <=  8'h00;      memory[62635] <=  8'h00;      memory[62636] <=  8'h00;      memory[62637] <=  8'h00;      memory[62638] <=  8'h00;      memory[62639] <=  8'h00;      memory[62640] <=  8'h00;      memory[62641] <=  8'h00;      memory[62642] <=  8'h00;      memory[62643] <=  8'h00;      memory[62644] <=  8'h00;      memory[62645] <=  8'h00;      memory[62646] <=  8'h00;      memory[62647] <=  8'h00;      memory[62648] <=  8'h00;      memory[62649] <=  8'h00;      memory[62650] <=  8'h00;      memory[62651] <=  8'h00;      memory[62652] <=  8'h00;      memory[62653] <=  8'h00;      memory[62654] <=  8'h00;      memory[62655] <=  8'h00;      memory[62656] <=  8'h00;      memory[62657] <=  8'h00;      memory[62658] <=  8'h00;      memory[62659] <=  8'h00;      memory[62660] <=  8'h00;      memory[62661] <=  8'h00;      memory[62662] <=  8'h00;      memory[62663] <=  8'h00;      memory[62664] <=  8'h00;      memory[62665] <=  8'h00;      memory[62666] <=  8'h00;      memory[62667] <=  8'h00;      memory[62668] <=  8'h00;      memory[62669] <=  8'h00;      memory[62670] <=  8'h00;      memory[62671] <=  8'h00;      memory[62672] <=  8'h00;      memory[62673] <=  8'h00;      memory[62674] <=  8'h00;      memory[62675] <=  8'h00;      memory[62676] <=  8'h00;      memory[62677] <=  8'h00;      memory[62678] <=  8'h00;      memory[62679] <=  8'h00;      memory[62680] <=  8'h00;      memory[62681] <=  8'h00;      memory[62682] <=  8'h00;      memory[62683] <=  8'h00;      memory[62684] <=  8'h00;      memory[62685] <=  8'h00;      memory[62686] <=  8'h00;      memory[62687] <=  8'h00;      memory[62688] <=  8'h00;      memory[62689] <=  8'h00;      memory[62690] <=  8'h00;      memory[62691] <=  8'h00;      memory[62692] <=  8'h00;      memory[62693] <=  8'h00;      memory[62694] <=  8'h00;      memory[62695] <=  8'h00;      memory[62696] <=  8'h00;      memory[62697] <=  8'h00;      memory[62698] <=  8'h00;      memory[62699] <=  8'h00;      memory[62700] <=  8'h00;      memory[62701] <=  8'h00;      memory[62702] <=  8'h00;      memory[62703] <=  8'h00;      memory[62704] <=  8'h00;      memory[62705] <=  8'h00;      memory[62706] <=  8'h00;      memory[62707] <=  8'h00;      memory[62708] <=  8'h00;      memory[62709] <=  8'h00;      memory[62710] <=  8'h00;      memory[62711] <=  8'h00;      memory[62712] <=  8'h00;      memory[62713] <=  8'h00;      memory[62714] <=  8'h00;      memory[62715] <=  8'h00;      memory[62716] <=  8'h00;      memory[62717] <=  8'h00;      memory[62718] <=  8'h00;      memory[62719] <=  8'h00;      memory[62720] <=  8'h00;      memory[62721] <=  8'h00;      memory[62722] <=  8'h00;      memory[62723] <=  8'h00;      memory[62724] <=  8'h00;      memory[62725] <=  8'h00;      memory[62726] <=  8'h00;      memory[62727] <=  8'h00;      memory[62728] <=  8'h00;      memory[62729] <=  8'h00;      memory[62730] <=  8'h00;      memory[62731] <=  8'h00;      memory[62732] <=  8'h00;      memory[62733] <=  8'h00;      memory[62734] <=  8'h00;      memory[62735] <=  8'h00;      memory[62736] <=  8'h00;      memory[62737] <=  8'h00;      memory[62738] <=  8'h00;      memory[62739] <=  8'h00;      memory[62740] <=  8'h00;      memory[62741] <=  8'h00;      memory[62742] <=  8'h00;      memory[62743] <=  8'h00;      memory[62744] <=  8'h00;      memory[62745] <=  8'h00;      memory[62746] <=  8'h00;      memory[62747] <=  8'h00;      memory[62748] <=  8'h00;      memory[62749] <=  8'h00;      memory[62750] <=  8'h00;      memory[62751] <=  8'h00;      memory[62752] <=  8'h00;      memory[62753] <=  8'h00;      memory[62754] <=  8'h00;      memory[62755] <=  8'h00;      memory[62756] <=  8'h00;      memory[62757] <=  8'h00;      memory[62758] <=  8'h00;      memory[62759] <=  8'h00;      memory[62760] <=  8'h00;      memory[62761] <=  8'h00;      memory[62762] <=  8'h00;      memory[62763] <=  8'h00;      memory[62764] <=  8'h00;      memory[62765] <=  8'h00;      memory[62766] <=  8'h00;      memory[62767] <=  8'h00;      memory[62768] <=  8'h00;      memory[62769] <=  8'h00;      memory[62770] <=  8'h00;      memory[62771] <=  8'h00;      memory[62772] <=  8'h00;      memory[62773] <=  8'h00;      memory[62774] <=  8'h00;      memory[62775] <=  8'h00;      memory[62776] <=  8'h00;      memory[62777] <=  8'h00;      memory[62778] <=  8'h00;      memory[62779] <=  8'h00;      memory[62780] <=  8'h00;      memory[62781] <=  8'h00;      memory[62782] <=  8'h00;      memory[62783] <=  8'h00;      memory[62784] <=  8'h00;      memory[62785] <=  8'h00;      memory[62786] <=  8'h00;      memory[62787] <=  8'h00;      memory[62788] <=  8'h00;      memory[62789] <=  8'h00;      memory[62790] <=  8'h00;      memory[62791] <=  8'h00;      memory[62792] <=  8'h00;      memory[62793] <=  8'h00;      memory[62794] <=  8'h00;      memory[62795] <=  8'h00;      memory[62796] <=  8'h00;      memory[62797] <=  8'h00;      memory[62798] <=  8'h00;      memory[62799] <=  8'h00;      memory[62800] <=  8'h00;      memory[62801] <=  8'h00;      memory[62802] <=  8'h00;      memory[62803] <=  8'h00;      memory[62804] <=  8'h00;      memory[62805] <=  8'h00;      memory[62806] <=  8'h00;      memory[62807] <=  8'h00;      memory[62808] <=  8'h00;      memory[62809] <=  8'h00;      memory[62810] <=  8'h00;      memory[62811] <=  8'h00;      memory[62812] <=  8'h00;      memory[62813] <=  8'h00;      memory[62814] <=  8'h00;      memory[62815] <=  8'h00;      memory[62816] <=  8'h00;      memory[62817] <=  8'h00;      memory[62818] <=  8'h00;      memory[62819] <=  8'h00;      memory[62820] <=  8'h00;      memory[62821] <=  8'h00;      memory[62822] <=  8'h00;      memory[62823] <=  8'h00;      memory[62824] <=  8'h00;      memory[62825] <=  8'h00;      memory[62826] <=  8'h00;      memory[62827] <=  8'h00;      memory[62828] <=  8'h00;      memory[62829] <=  8'h00;      memory[62830] <=  8'h00;      memory[62831] <=  8'h00;      memory[62832] <=  8'h00;      memory[62833] <=  8'h00;      memory[62834] <=  8'h00;      memory[62835] <=  8'h00;      memory[62836] <=  8'h00;      memory[62837] <=  8'h00;      memory[62838] <=  8'h00;      memory[62839] <=  8'h00;      memory[62840] <=  8'h00;      memory[62841] <=  8'h00;      memory[62842] <=  8'h00;      memory[62843] <=  8'h00;      memory[62844] <=  8'h00;      memory[62845] <=  8'h00;      memory[62846] <=  8'h00;      memory[62847] <=  8'h00;      memory[62848] <=  8'h00;      memory[62849] <=  8'h00;      memory[62850] <=  8'h00;      memory[62851] <=  8'h00;      memory[62852] <=  8'h00;      memory[62853] <=  8'h00;      memory[62854] <=  8'h00;      memory[62855] <=  8'h00;      memory[62856] <=  8'h00;      memory[62857] <=  8'h00;      memory[62858] <=  8'h00;      memory[62859] <=  8'h00;      memory[62860] <=  8'h00;      memory[62861] <=  8'h00;      memory[62862] <=  8'h00;      memory[62863] <=  8'h00;      memory[62864] <=  8'h00;      memory[62865] <=  8'h00;      memory[62866] <=  8'h00;      memory[62867] <=  8'h00;      memory[62868] <=  8'h00;      memory[62869] <=  8'h00;      memory[62870] <=  8'h00;      memory[62871] <=  8'h00;      memory[62872] <=  8'h00;      memory[62873] <=  8'h00;      memory[62874] <=  8'h00;      memory[62875] <=  8'h00;      memory[62876] <=  8'h00;      memory[62877] <=  8'h00;      memory[62878] <=  8'h00;      memory[62879] <=  8'h00;      memory[62880] <=  8'h00;      memory[62881] <=  8'h00;      memory[62882] <=  8'h00;      memory[62883] <=  8'h00;      memory[62884] <=  8'h00;      memory[62885] <=  8'h00;      memory[62886] <=  8'h00;      memory[62887] <=  8'h00;      memory[62888] <=  8'h00;      memory[62889] <=  8'h00;      memory[62890] <=  8'h00;      memory[62891] <=  8'h00;      memory[62892] <=  8'h00;      memory[62893] <=  8'h00;      memory[62894] <=  8'h00;      memory[62895] <=  8'h00;      memory[62896] <=  8'h00;      memory[62897] <=  8'h00;      memory[62898] <=  8'h00;      memory[62899] <=  8'h00;      memory[62900] <=  8'h00;      memory[62901] <=  8'h00;      memory[62902] <=  8'h00;      memory[62903] <=  8'h00;      memory[62904] <=  8'h00;      memory[62905] <=  8'h00;      memory[62906] <=  8'h00;      memory[62907] <=  8'h00;      memory[62908] <=  8'h00;      memory[62909] <=  8'h00;      memory[62910] <=  8'h00;      memory[62911] <=  8'h00;      memory[62912] <=  8'h00;      memory[62913] <=  8'h00;      memory[62914] <=  8'h00;      memory[62915] <=  8'h00;      memory[62916] <=  8'h00;      memory[62917] <=  8'h00;      memory[62918] <=  8'h00;      memory[62919] <=  8'h00;      memory[62920] <=  8'h00;      memory[62921] <=  8'h00;      memory[62922] <=  8'h00;      memory[62923] <=  8'h00;      memory[62924] <=  8'h00;      memory[62925] <=  8'h00;      memory[62926] <=  8'h00;      memory[62927] <=  8'h00;      memory[62928] <=  8'h00;      memory[62929] <=  8'h00;      memory[62930] <=  8'h00;      memory[62931] <=  8'h00;      memory[62932] <=  8'h00;      memory[62933] <=  8'h00;      memory[62934] <=  8'h00;      memory[62935] <=  8'h00;      memory[62936] <=  8'h00;      memory[62937] <=  8'h00;      memory[62938] <=  8'h00;      memory[62939] <=  8'h00;      memory[62940] <=  8'h00;      memory[62941] <=  8'h00;      memory[62942] <=  8'h00;      memory[62943] <=  8'h00;      memory[62944] <=  8'h00;      memory[62945] <=  8'h00;      memory[62946] <=  8'h00;      memory[62947] <=  8'h00;      memory[62948] <=  8'h00;      memory[62949] <=  8'h00;      memory[62950] <=  8'h00;      memory[62951] <=  8'h00;      memory[62952] <=  8'h00;      memory[62953] <=  8'h00;      memory[62954] <=  8'h00;      memory[62955] <=  8'h00;      memory[62956] <=  8'h00;      memory[62957] <=  8'h00;      memory[62958] <=  8'h00;      memory[62959] <=  8'h00;      memory[62960] <=  8'h00;      memory[62961] <=  8'h00;      memory[62962] <=  8'h00;      memory[62963] <=  8'h00;      memory[62964] <=  8'h00;      memory[62965] <=  8'h00;      memory[62966] <=  8'h00;      memory[62967] <=  8'h00;      memory[62968] <=  8'h00;      memory[62969] <=  8'h00;      memory[62970] <=  8'h00;      memory[62971] <=  8'h00;      memory[62972] <=  8'h00;      memory[62973] <=  8'h00;      memory[62974] <=  8'h00;      memory[62975] <=  8'h00;      memory[62976] <=  8'h00;      memory[62977] <=  8'h00;      memory[62978] <=  8'h00;      memory[62979] <=  8'h00;      memory[62980] <=  8'h00;      memory[62981] <=  8'h00;      memory[62982] <=  8'h00;      memory[62983] <=  8'h00;      memory[62984] <=  8'h00;      memory[62985] <=  8'h00;      memory[62986] <=  8'h00;      memory[62987] <=  8'h00;      memory[62988] <=  8'h00;      memory[62989] <=  8'h00;      memory[62990] <=  8'h00;      memory[62991] <=  8'h00;      memory[62992] <=  8'h00;      memory[62993] <=  8'h00;      memory[62994] <=  8'h00;      memory[62995] <=  8'h00;      memory[62996] <=  8'h00;      memory[62997] <=  8'h00;      memory[62998] <=  8'h00;      memory[62999] <=  8'h00;      memory[63000] <=  8'h00;      memory[63001] <=  8'h00;      memory[63002] <=  8'h00;      memory[63003] <=  8'h00;      memory[63004] <=  8'h00;      memory[63005] <=  8'h00;      memory[63006] <=  8'h00;      memory[63007] <=  8'h00;      memory[63008] <=  8'h00;      memory[63009] <=  8'h00;      memory[63010] <=  8'h00;      memory[63011] <=  8'h00;      memory[63012] <=  8'h00;      memory[63013] <=  8'h00;      memory[63014] <=  8'h00;      memory[63015] <=  8'h00;      memory[63016] <=  8'h00;      memory[63017] <=  8'h00;      memory[63018] <=  8'h00;      memory[63019] <=  8'h00;      memory[63020] <=  8'h00;      memory[63021] <=  8'h00;      memory[63022] <=  8'h00;      memory[63023] <=  8'h00;      memory[63024] <=  8'h00;      memory[63025] <=  8'h00;      memory[63026] <=  8'h00;      memory[63027] <=  8'h00;      memory[63028] <=  8'h00;      memory[63029] <=  8'h00;      memory[63030] <=  8'h00;      memory[63031] <=  8'h00;      memory[63032] <=  8'h00;      memory[63033] <=  8'h00;      memory[63034] <=  8'h00;      memory[63035] <=  8'h00;      memory[63036] <=  8'h00;      memory[63037] <=  8'h00;      memory[63038] <=  8'h00;      memory[63039] <=  8'h00;      memory[63040] <=  8'h00;      memory[63041] <=  8'h00;      memory[63042] <=  8'h00;      memory[63043] <=  8'h00;      memory[63044] <=  8'h00;      memory[63045] <=  8'h00;      memory[63046] <=  8'h00;      memory[63047] <=  8'h00;      memory[63048] <=  8'h00;      memory[63049] <=  8'h00;      memory[63050] <=  8'h00;      memory[63051] <=  8'h00;      memory[63052] <=  8'h00;      memory[63053] <=  8'h00;      memory[63054] <=  8'h00;      memory[63055] <=  8'h00;      memory[63056] <=  8'h00;      memory[63057] <=  8'h00;      memory[63058] <=  8'h00;      memory[63059] <=  8'h00;      memory[63060] <=  8'h00;      memory[63061] <=  8'h00;      memory[63062] <=  8'h00;      memory[63063] <=  8'h00;      memory[63064] <=  8'h00;      memory[63065] <=  8'h00;      memory[63066] <=  8'h00;      memory[63067] <=  8'h00;      memory[63068] <=  8'h00;      memory[63069] <=  8'h00;      memory[63070] <=  8'h00;      memory[63071] <=  8'h00;      memory[63072] <=  8'h00;      memory[63073] <=  8'h00;      memory[63074] <=  8'h00;      memory[63075] <=  8'h00;      memory[63076] <=  8'h00;      memory[63077] <=  8'h00;      memory[63078] <=  8'h00;      memory[63079] <=  8'h00;      memory[63080] <=  8'h00;      memory[63081] <=  8'h00;      memory[63082] <=  8'h00;      memory[63083] <=  8'h00;      memory[63084] <=  8'h00;      memory[63085] <=  8'h00;      memory[63086] <=  8'h00;      memory[63087] <=  8'h00;      memory[63088] <=  8'h00;      memory[63089] <=  8'h00;      memory[63090] <=  8'h00;      memory[63091] <=  8'h00;      memory[63092] <=  8'h00;      memory[63093] <=  8'h00;      memory[63094] <=  8'h00;      memory[63095] <=  8'h00;      memory[63096] <=  8'h00;      memory[63097] <=  8'h00;      memory[63098] <=  8'h00;      memory[63099] <=  8'h00;      memory[63100] <=  8'h00;      memory[63101] <=  8'h00;      memory[63102] <=  8'h00;      memory[63103] <=  8'h00;      memory[63104] <=  8'h00;      memory[63105] <=  8'h00;      memory[63106] <=  8'h00;      memory[63107] <=  8'h00;      memory[63108] <=  8'h00;      memory[63109] <=  8'h00;      memory[63110] <=  8'h00;      memory[63111] <=  8'h00;      memory[63112] <=  8'h00;      memory[63113] <=  8'h00;      memory[63114] <=  8'h00;      memory[63115] <=  8'h00;      memory[63116] <=  8'h00;      memory[63117] <=  8'h00;      memory[63118] <=  8'h00;      memory[63119] <=  8'h00;      memory[63120] <=  8'h00;      memory[63121] <=  8'h00;      memory[63122] <=  8'h00;      memory[63123] <=  8'h00;      memory[63124] <=  8'h00;      memory[63125] <=  8'h00;      memory[63126] <=  8'h00;      memory[63127] <=  8'h00;      memory[63128] <=  8'h00;      memory[63129] <=  8'h00;      memory[63130] <=  8'h00;      memory[63131] <=  8'h00;      memory[63132] <=  8'h00;      memory[63133] <=  8'h00;      memory[63134] <=  8'h00;      memory[63135] <=  8'h00;      memory[63136] <=  8'h00;      memory[63137] <=  8'h00;      memory[63138] <=  8'h00;      memory[63139] <=  8'h00;      memory[63140] <=  8'h00;      memory[63141] <=  8'h00;      memory[63142] <=  8'h00;      memory[63143] <=  8'h00;      memory[63144] <=  8'h00;      memory[63145] <=  8'h00;      memory[63146] <=  8'h00;      memory[63147] <=  8'h00;      memory[63148] <=  8'h00;      memory[63149] <=  8'h00;      memory[63150] <=  8'h00;      memory[63151] <=  8'h00;      memory[63152] <=  8'h00;      memory[63153] <=  8'h00;      memory[63154] <=  8'h00;      memory[63155] <=  8'h00;      memory[63156] <=  8'h00;      memory[63157] <=  8'h00;      memory[63158] <=  8'h00;      memory[63159] <=  8'h00;      memory[63160] <=  8'h00;      memory[63161] <=  8'h00;      memory[63162] <=  8'h00;      memory[63163] <=  8'h00;      memory[63164] <=  8'h00;      memory[63165] <=  8'h00;      memory[63166] <=  8'h00;      memory[63167] <=  8'h00;      memory[63168] <=  8'h00;      memory[63169] <=  8'h00;      memory[63170] <=  8'h00;      memory[63171] <=  8'h00;      memory[63172] <=  8'h00;      memory[63173] <=  8'h00;      memory[63174] <=  8'h00;      memory[63175] <=  8'h00;      memory[63176] <=  8'h00;      memory[63177] <=  8'h00;      memory[63178] <=  8'h00;      memory[63179] <=  8'h00;      memory[63180] <=  8'h00;      memory[63181] <=  8'h00;      memory[63182] <=  8'h00;      memory[63183] <=  8'h00;      memory[63184] <=  8'h00;      memory[63185] <=  8'h00;      memory[63186] <=  8'h00;      memory[63187] <=  8'h00;      memory[63188] <=  8'h00;      memory[63189] <=  8'h00;      memory[63190] <=  8'h00;      memory[63191] <=  8'h00;      memory[63192] <=  8'h00;      memory[63193] <=  8'h00;      memory[63194] <=  8'h00;      memory[63195] <=  8'h00;      memory[63196] <=  8'h00;      memory[63197] <=  8'h00;      memory[63198] <=  8'h00;      memory[63199] <=  8'h00;      memory[63200] <=  8'h00;      memory[63201] <=  8'h00;      memory[63202] <=  8'h00;      memory[63203] <=  8'h00;      memory[63204] <=  8'h00;      memory[63205] <=  8'h00;      memory[63206] <=  8'h00;      memory[63207] <=  8'h00;      memory[63208] <=  8'h00;      memory[63209] <=  8'h00;      memory[63210] <=  8'h00;      memory[63211] <=  8'h00;      memory[63212] <=  8'h00;      memory[63213] <=  8'h00;      memory[63214] <=  8'h00;      memory[63215] <=  8'h00;      memory[63216] <=  8'h00;      memory[63217] <=  8'h00;      memory[63218] <=  8'h00;      memory[63219] <=  8'h00;      memory[63220] <=  8'h00;      memory[63221] <=  8'h00;      memory[63222] <=  8'h00;      memory[63223] <=  8'h00;      memory[63224] <=  8'h00;      memory[63225] <=  8'h00;      memory[63226] <=  8'h00;      memory[63227] <=  8'h00;      memory[63228] <=  8'h00;      memory[63229] <=  8'h00;      memory[63230] <=  8'h00;      memory[63231] <=  8'h00;      memory[63232] <=  8'h00;      memory[63233] <=  8'h00;      memory[63234] <=  8'h00;      memory[63235] <=  8'h00;      memory[63236] <=  8'h00;      memory[63237] <=  8'h00;      memory[63238] <=  8'h00;      memory[63239] <=  8'h00;      memory[63240] <=  8'h00;      memory[63241] <=  8'h00;      memory[63242] <=  8'h00;      memory[63243] <=  8'h00;      memory[63244] <=  8'h00;      memory[63245] <=  8'h00;      memory[63246] <=  8'h00;      memory[63247] <=  8'h00;      memory[63248] <=  8'h00;      memory[63249] <=  8'h00;      memory[63250] <=  8'h00;      memory[63251] <=  8'h00;      memory[63252] <=  8'h00;      memory[63253] <=  8'h00;      memory[63254] <=  8'h00;      memory[63255] <=  8'h00;      memory[63256] <=  8'h00;      memory[63257] <=  8'h00;      memory[63258] <=  8'h00;      memory[63259] <=  8'h00;      memory[63260] <=  8'h00;      memory[63261] <=  8'h00;      memory[63262] <=  8'h00;      memory[63263] <=  8'h00;      memory[63264] <=  8'h00;      memory[63265] <=  8'h00;      memory[63266] <=  8'h00;      memory[63267] <=  8'h00;      memory[63268] <=  8'h00;      memory[63269] <=  8'h00;      memory[63270] <=  8'h00;      memory[63271] <=  8'h00;      memory[63272] <=  8'h00;      memory[63273] <=  8'h00;      memory[63274] <=  8'h00;      memory[63275] <=  8'h00;      memory[63276] <=  8'h00;      memory[63277] <=  8'h00;      memory[63278] <=  8'h00;      memory[63279] <=  8'h00;      memory[63280] <=  8'h00;      memory[63281] <=  8'h00;      memory[63282] <=  8'h00;      memory[63283] <=  8'h00;      memory[63284] <=  8'h00;      memory[63285] <=  8'h00;      memory[63286] <=  8'h00;      memory[63287] <=  8'h00;      memory[63288] <=  8'h00;      memory[63289] <=  8'h00;      memory[63290] <=  8'h00;      memory[63291] <=  8'h00;      memory[63292] <=  8'h00;      memory[63293] <=  8'h00;      memory[63294] <=  8'h00;      memory[63295] <=  8'h00;      memory[63296] <=  8'h00;      memory[63297] <=  8'h00;      memory[63298] <=  8'h00;      memory[63299] <=  8'h00;      memory[63300] <=  8'h00;      memory[63301] <=  8'h00;      memory[63302] <=  8'h00;      memory[63303] <=  8'h00;      memory[63304] <=  8'h00;      memory[63305] <=  8'h00;      memory[63306] <=  8'h00;      memory[63307] <=  8'h00;      memory[63308] <=  8'h00;      memory[63309] <=  8'h00;      memory[63310] <=  8'h00;      memory[63311] <=  8'h00;      memory[63312] <=  8'h00;      memory[63313] <=  8'h00;      memory[63314] <=  8'h00;      memory[63315] <=  8'h00;      memory[63316] <=  8'h00;      memory[63317] <=  8'h00;      memory[63318] <=  8'h00;      memory[63319] <=  8'h00;      memory[63320] <=  8'h00;      memory[63321] <=  8'h00;      memory[63322] <=  8'h00;      memory[63323] <=  8'h00;      memory[63324] <=  8'h00;      memory[63325] <=  8'h00;      memory[63326] <=  8'h00;      memory[63327] <=  8'h00;      memory[63328] <=  8'h00;      memory[63329] <=  8'h00;      memory[63330] <=  8'h00;      memory[63331] <=  8'h00;      memory[63332] <=  8'h00;      memory[63333] <=  8'h00;      memory[63334] <=  8'h00;      memory[63335] <=  8'h00;      memory[63336] <=  8'h00;      memory[63337] <=  8'h00;      memory[63338] <=  8'h00;      memory[63339] <=  8'h00;      memory[63340] <=  8'h00;      memory[63341] <=  8'h00;      memory[63342] <=  8'h00;      memory[63343] <=  8'h00;      memory[63344] <=  8'h00;      memory[63345] <=  8'h00;      memory[63346] <=  8'h00;      memory[63347] <=  8'h00;      memory[63348] <=  8'h00;      memory[63349] <=  8'h00;      memory[63350] <=  8'h00;      memory[63351] <=  8'h00;      memory[63352] <=  8'h00;      memory[63353] <=  8'h00;      memory[63354] <=  8'h00;      memory[63355] <=  8'h00;      memory[63356] <=  8'h00;      memory[63357] <=  8'h00;      memory[63358] <=  8'h00;      memory[63359] <=  8'h00;      memory[63360] <=  8'h00;      memory[63361] <=  8'h00;      memory[63362] <=  8'h00;      memory[63363] <=  8'h00;      memory[63364] <=  8'h00;      memory[63365] <=  8'h00;      memory[63366] <=  8'h00;      memory[63367] <=  8'h00;      memory[63368] <=  8'h00;      memory[63369] <=  8'h00;      memory[63370] <=  8'h00;      memory[63371] <=  8'h00;      memory[63372] <=  8'h00;      memory[63373] <=  8'h00;      memory[63374] <=  8'h00;      memory[63375] <=  8'h00;      memory[63376] <=  8'h00;      memory[63377] <=  8'h00;      memory[63378] <=  8'h00;      memory[63379] <=  8'h00;      memory[63380] <=  8'h00;      memory[63381] <=  8'h00;      memory[63382] <=  8'h00;      memory[63383] <=  8'h00;      memory[63384] <=  8'h00;      memory[63385] <=  8'h00;      memory[63386] <=  8'h00;      memory[63387] <=  8'h00;      memory[63388] <=  8'h00;      memory[63389] <=  8'h00;      memory[63390] <=  8'h00;      memory[63391] <=  8'h00;      memory[63392] <=  8'h00;      memory[63393] <=  8'h00;      memory[63394] <=  8'h00;      memory[63395] <=  8'h00;      memory[63396] <=  8'h00;      memory[63397] <=  8'h00;      memory[63398] <=  8'h00;      memory[63399] <=  8'h00;      memory[63400] <=  8'h00;      memory[63401] <=  8'h00;      memory[63402] <=  8'h00;      memory[63403] <=  8'h00;      memory[63404] <=  8'h00;      memory[63405] <=  8'h00;      memory[63406] <=  8'h00;      memory[63407] <=  8'h00;      memory[63408] <=  8'h00;      memory[63409] <=  8'h00;      memory[63410] <=  8'h00;      memory[63411] <=  8'h00;      memory[63412] <=  8'h00;      memory[63413] <=  8'h00;      memory[63414] <=  8'h00;      memory[63415] <=  8'h00;      memory[63416] <=  8'h00;      memory[63417] <=  8'h00;      memory[63418] <=  8'h00;      memory[63419] <=  8'h00;      memory[63420] <=  8'h00;      memory[63421] <=  8'h00;      memory[63422] <=  8'h00;      memory[63423] <=  8'h00;      memory[63424] <=  8'h00;      memory[63425] <=  8'h00;      memory[63426] <=  8'h00;      memory[63427] <=  8'h00;      memory[63428] <=  8'h00;      memory[63429] <=  8'h00;      memory[63430] <=  8'h00;      memory[63431] <=  8'h00;      memory[63432] <=  8'h00;      memory[63433] <=  8'h00;      memory[63434] <=  8'h00;      memory[63435] <=  8'h00;      memory[63436] <=  8'h00;      memory[63437] <=  8'h00;      memory[63438] <=  8'h00;      memory[63439] <=  8'h00;      memory[63440] <=  8'h00;      memory[63441] <=  8'h00;      memory[63442] <=  8'h00;      memory[63443] <=  8'h00;      memory[63444] <=  8'h00;      memory[63445] <=  8'h00;      memory[63446] <=  8'h00;      memory[63447] <=  8'h00;      memory[63448] <=  8'h00;      memory[63449] <=  8'h00;      memory[63450] <=  8'h00;      memory[63451] <=  8'h00;      memory[63452] <=  8'h00;      memory[63453] <=  8'h00;      memory[63454] <=  8'h00;      memory[63455] <=  8'h00;      memory[63456] <=  8'h00;      memory[63457] <=  8'h00;      memory[63458] <=  8'h00;      memory[63459] <=  8'h00;      memory[63460] <=  8'h00;      memory[63461] <=  8'h00;      memory[63462] <=  8'h00;      memory[63463] <=  8'h00;      memory[63464] <=  8'h00;      memory[63465] <=  8'h00;      memory[63466] <=  8'h00;      memory[63467] <=  8'h00;      memory[63468] <=  8'h00;      memory[63469] <=  8'h00;      memory[63470] <=  8'h00;      memory[63471] <=  8'h00;      memory[63472] <=  8'h00;      memory[63473] <=  8'h00;      memory[63474] <=  8'h00;      memory[63475] <=  8'h00;      memory[63476] <=  8'h00;      memory[63477] <=  8'h00;      memory[63478] <=  8'h00;      memory[63479] <=  8'h00;      memory[63480] <=  8'h00;      memory[63481] <=  8'h00;      memory[63482] <=  8'h00;      memory[63483] <=  8'h00;      memory[63484] <=  8'h00;      memory[63485] <=  8'h00;      memory[63486] <=  8'h00;      memory[63487] <=  8'h00;      memory[63488] <=  8'h00;      memory[63489] <=  8'h00;      memory[63490] <=  8'h00;      memory[63491] <=  8'h00;      memory[63492] <=  8'h00;      memory[63493] <=  8'h00;      memory[63494] <=  8'h00;      memory[63495] <=  8'h00;      memory[63496] <=  8'h00;      memory[63497] <=  8'h00;      memory[63498] <=  8'h00;      memory[63499] <=  8'h00;      memory[63500] <=  8'h00;      memory[63501] <=  8'h00;      memory[63502] <=  8'h00;      memory[63503] <=  8'h00;      memory[63504] <=  8'h00;      memory[63505] <=  8'h00;      memory[63506] <=  8'h00;      memory[63507] <=  8'h00;      memory[63508] <=  8'h00;      memory[63509] <=  8'h00;      memory[63510] <=  8'h00;      memory[63511] <=  8'h00;      memory[63512] <=  8'h00;      memory[63513] <=  8'h00;      memory[63514] <=  8'h00;      memory[63515] <=  8'h00;      memory[63516] <=  8'h00;      memory[63517] <=  8'h00;      memory[63518] <=  8'h00;      memory[63519] <=  8'h00;      memory[63520] <=  8'h00;      memory[63521] <=  8'h00;      memory[63522] <=  8'h00;      memory[63523] <=  8'h00;      memory[63524] <=  8'h00;      memory[63525] <=  8'h00;      memory[63526] <=  8'h00;      memory[63527] <=  8'h00;      memory[63528] <=  8'h00;      memory[63529] <=  8'h00;      memory[63530] <=  8'h00;      memory[63531] <=  8'h00;      memory[63532] <=  8'h00;      memory[63533] <=  8'h00;      memory[63534] <=  8'h00;      memory[63535] <=  8'h00;      memory[63536] <=  8'h00;      memory[63537] <=  8'h00;      memory[63538] <=  8'h00;      memory[63539] <=  8'h00;      memory[63540] <=  8'h00;      memory[63541] <=  8'h00;      memory[63542] <=  8'h00;      memory[63543] <=  8'h00;      memory[63544] <=  8'h00;      memory[63545] <=  8'h00;      memory[63546] <=  8'h00;      memory[63547] <=  8'h00;      memory[63548] <=  8'h00;      memory[63549] <=  8'h00;      memory[63550] <=  8'h00;      memory[63551] <=  8'h00;      memory[63552] <=  8'h00;      memory[63553] <=  8'h00;      memory[63554] <=  8'h00;      memory[63555] <=  8'h00;      memory[63556] <=  8'h00;      memory[63557] <=  8'h00;      memory[63558] <=  8'h00;      memory[63559] <=  8'h00;      memory[63560] <=  8'h00;      memory[63561] <=  8'h00;      memory[63562] <=  8'h00;      memory[63563] <=  8'h00;      memory[63564] <=  8'h00;      memory[63565] <=  8'h00;      memory[63566] <=  8'h00;      memory[63567] <=  8'h00;      memory[63568] <=  8'h00;      memory[63569] <=  8'h00;      memory[63570] <=  8'h00;      memory[63571] <=  8'h00;      memory[63572] <=  8'h00;      memory[63573] <=  8'h00;      memory[63574] <=  8'h00;      memory[63575] <=  8'h00;      memory[63576] <=  8'h00;      memory[63577] <=  8'h00;      memory[63578] <=  8'h00;      memory[63579] <=  8'h00;      memory[63580] <=  8'h00;      memory[63581] <=  8'h00;      memory[63582] <=  8'h00;      memory[63583] <=  8'h00;      memory[63584] <=  8'h00;      memory[63585] <=  8'h00;      memory[63586] <=  8'h00;      memory[63587] <=  8'h00;      memory[63588] <=  8'h00;      memory[63589] <=  8'h00;      memory[63590] <=  8'h00;      memory[63591] <=  8'h00;      memory[63592] <=  8'h00;      memory[63593] <=  8'h00;      memory[63594] <=  8'h00;      memory[63595] <=  8'h00;      memory[63596] <=  8'h00;      memory[63597] <=  8'h00;      memory[63598] <=  8'h00;      memory[63599] <=  8'h00;      memory[63600] <=  8'h00;      memory[63601] <=  8'h00;      memory[63602] <=  8'h00;      memory[63603] <=  8'h00;      memory[63604] <=  8'h00;      memory[63605] <=  8'h00;      memory[63606] <=  8'h00;      memory[63607] <=  8'h00;      memory[63608] <=  8'h00;      memory[63609] <=  8'h00;      memory[63610] <=  8'h00;      memory[63611] <=  8'h00;      memory[63612] <=  8'h00;      memory[63613] <=  8'h00;      memory[63614] <=  8'h00;      memory[63615] <=  8'h00;      memory[63616] <=  8'h00;      memory[63617] <=  8'h00;      memory[63618] <=  8'h00;      memory[63619] <=  8'h00;      memory[63620] <=  8'h00;      memory[63621] <=  8'h00;      memory[63622] <=  8'h00;      memory[63623] <=  8'h00;      memory[63624] <=  8'h00;      memory[63625] <=  8'h00;      memory[63626] <=  8'h00;      memory[63627] <=  8'h00;      memory[63628] <=  8'h00;      memory[63629] <=  8'h00;      memory[63630] <=  8'h00;      memory[63631] <=  8'h00;      memory[63632] <=  8'h00;      memory[63633] <=  8'h00;      memory[63634] <=  8'h00;      memory[63635] <=  8'h00;      memory[63636] <=  8'h00;      memory[63637] <=  8'h00;      memory[63638] <=  8'h00;      memory[63639] <=  8'h00;      memory[63640] <=  8'h00;      memory[63641] <=  8'h00;      memory[63642] <=  8'h00;      memory[63643] <=  8'h00;      memory[63644] <=  8'h00;      memory[63645] <=  8'h00;      memory[63646] <=  8'h00;      memory[63647] <=  8'h00;      memory[63648] <=  8'h00;      memory[63649] <=  8'h00;      memory[63650] <=  8'h00;      memory[63651] <=  8'h00;      memory[63652] <=  8'h00;      memory[63653] <=  8'h00;      memory[63654] <=  8'h00;      memory[63655] <=  8'h00;      memory[63656] <=  8'h00;      memory[63657] <=  8'h00;      memory[63658] <=  8'h00;      memory[63659] <=  8'h00;      memory[63660] <=  8'h00;      memory[63661] <=  8'h00;      memory[63662] <=  8'h00;      memory[63663] <=  8'h00;      memory[63664] <=  8'h00;      memory[63665] <=  8'h00;      memory[63666] <=  8'h00;      memory[63667] <=  8'h00;      memory[63668] <=  8'h00;      memory[63669] <=  8'h00;      memory[63670] <=  8'h00;      memory[63671] <=  8'h00;      memory[63672] <=  8'h00;      memory[63673] <=  8'h00;      memory[63674] <=  8'h00;      memory[63675] <=  8'h00;      memory[63676] <=  8'h00;      memory[63677] <=  8'h00;      memory[63678] <=  8'h00;      memory[63679] <=  8'h00;      memory[63680] <=  8'h00;      memory[63681] <=  8'h00;      memory[63682] <=  8'h00;      memory[63683] <=  8'h00;      memory[63684] <=  8'h00;      memory[63685] <=  8'h00;      memory[63686] <=  8'h00;      memory[63687] <=  8'h00;      memory[63688] <=  8'h00;      memory[63689] <=  8'h00;      memory[63690] <=  8'h00;      memory[63691] <=  8'h00;      memory[63692] <=  8'h00;      memory[63693] <=  8'h00;      memory[63694] <=  8'h00;      memory[63695] <=  8'h00;      memory[63696] <=  8'h00;      memory[63697] <=  8'h00;      memory[63698] <=  8'h00;      memory[63699] <=  8'h00;      memory[63700] <=  8'h00;      memory[63701] <=  8'h00;      memory[63702] <=  8'h00;      memory[63703] <=  8'h00;      memory[63704] <=  8'h00;      memory[63705] <=  8'h00;      memory[63706] <=  8'h00;      memory[63707] <=  8'h00;      memory[63708] <=  8'h00;      memory[63709] <=  8'h00;      memory[63710] <=  8'h00;      memory[63711] <=  8'h00;      memory[63712] <=  8'h00;      memory[63713] <=  8'h00;      memory[63714] <=  8'h00;      memory[63715] <=  8'h00;      memory[63716] <=  8'h00;      memory[63717] <=  8'h00;      memory[63718] <=  8'h00;      memory[63719] <=  8'h00;      memory[63720] <=  8'h00;      memory[63721] <=  8'h00;      memory[63722] <=  8'h00;      memory[63723] <=  8'h00;      memory[63724] <=  8'h00;      memory[63725] <=  8'h00;      memory[63726] <=  8'h00;      memory[63727] <=  8'h00;      memory[63728] <=  8'h00;      memory[63729] <=  8'h00;      memory[63730] <=  8'h00;      memory[63731] <=  8'h00;      memory[63732] <=  8'h00;      memory[63733] <=  8'h00;      memory[63734] <=  8'h00;      memory[63735] <=  8'h00;      memory[63736] <=  8'h00;      memory[63737] <=  8'h00;      memory[63738] <=  8'h00;      memory[63739] <=  8'h00;      memory[63740] <=  8'h00;      memory[63741] <=  8'h00;      memory[63742] <=  8'h00;      memory[63743] <=  8'h00;      memory[63744] <=  8'h00;      memory[63745] <=  8'h00;      memory[63746] <=  8'h00;      memory[63747] <=  8'h00;      memory[63748] <=  8'h00;      memory[63749] <=  8'h00;      memory[63750] <=  8'h00;      memory[63751] <=  8'h00;      memory[63752] <=  8'h00;      memory[63753] <=  8'h00;      memory[63754] <=  8'h00;      memory[63755] <=  8'h00;      memory[63756] <=  8'h00;      memory[63757] <=  8'h00;      memory[63758] <=  8'h00;      memory[63759] <=  8'h00;      memory[63760] <=  8'h00;      memory[63761] <=  8'h00;      memory[63762] <=  8'h00;      memory[63763] <=  8'h00;      memory[63764] <=  8'h00;      memory[63765] <=  8'h00;      memory[63766] <=  8'h00;      memory[63767] <=  8'h00;      memory[63768] <=  8'h00;      memory[63769] <=  8'h00;      memory[63770] <=  8'h00;      memory[63771] <=  8'h00;      memory[63772] <=  8'h00;      memory[63773] <=  8'h00;      memory[63774] <=  8'h00;      memory[63775] <=  8'h00;      memory[63776] <=  8'h00;      memory[63777] <=  8'h00;      memory[63778] <=  8'h00;      memory[63779] <=  8'h00;      memory[63780] <=  8'h00;      memory[63781] <=  8'h00;      memory[63782] <=  8'h00;      memory[63783] <=  8'h00;      memory[63784] <=  8'h00;      memory[63785] <=  8'h00;      memory[63786] <=  8'h00;      memory[63787] <=  8'h00;      memory[63788] <=  8'h00;      memory[63789] <=  8'h00;      memory[63790] <=  8'h00;      memory[63791] <=  8'h00;      memory[63792] <=  8'h00;      memory[63793] <=  8'h00;      memory[63794] <=  8'h00;      memory[63795] <=  8'h00;      memory[63796] <=  8'h00;      memory[63797] <=  8'h00;      memory[63798] <=  8'h00;      memory[63799] <=  8'h00;      memory[63800] <=  8'h00;      memory[63801] <=  8'h00;      memory[63802] <=  8'h00;      memory[63803] <=  8'h00;      memory[63804] <=  8'h00;      memory[63805] <=  8'h00;      memory[63806] <=  8'h00;      memory[63807] <=  8'h00;      memory[63808] <=  8'h00;      memory[63809] <=  8'h00;      memory[63810] <=  8'h00;      memory[63811] <=  8'h00;      memory[63812] <=  8'h00;      memory[63813] <=  8'h00;      memory[63814] <=  8'h00;      memory[63815] <=  8'h00;      memory[63816] <=  8'h00;      memory[63817] <=  8'h00;      memory[63818] <=  8'h00;      memory[63819] <=  8'h00;      memory[63820] <=  8'h00;      memory[63821] <=  8'h00;      memory[63822] <=  8'h00;      memory[63823] <=  8'h00;      memory[63824] <=  8'h00;      memory[63825] <=  8'h00;      memory[63826] <=  8'h00;      memory[63827] <=  8'h00;      memory[63828] <=  8'h00;      memory[63829] <=  8'h00;      memory[63830] <=  8'h00;      memory[63831] <=  8'h00;      memory[63832] <=  8'h00;      memory[63833] <=  8'h00;      memory[63834] <=  8'h00;      memory[63835] <=  8'h00;      memory[63836] <=  8'h00;      memory[63837] <=  8'h00;      memory[63838] <=  8'h00;      memory[63839] <=  8'h00;      memory[63840] <=  8'h00;      memory[63841] <=  8'h00;      memory[63842] <=  8'h00;      memory[63843] <=  8'h00;      memory[63844] <=  8'h00;      memory[63845] <=  8'h00;      memory[63846] <=  8'h00;      memory[63847] <=  8'h00;      memory[63848] <=  8'h00;      memory[63849] <=  8'h00;      memory[63850] <=  8'h00;      memory[63851] <=  8'h00;      memory[63852] <=  8'h00;      memory[63853] <=  8'h00;      memory[63854] <=  8'h00;      memory[63855] <=  8'h00;      memory[63856] <=  8'h00;      memory[63857] <=  8'h00;      memory[63858] <=  8'h00;      memory[63859] <=  8'h00;      memory[63860] <=  8'h00;      memory[63861] <=  8'h00;      memory[63862] <=  8'h00;      memory[63863] <=  8'h00;      memory[63864] <=  8'h00;      memory[63865] <=  8'h00;      memory[63866] <=  8'h00;      memory[63867] <=  8'h00;      memory[63868] <=  8'h00;      memory[63869] <=  8'h00;      memory[63870] <=  8'h00;      memory[63871] <=  8'h00;      memory[63872] <=  8'h00;      memory[63873] <=  8'h00;      memory[63874] <=  8'h00;      memory[63875] <=  8'h00;      memory[63876] <=  8'h00;      memory[63877] <=  8'h00;      memory[63878] <=  8'h00;      memory[63879] <=  8'h00;      memory[63880] <=  8'h00;      memory[63881] <=  8'h00;      memory[63882] <=  8'h00;      memory[63883] <=  8'h00;      memory[63884] <=  8'h00;      memory[63885] <=  8'h00;      memory[63886] <=  8'h00;      memory[63887] <=  8'h00;      memory[63888] <=  8'h00;      memory[63889] <=  8'h00;      memory[63890] <=  8'h00;      memory[63891] <=  8'h00;      memory[63892] <=  8'h00;      memory[63893] <=  8'h00;      memory[63894] <=  8'h00;      memory[63895] <=  8'h00;      memory[63896] <=  8'h00;      memory[63897] <=  8'h00;      memory[63898] <=  8'h00;      memory[63899] <=  8'h00;      memory[63900] <=  8'h00;      memory[63901] <=  8'h00;      memory[63902] <=  8'h00;      memory[63903] <=  8'h00;      memory[63904] <=  8'h00;      memory[63905] <=  8'h00;      memory[63906] <=  8'h00;      memory[63907] <=  8'h00;      memory[63908] <=  8'h00;      memory[63909] <=  8'h00;      memory[63910] <=  8'h00;      memory[63911] <=  8'h00;      memory[63912] <=  8'h00;      memory[63913] <=  8'h00;      memory[63914] <=  8'h00;      memory[63915] <=  8'h00;      memory[63916] <=  8'h00;      memory[63917] <=  8'h00;      memory[63918] <=  8'h00;      memory[63919] <=  8'h00;      memory[63920] <=  8'h00;      memory[63921] <=  8'h00;      memory[63922] <=  8'h00;      memory[63923] <=  8'h00;      memory[63924] <=  8'h00;      memory[63925] <=  8'h00;      memory[63926] <=  8'h00;      memory[63927] <=  8'h00;      memory[63928] <=  8'h00;      memory[63929] <=  8'h00;      memory[63930] <=  8'h00;      memory[63931] <=  8'h00;      memory[63932] <=  8'h00;      memory[63933] <=  8'h00;      memory[63934] <=  8'h00;      memory[63935] <=  8'h00;      memory[63936] <=  8'h00;      memory[63937] <=  8'h00;      memory[63938] <=  8'h00;      memory[63939] <=  8'h00;      memory[63940] <=  8'h00;      memory[63941] <=  8'h00;      memory[63942] <=  8'h00;      memory[63943] <=  8'h00;      memory[63944] <=  8'h00;      memory[63945] <=  8'h00;      memory[63946] <=  8'h00;      memory[63947] <=  8'h00;      memory[63948] <=  8'h00;      memory[63949] <=  8'h00;      memory[63950] <=  8'h00;      memory[63951] <=  8'h00;      memory[63952] <=  8'h00;      memory[63953] <=  8'h00;      memory[63954] <=  8'h00;      memory[63955] <=  8'h00;      memory[63956] <=  8'h00;      memory[63957] <=  8'h00;      memory[63958] <=  8'h00;      memory[63959] <=  8'h00;      memory[63960] <=  8'h00;      memory[63961] <=  8'h00;      memory[63962] <=  8'h00;      memory[63963] <=  8'h00;      memory[63964] <=  8'h00;      memory[63965] <=  8'h00;      memory[63966] <=  8'h00;      memory[63967] <=  8'h00;      memory[63968] <=  8'h00;      memory[63969] <=  8'h00;      memory[63970] <=  8'h00;      memory[63971] <=  8'h00;      memory[63972] <=  8'h00;      memory[63973] <=  8'h00;      memory[63974] <=  8'h00;      memory[63975] <=  8'h00;      memory[63976] <=  8'h00;      memory[63977] <=  8'h00;      memory[63978] <=  8'h00;      memory[63979] <=  8'h00;      memory[63980] <=  8'h00;      memory[63981] <=  8'h00;      memory[63982] <=  8'h00;      memory[63983] <=  8'h00;      memory[63984] <=  8'h00;      memory[63985] <=  8'h00;      memory[63986] <=  8'h00;      memory[63987] <=  8'h00;      memory[63988] <=  8'h00;      memory[63989] <=  8'h00;      memory[63990] <=  8'h00;      memory[63991] <=  8'h00;      memory[63992] <=  8'h00;      memory[63993] <=  8'h00;      memory[63994] <=  8'h00;      memory[63995] <=  8'h00;      memory[63996] <=  8'h00;      memory[63997] <=  8'h00;      memory[63998] <=  8'h00;      memory[63999] <=  8'h00;      memory[64000] <=  8'h00;      memory[64001] <=  8'h00;      memory[64002] <=  8'h00;      memory[64003] <=  8'h00;      memory[64004] <=  8'h00;      memory[64005] <=  8'h00;      memory[64006] <=  8'h00;      memory[64007] <=  8'h00;      memory[64008] <=  8'h00;      memory[64009] <=  8'h00;      memory[64010] <=  8'h00;      memory[64011] <=  8'h00;      memory[64012] <=  8'h00;      memory[64013] <=  8'h00;      memory[64014] <=  8'h00;      memory[64015] <=  8'h00;      memory[64016] <=  8'h00;      memory[64017] <=  8'h00;      memory[64018] <=  8'h00;      memory[64019] <=  8'h00;      memory[64020] <=  8'h00;      memory[64021] <=  8'h00;      memory[64022] <=  8'h00;      memory[64023] <=  8'h00;      memory[64024] <=  8'h00;      memory[64025] <=  8'h00;      memory[64026] <=  8'h00;      memory[64027] <=  8'h00;      memory[64028] <=  8'h00;      memory[64029] <=  8'h00;      memory[64030] <=  8'h00;      memory[64031] <=  8'h00;      memory[64032] <=  8'h00;      memory[64033] <=  8'h00;      memory[64034] <=  8'h00;      memory[64035] <=  8'h00;      memory[64036] <=  8'h00;      memory[64037] <=  8'h00;      memory[64038] <=  8'h00;      memory[64039] <=  8'h00;      memory[64040] <=  8'h00;      memory[64041] <=  8'h00;      memory[64042] <=  8'h00;      memory[64043] <=  8'h00;      memory[64044] <=  8'h00;      memory[64045] <=  8'h00;      memory[64046] <=  8'h00;      memory[64047] <=  8'h00;      memory[64048] <=  8'h00;      memory[64049] <=  8'h00;      memory[64050] <=  8'h00;      memory[64051] <=  8'h00;      memory[64052] <=  8'h00;      memory[64053] <=  8'h00;      memory[64054] <=  8'h00;      memory[64055] <=  8'h00;      memory[64056] <=  8'h00;      memory[64057] <=  8'h00;      memory[64058] <=  8'h00;      memory[64059] <=  8'h00;      memory[64060] <=  8'h00;      memory[64061] <=  8'h00;      memory[64062] <=  8'h00;      memory[64063] <=  8'h00;      memory[64064] <=  8'h00;      memory[64065] <=  8'h00;      memory[64066] <=  8'h00;      memory[64067] <=  8'h00;      memory[64068] <=  8'h00;      memory[64069] <=  8'h00;      memory[64070] <=  8'h00;      memory[64071] <=  8'h00;      memory[64072] <=  8'h00;      memory[64073] <=  8'h00;      memory[64074] <=  8'h00;      memory[64075] <=  8'h00;      memory[64076] <=  8'h00;      memory[64077] <=  8'h00;      memory[64078] <=  8'h00;      memory[64079] <=  8'h00;      memory[64080] <=  8'h00;      memory[64081] <=  8'h00;      memory[64082] <=  8'h00;      memory[64083] <=  8'h00;      memory[64084] <=  8'h00;      memory[64085] <=  8'h00;      memory[64086] <=  8'h00;      memory[64087] <=  8'h00;      memory[64088] <=  8'h00;      memory[64089] <=  8'h00;      memory[64090] <=  8'h00;      memory[64091] <=  8'h00;      memory[64092] <=  8'h00;      memory[64093] <=  8'h00;      memory[64094] <=  8'h00;      memory[64095] <=  8'h00;      memory[64096] <=  8'h00;      memory[64097] <=  8'h00;      memory[64098] <=  8'h00;      memory[64099] <=  8'h00;      memory[64100] <=  8'h00;      memory[64101] <=  8'h00;      memory[64102] <=  8'h00;      memory[64103] <=  8'h00;      memory[64104] <=  8'h00;      memory[64105] <=  8'h00;      memory[64106] <=  8'h00;      memory[64107] <=  8'h00;      memory[64108] <=  8'h00;      memory[64109] <=  8'h00;      memory[64110] <=  8'h00;      memory[64111] <=  8'h00;      memory[64112] <=  8'h00;      memory[64113] <=  8'h00;      memory[64114] <=  8'h00;      memory[64115] <=  8'h00;      memory[64116] <=  8'h00;      memory[64117] <=  8'h00;      memory[64118] <=  8'h00;      memory[64119] <=  8'h00;      memory[64120] <=  8'h00;      memory[64121] <=  8'h00;      memory[64122] <=  8'h00;      memory[64123] <=  8'h00;      memory[64124] <=  8'h00;      memory[64125] <=  8'h00;      memory[64126] <=  8'h00;      memory[64127] <=  8'h00;      memory[64128] <=  8'h00;      memory[64129] <=  8'h00;      memory[64130] <=  8'h00;      memory[64131] <=  8'h00;      memory[64132] <=  8'h00;      memory[64133] <=  8'h00;      memory[64134] <=  8'h00;      memory[64135] <=  8'h00;      memory[64136] <=  8'h00;      memory[64137] <=  8'h00;      memory[64138] <=  8'h00;      memory[64139] <=  8'h00;      memory[64140] <=  8'h00;      memory[64141] <=  8'h00;      memory[64142] <=  8'h00;      memory[64143] <=  8'h00;      memory[64144] <=  8'h00;      memory[64145] <=  8'h00;      memory[64146] <=  8'h00;      memory[64147] <=  8'h00;      memory[64148] <=  8'h00;      memory[64149] <=  8'h00;      memory[64150] <=  8'h00;      memory[64151] <=  8'h00;      memory[64152] <=  8'h00;      memory[64153] <=  8'h00;      memory[64154] <=  8'h00;      memory[64155] <=  8'h00;      memory[64156] <=  8'h00;      memory[64157] <=  8'h00;      memory[64158] <=  8'h00;      memory[64159] <=  8'h00;      memory[64160] <=  8'h00;      memory[64161] <=  8'h00;      memory[64162] <=  8'h00;      memory[64163] <=  8'h00;      memory[64164] <=  8'h00;      memory[64165] <=  8'h00;      memory[64166] <=  8'h00;      memory[64167] <=  8'h00;      memory[64168] <=  8'h00;      memory[64169] <=  8'h00;      memory[64170] <=  8'h00;      memory[64171] <=  8'h00;      memory[64172] <=  8'h00;      memory[64173] <=  8'h00;      memory[64174] <=  8'h00;      memory[64175] <=  8'h00;      memory[64176] <=  8'h00;      memory[64177] <=  8'h00;      memory[64178] <=  8'h00;      memory[64179] <=  8'h00;      memory[64180] <=  8'h00;      memory[64181] <=  8'h00;      memory[64182] <=  8'h00;      memory[64183] <=  8'h00;      memory[64184] <=  8'h00;      memory[64185] <=  8'h00;      memory[64186] <=  8'h00;      memory[64187] <=  8'h00;      memory[64188] <=  8'h00;      memory[64189] <=  8'h00;      memory[64190] <=  8'h00;      memory[64191] <=  8'h00;      memory[64192] <=  8'h00;      memory[64193] <=  8'h00;      memory[64194] <=  8'h00;      memory[64195] <=  8'h00;      memory[64196] <=  8'h00;      memory[64197] <=  8'h00;      memory[64198] <=  8'h00;      memory[64199] <=  8'h00;      memory[64200] <=  8'h00;      memory[64201] <=  8'h00;      memory[64202] <=  8'h00;      memory[64203] <=  8'h00;      memory[64204] <=  8'h00;      memory[64205] <=  8'h00;      memory[64206] <=  8'h00;      memory[64207] <=  8'h00;      memory[64208] <=  8'h00;      memory[64209] <=  8'h00;      memory[64210] <=  8'h00;      memory[64211] <=  8'h00;      memory[64212] <=  8'h00;      memory[64213] <=  8'h00;      memory[64214] <=  8'h00;      memory[64215] <=  8'h00;      memory[64216] <=  8'h00;      memory[64217] <=  8'h00;      memory[64218] <=  8'h00;      memory[64219] <=  8'h00;      memory[64220] <=  8'h00;      memory[64221] <=  8'h00;      memory[64222] <=  8'h00;      memory[64223] <=  8'h00;      memory[64224] <=  8'h00;      memory[64225] <=  8'h00;      memory[64226] <=  8'h00;      memory[64227] <=  8'h00;      memory[64228] <=  8'h00;      memory[64229] <=  8'h00;      memory[64230] <=  8'h00;      memory[64231] <=  8'h00;      memory[64232] <=  8'h00;      memory[64233] <=  8'h00;      memory[64234] <=  8'h00;      memory[64235] <=  8'h00;      memory[64236] <=  8'h00;      memory[64237] <=  8'h00;      memory[64238] <=  8'h00;      memory[64239] <=  8'h00;      memory[64240] <=  8'h00;      memory[64241] <=  8'h00;      memory[64242] <=  8'h00;      memory[64243] <=  8'h00;      memory[64244] <=  8'h00;      memory[64245] <=  8'h00;      memory[64246] <=  8'h00;      memory[64247] <=  8'h00;      memory[64248] <=  8'h00;      memory[64249] <=  8'h00;      memory[64250] <=  8'h00;      memory[64251] <=  8'h00;      memory[64252] <=  8'h00;      memory[64253] <=  8'h00;      memory[64254] <=  8'h00;      memory[64255] <=  8'h00;      memory[64256] <=  8'h00;      memory[64257] <=  8'h00;      memory[64258] <=  8'h00;      memory[64259] <=  8'h00;      memory[64260] <=  8'h00;      memory[64261] <=  8'h00;      memory[64262] <=  8'h00;      memory[64263] <=  8'h00;      memory[64264] <=  8'h00;      memory[64265] <=  8'h00;      memory[64266] <=  8'h00;      memory[64267] <=  8'h00;      memory[64268] <=  8'h00;      memory[64269] <=  8'h00;      memory[64270] <=  8'h00;      memory[64271] <=  8'h00;      memory[64272] <=  8'h00;      memory[64273] <=  8'h00;      memory[64274] <=  8'h00;      memory[64275] <=  8'h00;      memory[64276] <=  8'h00;      memory[64277] <=  8'h00;      memory[64278] <=  8'h00;      memory[64279] <=  8'h00;      memory[64280] <=  8'h00;      memory[64281] <=  8'h00;      memory[64282] <=  8'h00;      memory[64283] <=  8'h00;      memory[64284] <=  8'h00;      memory[64285] <=  8'h00;      memory[64286] <=  8'h00;      memory[64287] <=  8'h00;      memory[64288] <=  8'h00;      memory[64289] <=  8'h00;      memory[64290] <=  8'h00;      memory[64291] <=  8'h00;      memory[64292] <=  8'h00;      memory[64293] <=  8'h00;      memory[64294] <=  8'h00;      memory[64295] <=  8'h00;      memory[64296] <=  8'h00;      memory[64297] <=  8'h00;      memory[64298] <=  8'h00;      memory[64299] <=  8'h00;      memory[64300] <=  8'h00;      memory[64301] <=  8'h00;      memory[64302] <=  8'h00;      memory[64303] <=  8'h00;      memory[64304] <=  8'h00;      memory[64305] <=  8'h00;      memory[64306] <=  8'h00;      memory[64307] <=  8'h00;      memory[64308] <=  8'h00;      memory[64309] <=  8'h00;      memory[64310] <=  8'h00;      memory[64311] <=  8'h00;      memory[64312] <=  8'h00;      memory[64313] <=  8'h00;      memory[64314] <=  8'h00;      memory[64315] <=  8'h00;      memory[64316] <=  8'h00;      memory[64317] <=  8'h00;      memory[64318] <=  8'h00;      memory[64319] <=  8'h00;      memory[64320] <=  8'h00;      memory[64321] <=  8'h00;      memory[64322] <=  8'h00;      memory[64323] <=  8'h00;      memory[64324] <=  8'h00;      memory[64325] <=  8'h00;      memory[64326] <=  8'h00;      memory[64327] <=  8'h00;      memory[64328] <=  8'h00;      memory[64329] <=  8'h00;      memory[64330] <=  8'h00;      memory[64331] <=  8'h00;      memory[64332] <=  8'h00;      memory[64333] <=  8'h00;      memory[64334] <=  8'h00;      memory[64335] <=  8'h00;      memory[64336] <=  8'h00;      memory[64337] <=  8'h00;      memory[64338] <=  8'h00;      memory[64339] <=  8'h00;      memory[64340] <=  8'h00;      memory[64341] <=  8'h00;      memory[64342] <=  8'h00;      memory[64343] <=  8'h00;      memory[64344] <=  8'h00;      memory[64345] <=  8'h00;      memory[64346] <=  8'h00;      memory[64347] <=  8'h00;      memory[64348] <=  8'h00;      memory[64349] <=  8'h00;      memory[64350] <=  8'h00;      memory[64351] <=  8'h00;      memory[64352] <=  8'h00;      memory[64353] <=  8'h00;      memory[64354] <=  8'h00;      memory[64355] <=  8'h00;      memory[64356] <=  8'h00;      memory[64357] <=  8'h00;      memory[64358] <=  8'h00;      memory[64359] <=  8'h00;      memory[64360] <=  8'h00;      memory[64361] <=  8'h00;      memory[64362] <=  8'h00;      memory[64363] <=  8'h00;      memory[64364] <=  8'h00;      memory[64365] <=  8'h00;      memory[64366] <=  8'h00;      memory[64367] <=  8'h00;      memory[64368] <=  8'h00;      memory[64369] <=  8'h00;      memory[64370] <=  8'h00;      memory[64371] <=  8'h00;      memory[64372] <=  8'h00;      memory[64373] <=  8'h00;      memory[64374] <=  8'h00;      memory[64375] <=  8'h00;      memory[64376] <=  8'h00;      memory[64377] <=  8'h00;      memory[64378] <=  8'h00;      memory[64379] <=  8'h00;      memory[64380] <=  8'h00;      memory[64381] <=  8'h00;      memory[64382] <=  8'h00;      memory[64383] <=  8'h00;      memory[64384] <=  8'h00;      memory[64385] <=  8'h00;      memory[64386] <=  8'h00;      memory[64387] <=  8'h00;      memory[64388] <=  8'h00;      memory[64389] <=  8'h00;      memory[64390] <=  8'h00;      memory[64391] <=  8'h00;      memory[64392] <=  8'h00;      memory[64393] <=  8'h00;      memory[64394] <=  8'h00;      memory[64395] <=  8'h00;      memory[64396] <=  8'h00;      memory[64397] <=  8'h00;      memory[64398] <=  8'h00;      memory[64399] <=  8'h00;      memory[64400] <=  8'h00;      memory[64401] <=  8'h00;      memory[64402] <=  8'h00;      memory[64403] <=  8'h00;      memory[64404] <=  8'h00;      memory[64405] <=  8'h00;      memory[64406] <=  8'h00;      memory[64407] <=  8'h00;      memory[64408] <=  8'h00;      memory[64409] <=  8'h00;      memory[64410] <=  8'h00;      memory[64411] <=  8'h00;      memory[64412] <=  8'h00;      memory[64413] <=  8'h00;      memory[64414] <=  8'h00;      memory[64415] <=  8'h00;      memory[64416] <=  8'h00;      memory[64417] <=  8'h00;      memory[64418] <=  8'h00;      memory[64419] <=  8'h00;      memory[64420] <=  8'h00;      memory[64421] <=  8'h00;      memory[64422] <=  8'h00;      memory[64423] <=  8'h00;      memory[64424] <=  8'h00;      memory[64425] <=  8'h00;      memory[64426] <=  8'h00;      memory[64427] <=  8'h00;      memory[64428] <=  8'h00;      memory[64429] <=  8'h00;      memory[64430] <=  8'h00;      memory[64431] <=  8'h00;      memory[64432] <=  8'h00;      memory[64433] <=  8'h00;      memory[64434] <=  8'h00;      memory[64435] <=  8'h00;      memory[64436] <=  8'h00;      memory[64437] <=  8'h00;      memory[64438] <=  8'h00;      memory[64439] <=  8'h00;      memory[64440] <=  8'h00;      memory[64441] <=  8'h00;      memory[64442] <=  8'h00;      memory[64443] <=  8'h00;      memory[64444] <=  8'h00;      memory[64445] <=  8'h00;      memory[64446] <=  8'h00;      memory[64447] <=  8'h00;      memory[64448] <=  8'h00;      memory[64449] <=  8'h00;      memory[64450] <=  8'h00;      memory[64451] <=  8'h00;      memory[64452] <=  8'h00;      memory[64453] <=  8'h00;      memory[64454] <=  8'h00;      memory[64455] <=  8'h00;      memory[64456] <=  8'h00;      memory[64457] <=  8'h00;      memory[64458] <=  8'h00;      memory[64459] <=  8'h00;      memory[64460] <=  8'h00;      memory[64461] <=  8'h00;      memory[64462] <=  8'h00;      memory[64463] <=  8'h00;      memory[64464] <=  8'h00;      memory[64465] <=  8'h00;      memory[64466] <=  8'h00;      memory[64467] <=  8'h00;      memory[64468] <=  8'h00;      memory[64469] <=  8'h00;      memory[64470] <=  8'h00;      memory[64471] <=  8'h00;      memory[64472] <=  8'h00;      memory[64473] <=  8'h00;      memory[64474] <=  8'h00;      memory[64475] <=  8'h00;      memory[64476] <=  8'h00;      memory[64477] <=  8'h00;      memory[64478] <=  8'h00;      memory[64479] <=  8'h00;      memory[64480] <=  8'h00;      memory[64481] <=  8'h00;      memory[64482] <=  8'h00;      memory[64483] <=  8'h00;      memory[64484] <=  8'h00;      memory[64485] <=  8'h00;      memory[64486] <=  8'h00;      memory[64487] <=  8'h00;      memory[64488] <=  8'h00;      memory[64489] <=  8'h00;      memory[64490] <=  8'h00;      memory[64491] <=  8'h00;      memory[64492] <=  8'h00;      memory[64493] <=  8'h00;      memory[64494] <=  8'h00;      memory[64495] <=  8'h00;      memory[64496] <=  8'h00;      memory[64497] <=  8'h00;      memory[64498] <=  8'h00;      memory[64499] <=  8'h00;      memory[64500] <=  8'h00;      memory[64501] <=  8'h00;      memory[64502] <=  8'h00;      memory[64503] <=  8'h00;      memory[64504] <=  8'h00;      memory[64505] <=  8'h00;      memory[64506] <=  8'h00;      memory[64507] <=  8'h00;      memory[64508] <=  8'h00;      memory[64509] <=  8'h00;      memory[64510] <=  8'h00;      memory[64511] <=  8'h00;      memory[64512] <=  8'h00;      memory[64513] <=  8'h00;      memory[64514] <=  8'h00;      memory[64515] <=  8'h00;      memory[64516] <=  8'h00;      memory[64517] <=  8'h00;      memory[64518] <=  8'h00;      memory[64519] <=  8'h00;      memory[64520] <=  8'h00;      memory[64521] <=  8'h00;      memory[64522] <=  8'h00;      memory[64523] <=  8'h00;      memory[64524] <=  8'h00;      memory[64525] <=  8'h00;      memory[64526] <=  8'h00;      memory[64527] <=  8'h00;      memory[64528] <=  8'h00;      memory[64529] <=  8'h00;      memory[64530] <=  8'h00;      memory[64531] <=  8'h00;      memory[64532] <=  8'h00;      memory[64533] <=  8'h00;      memory[64534] <=  8'h00;      memory[64535] <=  8'h00;      memory[64536] <=  8'h00;      memory[64537] <=  8'h00;      memory[64538] <=  8'h00;      memory[64539] <=  8'h00;      memory[64540] <=  8'h00;      memory[64541] <=  8'h00;      memory[64542] <=  8'h00;      memory[64543] <=  8'h00;      memory[64544] <=  8'h00;      memory[64545] <=  8'h00;      memory[64546] <=  8'h00;      memory[64547] <=  8'h00;      memory[64548] <=  8'h00;      memory[64549] <=  8'h00;      memory[64550] <=  8'h00;      memory[64551] <=  8'h00;      memory[64552] <=  8'h00;      memory[64553] <=  8'h00;      memory[64554] <=  8'h00;      memory[64555] <=  8'h00;      memory[64556] <=  8'h00;      memory[64557] <=  8'h00;      memory[64558] <=  8'h00;      memory[64559] <=  8'h00;      memory[64560] <=  8'h00;      memory[64561] <=  8'h00;      memory[64562] <=  8'h00;      memory[64563] <=  8'h00;      memory[64564] <=  8'h00;      memory[64565] <=  8'h00;      memory[64566] <=  8'h00;      memory[64567] <=  8'h00;      memory[64568] <=  8'h00;      memory[64569] <=  8'h00;      memory[64570] <=  8'h00;      memory[64571] <=  8'h00;      memory[64572] <=  8'h00;      memory[64573] <=  8'h00;      memory[64574] <=  8'h00;      memory[64575] <=  8'h00;      memory[64576] <=  8'h00;      memory[64577] <=  8'h00;      memory[64578] <=  8'h00;      memory[64579] <=  8'h00;      memory[64580] <=  8'h00;      memory[64581] <=  8'h00;      memory[64582] <=  8'h00;      memory[64583] <=  8'h00;      memory[64584] <=  8'h00;      memory[64585] <=  8'h00;      memory[64586] <=  8'h00;      memory[64587] <=  8'h00;      memory[64588] <=  8'h00;      memory[64589] <=  8'h00;      memory[64590] <=  8'h00;      memory[64591] <=  8'h00;      memory[64592] <=  8'h00;      memory[64593] <=  8'h00;      memory[64594] <=  8'h00;      memory[64595] <=  8'h00;      memory[64596] <=  8'h00;      memory[64597] <=  8'h00;      memory[64598] <=  8'h00;      memory[64599] <=  8'h00;      memory[64600] <=  8'h00;      memory[64601] <=  8'h00;      memory[64602] <=  8'h00;      memory[64603] <=  8'h00;      memory[64604] <=  8'h00;      memory[64605] <=  8'h00;      memory[64606] <=  8'h00;      memory[64607] <=  8'h00;      memory[64608] <=  8'h00;      memory[64609] <=  8'h00;      memory[64610] <=  8'h00;      memory[64611] <=  8'h00;      memory[64612] <=  8'h00;      memory[64613] <=  8'h00;      memory[64614] <=  8'h00;      memory[64615] <=  8'h00;      memory[64616] <=  8'h00;      memory[64617] <=  8'h00;      memory[64618] <=  8'h00;      memory[64619] <=  8'h00;      memory[64620] <=  8'h00;      memory[64621] <=  8'h00;      memory[64622] <=  8'h00;      memory[64623] <=  8'h00;      memory[64624] <=  8'h00;      memory[64625] <=  8'h00;      memory[64626] <=  8'h00;      memory[64627] <=  8'h00;      memory[64628] <=  8'h00;      memory[64629] <=  8'h00;      memory[64630] <=  8'h00;      memory[64631] <=  8'h00;      memory[64632] <=  8'h00;      memory[64633] <=  8'h00;      memory[64634] <=  8'h00;      memory[64635] <=  8'h00;      memory[64636] <=  8'h00;      memory[64637] <=  8'h00;      memory[64638] <=  8'h00;      memory[64639] <=  8'h00;      memory[64640] <=  8'h00;      memory[64641] <=  8'h00;      memory[64642] <=  8'h00;      memory[64643] <=  8'h00;      memory[64644] <=  8'h00;      memory[64645] <=  8'h00;      memory[64646] <=  8'h00;      memory[64647] <=  8'h00;      memory[64648] <=  8'h00;      memory[64649] <=  8'h00;      memory[64650] <=  8'h00;      memory[64651] <=  8'h00;      memory[64652] <=  8'h00;      memory[64653] <=  8'h00;      memory[64654] <=  8'h00;      memory[64655] <=  8'h00;      memory[64656] <=  8'h00;      memory[64657] <=  8'h00;      memory[64658] <=  8'h00;      memory[64659] <=  8'h00;      memory[64660] <=  8'h00;      memory[64661] <=  8'h00;      memory[64662] <=  8'h00;      memory[64663] <=  8'h00;      memory[64664] <=  8'h00;      memory[64665] <=  8'h00;      memory[64666] <=  8'h00;      memory[64667] <=  8'h00;      memory[64668] <=  8'h00;      memory[64669] <=  8'h00;      memory[64670] <=  8'h00;      memory[64671] <=  8'h00;      memory[64672] <=  8'h00;      memory[64673] <=  8'h00;      memory[64674] <=  8'h00;      memory[64675] <=  8'h00;      memory[64676] <=  8'h00;      memory[64677] <=  8'h00;      memory[64678] <=  8'h00;      memory[64679] <=  8'h00;      memory[64680] <=  8'h00;      memory[64681] <=  8'h00;      memory[64682] <=  8'h00;      memory[64683] <=  8'h00;      memory[64684] <=  8'h00;      memory[64685] <=  8'h00;      memory[64686] <=  8'h00;      memory[64687] <=  8'h00;      memory[64688] <=  8'h00;      memory[64689] <=  8'h00;      memory[64690] <=  8'h00;      memory[64691] <=  8'h00;      memory[64692] <=  8'h00;      memory[64693] <=  8'h00;      memory[64694] <=  8'h00;      memory[64695] <=  8'h00;      memory[64696] <=  8'h00;      memory[64697] <=  8'h00;      memory[64698] <=  8'h00;      memory[64699] <=  8'h00;      memory[64700] <=  8'h00;      memory[64701] <=  8'h00;      memory[64702] <=  8'h00;      memory[64703] <=  8'h00;      memory[64704] <=  8'h00;      memory[64705] <=  8'h00;      memory[64706] <=  8'h00;      memory[64707] <=  8'h00;      memory[64708] <=  8'h00;      memory[64709] <=  8'h00;      memory[64710] <=  8'h00;      memory[64711] <=  8'h00;      memory[64712] <=  8'h00;      memory[64713] <=  8'h00;      memory[64714] <=  8'h00;      memory[64715] <=  8'h00;      memory[64716] <=  8'h00;      memory[64717] <=  8'h00;      memory[64718] <=  8'h00;      memory[64719] <=  8'h00;      memory[64720] <=  8'h00;      memory[64721] <=  8'h00;      memory[64722] <=  8'h00;      memory[64723] <=  8'h00;      memory[64724] <=  8'h00;      memory[64725] <=  8'h00;      memory[64726] <=  8'h00;      memory[64727] <=  8'h00;      memory[64728] <=  8'h00;      memory[64729] <=  8'h00;      memory[64730] <=  8'h00;      memory[64731] <=  8'h00;      memory[64732] <=  8'h00;      memory[64733] <=  8'h00;      memory[64734] <=  8'h00;      memory[64735] <=  8'h00;      memory[64736] <=  8'h00;      memory[64737] <=  8'h00;      memory[64738] <=  8'h00;      memory[64739] <=  8'h00;      memory[64740] <=  8'h00;      memory[64741] <=  8'h00;      memory[64742] <=  8'h00;      memory[64743] <=  8'h00;      memory[64744] <=  8'h00;      memory[64745] <=  8'h00;      memory[64746] <=  8'h00;      memory[64747] <=  8'h00;      memory[64748] <=  8'h00;      memory[64749] <=  8'h00;      memory[64750] <=  8'h00;      memory[64751] <=  8'h00;      memory[64752] <=  8'h00;      memory[64753] <=  8'h00;      memory[64754] <=  8'h00;      memory[64755] <=  8'h00;      memory[64756] <=  8'h00;      memory[64757] <=  8'h00;      memory[64758] <=  8'h00;      memory[64759] <=  8'h00;      memory[64760] <=  8'h00;      memory[64761] <=  8'h00;      memory[64762] <=  8'h00;      memory[64763] <=  8'h00;      memory[64764] <=  8'h00;      memory[64765] <=  8'h00;      memory[64766] <=  8'h00;      memory[64767] <=  8'h00;      memory[64768] <=  8'h00;      memory[64769] <=  8'h00;      memory[64770] <=  8'h00;      memory[64771] <=  8'h00;      memory[64772] <=  8'h00;      memory[64773] <=  8'h00;      memory[64774] <=  8'h00;      memory[64775] <=  8'h00;      memory[64776] <=  8'h00;      memory[64777] <=  8'h00;      memory[64778] <=  8'h00;      memory[64779] <=  8'h00;      memory[64780] <=  8'h00;      memory[64781] <=  8'h00;      memory[64782] <=  8'h00;      memory[64783] <=  8'h00;      memory[64784] <=  8'h00;      memory[64785] <=  8'h00;      memory[64786] <=  8'h00;      memory[64787] <=  8'h00;      memory[64788] <=  8'h00;      memory[64789] <=  8'h00;      memory[64790] <=  8'h00;      memory[64791] <=  8'h00;      memory[64792] <=  8'h00;      memory[64793] <=  8'h00;      memory[64794] <=  8'h00;      memory[64795] <=  8'h00;      memory[64796] <=  8'h00;      memory[64797] <=  8'h00;      memory[64798] <=  8'h00;      memory[64799] <=  8'h00;      memory[64800] <=  8'h00;      memory[64801] <=  8'h00;      memory[64802] <=  8'h00;      memory[64803] <=  8'h00;      memory[64804] <=  8'h00;      memory[64805] <=  8'h00;      memory[64806] <=  8'h00;      memory[64807] <=  8'h00;      memory[64808] <=  8'h00;      memory[64809] <=  8'h00;      memory[64810] <=  8'h00;      memory[64811] <=  8'h00;      memory[64812] <=  8'h00;      memory[64813] <=  8'h00;      memory[64814] <=  8'h00;      memory[64815] <=  8'h00;      memory[64816] <=  8'h00;      memory[64817] <=  8'h00;      memory[64818] <=  8'h00;      memory[64819] <=  8'h00;      memory[64820] <=  8'h00;      memory[64821] <=  8'h00;      memory[64822] <=  8'h00;      memory[64823] <=  8'h00;      memory[64824] <=  8'h00;      memory[64825] <=  8'h00;      memory[64826] <=  8'h00;      memory[64827] <=  8'h00;      memory[64828] <=  8'h00;      memory[64829] <=  8'h00;      memory[64830] <=  8'h00;      memory[64831] <=  8'h00;      memory[64832] <=  8'h00;      memory[64833] <=  8'h00;      memory[64834] <=  8'h00;      memory[64835] <=  8'h00;      memory[64836] <=  8'h00;      memory[64837] <=  8'h00;      memory[64838] <=  8'h00;      memory[64839] <=  8'h00;      memory[64840] <=  8'h00;      memory[64841] <=  8'h00;      memory[64842] <=  8'h00;      memory[64843] <=  8'h00;      memory[64844] <=  8'h00;      memory[64845] <=  8'h00;      memory[64846] <=  8'h00;      memory[64847] <=  8'h00;      memory[64848] <=  8'h00;      memory[64849] <=  8'h00;      memory[64850] <=  8'h00;      memory[64851] <=  8'h00;      memory[64852] <=  8'h00;      memory[64853] <=  8'h00;      memory[64854] <=  8'h00;      memory[64855] <=  8'h00;      memory[64856] <=  8'h00;      memory[64857] <=  8'h00;      memory[64858] <=  8'h00;      memory[64859] <=  8'h00;      memory[64860] <=  8'h00;      memory[64861] <=  8'h00;      memory[64862] <=  8'h00;      memory[64863] <=  8'h00;      memory[64864] <=  8'h00;      memory[64865] <=  8'h00;      memory[64866] <=  8'h00;      memory[64867] <=  8'h00;      memory[64868] <=  8'h00;      memory[64869] <=  8'h00;      memory[64870] <=  8'h00;      memory[64871] <=  8'h00;      memory[64872] <=  8'h00;      memory[64873] <=  8'h00;      memory[64874] <=  8'h00;      memory[64875] <=  8'h00;      memory[64876] <=  8'h00;      memory[64877] <=  8'h00;      memory[64878] <=  8'h00;      memory[64879] <=  8'h00;      memory[64880] <=  8'h00;      memory[64881] <=  8'h00;      memory[64882] <=  8'h00;      memory[64883] <=  8'h00;      memory[64884] <=  8'h00;      memory[64885] <=  8'h00;      memory[64886] <=  8'h00;      memory[64887] <=  8'h00;      memory[64888] <=  8'h00;      memory[64889] <=  8'h00;      memory[64890] <=  8'h00;      memory[64891] <=  8'h00;      memory[64892] <=  8'h00;      memory[64893] <=  8'h00;      memory[64894] <=  8'h00;      memory[64895] <=  8'h00;      memory[64896] <=  8'h00;      memory[64897] <=  8'h00;      memory[64898] <=  8'h00;      memory[64899] <=  8'h00;      memory[64900] <=  8'h00;      memory[64901] <=  8'h00;      memory[64902] <=  8'h00;      memory[64903] <=  8'h00;      memory[64904] <=  8'h00;      memory[64905] <=  8'h00;      memory[64906] <=  8'h00;      memory[64907] <=  8'h00;      memory[64908] <=  8'h00;      memory[64909] <=  8'h00;      memory[64910] <=  8'h00;      memory[64911] <=  8'h00;      memory[64912] <=  8'h00;      memory[64913] <=  8'h00;      memory[64914] <=  8'h00;      memory[64915] <=  8'h00;      memory[64916] <=  8'h00;      memory[64917] <=  8'h00;      memory[64918] <=  8'h00;      memory[64919] <=  8'h00;      memory[64920] <=  8'h00;      memory[64921] <=  8'h00;      memory[64922] <=  8'h00;      memory[64923] <=  8'h00;      memory[64924] <=  8'h00;      memory[64925] <=  8'h00;      memory[64926] <=  8'h00;      memory[64927] <=  8'h00;      memory[64928] <=  8'h00;      memory[64929] <=  8'h00;      memory[64930] <=  8'h00;      memory[64931] <=  8'h00;      memory[64932] <=  8'h00;      memory[64933] <=  8'h00;      memory[64934] <=  8'h00;      memory[64935] <=  8'h00;      memory[64936] <=  8'h00;      memory[64937] <=  8'h00;      memory[64938] <=  8'h00;      memory[64939] <=  8'h00;      memory[64940] <=  8'h00;      memory[64941] <=  8'h00;      memory[64942] <=  8'h00;      memory[64943] <=  8'h00;      memory[64944] <=  8'h00;      memory[64945] <=  8'h00;      memory[64946] <=  8'h00;      memory[64947] <=  8'h00;      memory[64948] <=  8'h00;      memory[64949] <=  8'h00;      memory[64950] <=  8'h00;      memory[64951] <=  8'h00;      memory[64952] <=  8'h00;      memory[64953] <=  8'h00;      memory[64954] <=  8'h00;      memory[64955] <=  8'h00;      memory[64956] <=  8'h00;      memory[64957] <=  8'h00;      memory[64958] <=  8'h00;      memory[64959] <=  8'h00;      memory[64960] <=  8'h00;      memory[64961] <=  8'h00;      memory[64962] <=  8'h00;      memory[64963] <=  8'h00;      memory[64964] <=  8'h00;      memory[64965] <=  8'h00;      memory[64966] <=  8'h00;      memory[64967] <=  8'h00;      memory[64968] <=  8'h00;      memory[64969] <=  8'h00;      memory[64970] <=  8'h00;      memory[64971] <=  8'h00;      memory[64972] <=  8'h00;      memory[64973] <=  8'h00;      memory[64974] <=  8'h00;      memory[64975] <=  8'h00;      memory[64976] <=  8'h00;      memory[64977] <=  8'h00;      memory[64978] <=  8'h00;      memory[64979] <=  8'h00;      memory[64980] <=  8'h00;      memory[64981] <=  8'h00;      memory[64982] <=  8'h00;      memory[64983] <=  8'h00;      memory[64984] <=  8'h00;      memory[64985] <=  8'h00;      memory[64986] <=  8'h00;      memory[64987] <=  8'h00;      memory[64988] <=  8'h00;      memory[64989] <=  8'h00;      memory[64990] <=  8'h00;      memory[64991] <=  8'h00;      memory[64992] <=  8'h00;      memory[64993] <=  8'h00;      memory[64994] <=  8'h00;      memory[64995] <=  8'h00;      memory[64996] <=  8'h00;      memory[64997] <=  8'h00;      memory[64998] <=  8'h00;      memory[64999] <=  8'h00;      memory[65000] <=  8'h00;      memory[65001] <=  8'h00;      memory[65002] <=  8'h00;      memory[65003] <=  8'h00;      memory[65004] <=  8'h00;      memory[65005] <=  8'h00;      memory[65006] <=  8'h00;      memory[65007] <=  8'h00;      memory[65008] <=  8'h00;      memory[65009] <=  8'h00;      memory[65010] <=  8'h00;      memory[65011] <=  8'h00;      memory[65012] <=  8'h00;      memory[65013] <=  8'h00;      memory[65014] <=  8'h00;      memory[65015] <=  8'h00;      memory[65016] <=  8'h00;      memory[65017] <=  8'h00;      memory[65018] <=  8'h00;      memory[65019] <=  8'h00;      memory[65020] <=  8'h00;      memory[65021] <=  8'h00;      memory[65022] <=  8'h00;      memory[65023] <=  8'h00;      memory[65024] <=  8'h00;      memory[65025] <=  8'h00;      memory[65026] <=  8'h00;      memory[65027] <=  8'h00;      memory[65028] <=  8'h00;      memory[65029] <=  8'h00;      memory[65030] <=  8'h00;      memory[65031] <=  8'h00;      memory[65032] <=  8'h00;      memory[65033] <=  8'h00;      memory[65034] <=  8'h00;      memory[65035] <=  8'h00;      memory[65036] <=  8'h00;      memory[65037] <=  8'h00;      memory[65038] <=  8'h00;      memory[65039] <=  8'h00;      memory[65040] <=  8'h00;      memory[65041] <=  8'h00;      memory[65042] <=  8'h00;      memory[65043] <=  8'h00;      memory[65044] <=  8'h00;      memory[65045] <=  8'h00;      memory[65046] <=  8'h00;      memory[65047] <=  8'h00;      memory[65048] <=  8'h00;      memory[65049] <=  8'h00;      memory[65050] <=  8'h00;      memory[65051] <=  8'h00;      memory[65052] <=  8'h00;      memory[65053] <=  8'h00;      memory[65054] <=  8'h00;      memory[65055] <=  8'h00;      memory[65056] <=  8'h00;      memory[65057] <=  8'h00;      memory[65058] <=  8'h00;      memory[65059] <=  8'h00;      memory[65060] <=  8'h00;      memory[65061] <=  8'h00;      memory[65062] <=  8'h00;      memory[65063] <=  8'h00;      memory[65064] <=  8'h00;      memory[65065] <=  8'h00;      memory[65066] <=  8'h00;      memory[65067] <=  8'h00;      memory[65068] <=  8'h00;      memory[65069] <=  8'h00;      memory[65070] <=  8'h00;      memory[65071] <=  8'h00;      memory[65072] <=  8'h00;      memory[65073] <=  8'h00;      memory[65074] <=  8'h00;      memory[65075] <=  8'h00;      memory[65076] <=  8'h00;      memory[65077] <=  8'h00;      memory[65078] <=  8'h00;      memory[65079] <=  8'h00;      memory[65080] <=  8'h00;      memory[65081] <=  8'h00;      memory[65082] <=  8'h00;      memory[65083] <=  8'h00;      memory[65084] <=  8'h00;      memory[65085] <=  8'h00;      memory[65086] <=  8'h00;      memory[65087] <=  8'h00;      memory[65088] <=  8'h00;      memory[65089] <=  8'h00;      memory[65090] <=  8'h00;      memory[65091] <=  8'h00;      memory[65092] <=  8'h00;      memory[65093] <=  8'h00;      memory[65094] <=  8'h00;      memory[65095] <=  8'h00;      memory[65096] <=  8'h00;      memory[65097] <=  8'h00;      memory[65098] <=  8'h00;      memory[65099] <=  8'h00;      memory[65100] <=  8'h00;      memory[65101] <=  8'h00;      memory[65102] <=  8'h00;      memory[65103] <=  8'h00;      memory[65104] <=  8'h00;      memory[65105] <=  8'h00;      memory[65106] <=  8'h00;      memory[65107] <=  8'h00;      memory[65108] <=  8'h00;      memory[65109] <=  8'h00;      memory[65110] <=  8'h00;      memory[65111] <=  8'h00;      memory[65112] <=  8'h00;      memory[65113] <=  8'h00;      memory[65114] <=  8'h00;      memory[65115] <=  8'h00;      memory[65116] <=  8'h00;      memory[65117] <=  8'h00;      memory[65118] <=  8'h00;      memory[65119] <=  8'h00;      memory[65120] <=  8'h00;      memory[65121] <=  8'h00;      memory[65122] <=  8'h00;      memory[65123] <=  8'h00;      memory[65124] <=  8'h00;      memory[65125] <=  8'h00;      memory[65126] <=  8'h00;      memory[65127] <=  8'h00;      memory[65128] <=  8'h00;      memory[65129] <=  8'h00;      memory[65130] <=  8'h00;      memory[65131] <=  8'h00;      memory[65132] <=  8'h00;      memory[65133] <=  8'h00;      memory[65134] <=  8'h00;      memory[65135] <=  8'h00;      memory[65136] <=  8'h00;      memory[65137] <=  8'h00;      memory[65138] <=  8'h00;      memory[65139] <=  8'h00;      memory[65140] <=  8'h00;      memory[65141] <=  8'h00;      memory[65142] <=  8'h00;      memory[65143] <=  8'h00;      memory[65144] <=  8'h00;      memory[65145] <=  8'h00;      memory[65146] <=  8'h00;      memory[65147] <=  8'h00;      memory[65148] <=  8'h00;      memory[65149] <=  8'h00;      memory[65150] <=  8'h00;      memory[65151] <=  8'h00;      memory[65152] <=  8'h00;      memory[65153] <=  8'h00;      memory[65154] <=  8'h00;      memory[65155] <=  8'h00;      memory[65156] <=  8'h00;      memory[65157] <=  8'h00;      memory[65158] <=  8'h00;      memory[65159] <=  8'h00;      memory[65160] <=  8'h00;      memory[65161] <=  8'h00;      memory[65162] <=  8'h00;      memory[65163] <=  8'h00;      memory[65164] <=  8'h00;      memory[65165] <=  8'h00;      memory[65166] <=  8'h00;      memory[65167] <=  8'h00;      memory[65168] <=  8'h00;      memory[65169] <=  8'h00;      memory[65170] <=  8'h00;      memory[65171] <=  8'h00;      memory[65172] <=  8'h00;      memory[65173] <=  8'h00;      memory[65174] <=  8'h00;      memory[65175] <=  8'h00;      memory[65176] <=  8'h00;      memory[65177] <=  8'h00;      memory[65178] <=  8'h00;      memory[65179] <=  8'h00;      memory[65180] <=  8'h00;      memory[65181] <=  8'h00;      memory[65182] <=  8'h00;      memory[65183] <=  8'h00;      memory[65184] <=  8'h00;      memory[65185] <=  8'h00;      memory[65186] <=  8'h00;      memory[65187] <=  8'h00;      memory[65188] <=  8'h00;      memory[65189] <=  8'h00;      memory[65190] <=  8'h00;      memory[65191] <=  8'h00;      memory[65192] <=  8'h00;      memory[65193] <=  8'h00;      memory[65194] <=  8'h00;      memory[65195] <=  8'h00;      memory[65196] <=  8'h00;      memory[65197] <=  8'h00;      memory[65198] <=  8'h00;      memory[65199] <=  8'h00;      memory[65200] <=  8'h00;      memory[65201] <=  8'h00;      memory[65202] <=  8'h00;      memory[65203] <=  8'h00;      memory[65204] <=  8'h00;      memory[65205] <=  8'h00;      memory[65206] <=  8'h00;      memory[65207] <=  8'h00;      memory[65208] <=  8'h00;      memory[65209] <=  8'h00;      memory[65210] <=  8'h00;      memory[65211] <=  8'h00;      memory[65212] <=  8'h00;      memory[65213] <=  8'h00;      memory[65214] <=  8'h00;      memory[65215] <=  8'h00;      memory[65216] <=  8'h00;      memory[65217] <=  8'h00;      memory[65218] <=  8'h00;      memory[65219] <=  8'h00;      memory[65220] <=  8'h00;      memory[65221] <=  8'h00;      memory[65222] <=  8'h00;      memory[65223] <=  8'h00;      memory[65224] <=  8'h00;      memory[65225] <=  8'h00;      memory[65226] <=  8'h00;      memory[65227] <=  8'h00;      memory[65228] <=  8'h00;      memory[65229] <=  8'h00;      memory[65230] <=  8'h00;      memory[65231] <=  8'h00;      memory[65232] <=  8'h00;      memory[65233] <=  8'h00;      memory[65234] <=  8'h00;      memory[65235] <=  8'h00;      memory[65236] <=  8'h00;      memory[65237] <=  8'h00;      memory[65238] <=  8'h00;      memory[65239] <=  8'h00;      memory[65240] <=  8'h00;      memory[65241] <=  8'h00;      memory[65242] <=  8'h00;      memory[65243] <=  8'h00;      memory[65244] <=  8'h00;      memory[65245] <=  8'h00;      memory[65246] <=  8'h00;      memory[65247] <=  8'h00;      memory[65248] <=  8'h00;      memory[65249] <=  8'h00;      memory[65250] <=  8'h00;      memory[65251] <=  8'h00;      memory[65252] <=  8'h00;      memory[65253] <=  8'h00;      memory[65254] <=  8'h00;      memory[65255] <=  8'h00;      memory[65256] <=  8'h00;      memory[65257] <=  8'h00;      memory[65258] <=  8'h00;      memory[65259] <=  8'h00;      memory[65260] <=  8'h00;      memory[65261] <=  8'h00;      memory[65262] <=  8'h00;      memory[65263] <=  8'h00;      memory[65264] <=  8'h00;      memory[65265] <=  8'h00;      memory[65266] <=  8'h00;      memory[65267] <=  8'h00;      memory[65268] <=  8'h00;      memory[65269] <=  8'h00;      memory[65270] <=  8'h00;      memory[65271] <=  8'h00;      memory[65272] <=  8'h00;      memory[65273] <=  8'h00;      memory[65274] <=  8'h00;      memory[65275] <=  8'h00;      memory[65276] <=  8'h00;      memory[65277] <=  8'h00;      memory[65278] <=  8'h00;      memory[65279] <=  8'h00;      memory[65280] <=  8'h00;      memory[65281] <=  8'h00;      memory[65282] <=  8'h00;      memory[65283] <=  8'h00;      memory[65284] <=  8'h00;      memory[65285] <=  8'h00;      memory[65286] <=  8'h00;      memory[65287] <=  8'h00;      memory[65288] <=  8'h00;      memory[65289] <=  8'h00;      memory[65290] <=  8'h00;      memory[65291] <=  8'h00;      memory[65292] <=  8'h00;      memory[65293] <=  8'h00;      memory[65294] <=  8'h00;      memory[65295] <=  8'h00;      memory[65296] <=  8'h00;      memory[65297] <=  8'h00;      memory[65298] <=  8'h00;      memory[65299] <=  8'h00;      memory[65300] <=  8'h00;      memory[65301] <=  8'h00;      memory[65302] <=  8'h00;      memory[65303] <=  8'h00;      memory[65304] <=  8'h00;      memory[65305] <=  8'h00;      memory[65306] <=  8'h00;      memory[65307] <=  8'h00;      memory[65308] <=  8'h00;      memory[65309] <=  8'h00;      memory[65310] <=  8'h00;      memory[65311] <=  8'h00;      memory[65312] <=  8'h00;      memory[65313] <=  8'h00;      memory[65314] <=  8'h00;      memory[65315] <=  8'h00;      memory[65316] <=  8'h00;      memory[65317] <=  8'h00;      memory[65318] <=  8'h00;      memory[65319] <=  8'h00;      memory[65320] <=  8'h00;      memory[65321] <=  8'h00;      memory[65322] <=  8'h00;      memory[65323] <=  8'h00;      memory[65324] <=  8'h00;      memory[65325] <=  8'h00;      memory[65326] <=  8'h00;      memory[65327] <=  8'h00;      memory[65328] <=  8'h00;      memory[65329] <=  8'h00;      memory[65330] <=  8'h00;      memory[65331] <=  8'h00;      memory[65332] <=  8'h00;      memory[65333] <=  8'h00;      memory[65334] <=  8'h00;      memory[65335] <=  8'h00;      memory[65336] <=  8'h00;      memory[65337] <=  8'h00;      memory[65338] <=  8'h00;      memory[65339] <=  8'h00;      memory[65340] <=  8'h00;      memory[65341] <=  8'h00;      memory[65342] <=  8'h00;      memory[65343] <=  8'h00;      memory[65344] <=  8'h00;      memory[65345] <=  8'h00;      memory[65346] <=  8'h00;      memory[65347] <=  8'h00;      memory[65348] <=  8'h00;      memory[65349] <=  8'h00;      memory[65350] <=  8'h00;      memory[65351] <=  8'h00;      memory[65352] <=  8'h00;      memory[65353] <=  8'h00;      memory[65354] <=  8'h00;      memory[65355] <=  8'h00;      memory[65356] <=  8'h00;      memory[65357] <=  8'h00;      memory[65358] <=  8'h00;      memory[65359] <=  8'h00;      memory[65360] <=  8'h00;      memory[65361] <=  8'h00;      memory[65362] <=  8'h00;      memory[65363] <=  8'h00;      memory[65364] <=  8'h00;      memory[65365] <=  8'h00;      memory[65366] <=  8'h00;      memory[65367] <=  8'h00;      memory[65368] <=  8'h00;      memory[65369] <=  8'h00;      memory[65370] <=  8'h00;      memory[65371] <=  8'h00;      memory[65372] <=  8'h00;      memory[65373] <=  8'h00;      memory[65374] <=  8'h00;      memory[65375] <=  8'h00;      memory[65376] <=  8'h00;      memory[65377] <=  8'h00;      memory[65378] <=  8'h00;      memory[65379] <=  8'h00;      memory[65380] <=  8'h00;      memory[65381] <=  8'h00;      memory[65382] <=  8'h00;      memory[65383] <=  8'h00;      memory[65384] <=  8'h00;      memory[65385] <=  8'h00;      memory[65386] <=  8'h00;      memory[65387] <=  8'h00;      memory[65388] <=  8'h00;      memory[65389] <=  8'h00;      memory[65390] <=  8'h00;      memory[65391] <=  8'h00;      memory[65392] <=  8'h00;      memory[65393] <=  8'h00;      memory[65394] <=  8'h00;      memory[65395] <=  8'h00;      memory[65396] <=  8'h00;      memory[65397] <=  8'h00;      memory[65398] <=  8'h00;      memory[65399] <=  8'h00;      memory[65400] <=  8'h00;      memory[65401] <=  8'h00;      memory[65402] <=  8'h00;      memory[65403] <=  8'h00;      memory[65404] <=  8'h00;      memory[65405] <=  8'h00;      memory[65406] <=  8'h00;      memory[65407] <=  8'h00;      memory[65408] <=  8'h00;      memory[65409] <=  8'h00;      memory[65410] <=  8'h00;      memory[65411] <=  8'h00;      memory[65412] <=  8'h00;      memory[65413] <=  8'h00;      memory[65414] <=  8'h00;      memory[65415] <=  8'h00;      memory[65416] <=  8'h00;      memory[65417] <=  8'h00;      memory[65418] <=  8'h00;      memory[65419] <=  8'h00;      memory[65420] <=  8'h00;      memory[65421] <=  8'h00;      memory[65422] <=  8'h00;      memory[65423] <=  8'h00;      memory[65424] <=  8'h00;      memory[65425] <=  8'h00;      memory[65426] <=  8'h00;      memory[65427] <=  8'h00;      memory[65428] <=  8'h00;      memory[65429] <=  8'h00;      memory[65430] <=  8'h00;      memory[65431] <=  8'h00;      memory[65432] <=  8'h00;      memory[65433] <=  8'h00;      memory[65434] <=  8'h00;      memory[65435] <=  8'h00;      memory[65436] <=  8'h00;      memory[65437] <=  8'h00;      memory[65438] <=  8'h00;      memory[65439] <=  8'h00;      memory[65440] <=  8'h00;      memory[65441] <=  8'h00;      memory[65442] <=  8'h00;      memory[65443] <=  8'h00;      memory[65444] <=  8'h00;      memory[65445] <=  8'h00;      memory[65446] <=  8'h00;      memory[65447] <=  8'h00;      memory[65448] <=  8'h00;      memory[65449] <=  8'h00;      memory[65450] <=  8'h00;      memory[65451] <=  8'h00;      memory[65452] <=  8'h00;      memory[65453] <=  8'h00;      memory[65454] <=  8'h00;      memory[65455] <=  8'h00;      memory[65456] <=  8'h00;      memory[65457] <=  8'h00;      memory[65458] <=  8'h00;      memory[65459] <=  8'h00;      memory[65460] <=  8'h00;      memory[65461] <=  8'h00;      memory[65462] <=  8'h00;      memory[65463] <=  8'h00;      memory[65464] <=  8'h00;      memory[65465] <=  8'h00;      memory[65466] <=  8'h00;      memory[65467] <=  8'h00;      memory[65468] <=  8'h00;      memory[65469] <=  8'h00;      memory[65470] <=  8'h00;      memory[65471] <=  8'h00;      memory[65472] <=  8'h00;      memory[65473] <=  8'h00;      memory[65474] <=  8'h00;      memory[65475] <=  8'h00;      memory[65476] <=  8'h00;      memory[65477] <=  8'h00;      memory[65478] <=  8'h00;      memory[65479] <=  8'h00;      memory[65480] <=  8'h00;      memory[65481] <=  8'h00;      memory[65482] <=  8'h00;      memory[65483] <=  8'h00;      memory[65484] <=  8'h00;      memory[65485] <=  8'h00;      memory[65486] <=  8'h00;      memory[65487] <=  8'h00;      memory[65488] <=  8'h00;      memory[65489] <=  8'h00;      memory[65490] <=  8'h00;      memory[65491] <=  8'h00;      memory[65492] <=  8'h00;      memory[65493] <=  8'h00;      memory[65494] <=  8'h00;      memory[65495] <=  8'h00;      memory[65496] <=  8'h00;      memory[65497] <=  8'h00;      memory[65498] <=  8'h00;      memory[65499] <=  8'h00;      memory[65500] <=  8'h00;      memory[65501] <=  8'h00;      memory[65502] <=  8'h00;      memory[65503] <=  8'h00;      memory[65504] <=  8'h00;      memory[65505] <=  8'h00;      memory[65506] <=  8'h00;      memory[65507] <=  8'h00;      memory[65508] <=  8'h00;      memory[65509] <=  8'h00;      memory[65510] <=  8'h00;      memory[65511] <=  8'h00;      memory[65512] <=  8'h00;      memory[65513] <=  8'h00;      memory[65514] <=  8'h00;      memory[65515] <=  8'h00;      memory[65516] <=  8'h00;      memory[65517] <=  8'h00;      memory[65518] <=  8'h00;      memory[65519] <=  8'h00;      memory[65520] <=  8'h00;      memory[65521] <=  8'h00;      memory[65522] <=  8'h00;      memory[65523] <=  8'h00;      memory[65524] <=  8'h00;      memory[65525] <=  8'h00;      memory[65526] <=  8'h00;      memory[65527] <=  8'h00;      memory[65528] <=  8'h00;      memory[65529] <=  8'h00;      memory[65530] <=  8'h00;      memory[65531] <=  8'h00;      memory[65532] <=  8'h00;      memory[65533] <=  8'h00;      memory[65534] <=  8'h00;      memory[65535] <=  8'h00;  
    end

    always @(posedge clk) begin
        if (enable) begin
            if (we) begin
                memory[addr] <= write_data; // Write operation when we and enable are high
                reg_last_written_data <= write_data;
                reg_last_written_addr <= addr;
            end
        read_data_buff2  <= memory[addr]; // Read operation when enable is high
            read_data_buff1  <= read_data_buff2; // Read operation when enable is high
            read_data <= read_data_buff1; // Read operation when enable is high

        end
    end
 
endmodule
